module fake_netlist_6_1850_n_1988 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1988);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1988;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1890;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g190 ( 
.A(n_54),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_18),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_8),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_93),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_41),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_14),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_52),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_66),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_69),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_34),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_106),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_1),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_99),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_64),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_23),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_71),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_33),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_92),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_10),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_78),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_124),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_90),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_128),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_87),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_169),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_68),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_139),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_89),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_112),
.Y(n_260)
);

BUFx8_ASAP7_75t_SL g261 ( 
.A(n_34),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_29),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_61),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_135),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_149),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_182),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_130),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_95),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_19),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_189),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_137),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_172),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_140),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_116),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_21),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_100),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_119),
.Y(n_281)
);

BUFx2_ASAP7_75t_R g282 ( 
.A(n_132),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_122),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_117),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_143),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_3),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_120),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_160),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_159),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_28),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_144),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_50),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_79),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_68),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_105),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_65),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_158),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_48),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_91),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_17),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_138),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_47),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_40),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_70),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_80),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_24),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_42),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_67),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_75),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_14),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_35),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_185),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_57),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_39),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_65),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_157),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_43),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_154),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_11),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_129),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_101),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_152),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_57),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_7),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_4),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_51),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_126),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_55),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_20),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_162),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_150),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_48),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_155),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_71),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_102),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_164),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_175),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_15),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_60),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_51),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_148),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_43),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_186),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_181),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_125),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_45),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_59),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_134),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_84),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_81),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_45),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_83),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_82),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_73),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_127),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_72),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_103),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_0),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_38),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_4),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_114),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_22),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_12),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_0),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_156),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_280),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_280),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_291),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_331),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_280),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_280),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_261),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_280),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_300),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_330),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_334),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_300),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_237),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_361),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_239),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_242),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_300),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_248),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_300),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_307),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_243),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_200),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_254),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_246),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_247),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_304),
.B(n_2),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_259),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_307),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_264),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_191),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_307),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_276),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_289),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_290),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_359),
.B(n_5),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_353),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_319),
.B(n_9),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_249),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_251),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_299),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_197),
.B(n_9),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_320),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_320),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_190),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_252),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_253),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_301),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_257),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_193),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_265),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_305),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_204),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_306),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_207),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_266),
.B(n_133),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_309),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_313),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_304),
.B(n_11),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_316),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_220),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_211),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_317),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_259),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_236),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_267),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_235),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_238),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_269),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_271),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_241),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_372),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_244),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_273),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_274),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_250),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_256),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_209),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_209),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_216),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_216),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_311),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_223),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_321),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_323),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_411),
.B(n_304),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_318),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_412),
.B(n_375),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_450),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_349),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_412),
.B(n_453),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_405),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_279),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_349),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_233),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_424),
.B(n_233),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_424),
.B(n_357),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_390),
.B(n_196),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_392),
.B(n_395),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_469),
.A2(n_342),
.B(n_311),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_469),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_470),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_471),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_472),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_421),
.B(n_282),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_382),
.B(n_245),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_386),
.B(n_319),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_260),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_466),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_454),
.B(n_196),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_421),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_384),
.A2(n_194),
.B1(n_201),
.B2(n_377),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_398),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_473),
.B(n_202),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_399),
.B(n_202),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_SL g555 ( 
.A(n_481),
.B(n_397),
.C(n_399),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_492),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_532),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_515),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_481),
.B(n_401),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_407),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_515),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_507),
.B(n_222),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_551),
.B(n_422),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_549),
.B(n_407),
.Y(n_567)
);

INVx6_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_414),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_554),
.B(n_408),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_522),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_492),
.B(n_383),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_522),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_529),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_536),
.B(n_417),
.C(n_414),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_477),
.B(n_245),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_515),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_494),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_491),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_517),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_491),
.B(n_417),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_494),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_517),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_552),
.A2(n_426),
.B1(n_427),
.B2(n_409),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_550),
.B(n_385),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_549),
.B(n_551),
.Y(n_593)
);

AND3x2_ASAP7_75t_L g594 ( 
.A(n_529),
.B(n_302),
.C(n_293),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_536),
.B(n_420),
.C(n_418),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_487),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_487),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_551),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_507),
.A2(n_342),
.B1(n_378),
.B2(n_341),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_491),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_532),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_532),
.Y(n_604)
);

AND3x2_ASAP7_75t_L g605 ( 
.A(n_518),
.B(n_302),
.C(n_293),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_303),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_507),
.B(n_303),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_491),
.B(n_507),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_518),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_503),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g615 ( 
.A1(n_548),
.A2(n_315),
.B1(n_327),
.B2(n_324),
.Y(n_615)
);

INVx8_ASAP7_75t_L g616 ( 
.A(n_504),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_552),
.B(n_554),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_488),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_552),
.B(n_461),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_552),
.A2(n_434),
.B1(n_437),
.B2(n_433),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_549),
.B(n_418),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_476),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_553),
.B(n_420),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_255),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_488),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_502),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_531),
.B(n_428),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_500),
.B(n_428),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_500),
.B(n_435),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_553),
.B(n_389),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_534),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_550),
.B(n_394),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_548),
.B(n_439),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_499),
.B(n_455),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_500),
.B(n_435),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_488),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_495),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_488),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_504),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_531),
.B(n_440),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_504),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_477),
.B(n_440),
.Y(n_656)
);

OAI21xp33_ASAP7_75t_SL g657 ( 
.A1(n_499),
.A2(n_270),
.B(n_262),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_477),
.A2(n_294),
.B1(n_278),
.B2(n_288),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_478),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_511),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_539),
.B(n_292),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_509),
.B(n_458),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_511),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_504),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_478),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_539),
.B(n_326),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_479),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_518),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_542),
.B(n_442),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_487),
.B(n_284),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_479),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_539),
.B(n_543),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_482),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_542),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_489),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_477),
.B(n_442),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_SL g680 ( 
.A(n_509),
.B(n_195),
.C(n_191),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_482),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_504),
.B(n_490),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_489),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_487),
.B(n_447),
.C(n_446),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_504),
.A2(n_345),
.B1(n_337),
.B2(n_352),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_542),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_482),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_483),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_543),
.A2(n_372),
.B1(n_368),
.B2(n_195),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_495),
.B(n_459),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_504),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_531),
.B(n_192),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_490),
.B(n_446),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_483),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_489),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_535),
.A2(n_436),
.B1(n_444),
.B2(n_463),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_516),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_504),
.B(n_447),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_483),
.Y(n_701)
);

AND2x6_ASAP7_75t_L g702 ( 
.A(n_490),
.B(n_255),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_504),
.B(n_449),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_535),
.A2(n_465),
.B1(n_464),
.B2(n_475),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_484),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_531),
.B(n_449),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_660),
.B(n_504),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_660),
.B(n_480),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_602),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_556),
.B(n_452),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_607),
.A2(n_277),
.B1(n_258),
.B2(n_224),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_587),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_580),
.B(n_220),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_618),
.A2(n_516),
.B1(n_452),
.B2(n_475),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_634),
.B(n_474),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_602),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_SL g718 ( 
.A(n_575),
.B(n_255),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_630),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_664),
.B(n_480),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_630),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_607),
.A2(n_474),
.B1(n_295),
.B2(n_287),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_580),
.B(n_220),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_612),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_612),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_255),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_664),
.B(n_480),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_675),
.B(n_539),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_636),
.B(n_535),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_579),
.B(n_537),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_582),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_627),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_568),
.Y(n_734)
);

AND2x2_ASAP7_75t_SL g735 ( 
.A(n_642),
.B(n_255),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_568),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_584),
.B(n_480),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_650),
.B(n_272),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_590),
.B(n_368),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_609),
.B(n_480),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_627),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_555),
.A2(n_332),
.B1(n_360),
.B2(n_363),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_687),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_SL g744 ( 
.A1(n_628),
.A2(n_339),
.B1(n_210),
.B2(n_212),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_568),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_568),
.Y(n_746)
);

O2A1O1Ixp5_ASAP7_75t_L g747 ( 
.A1(n_562),
.A2(n_486),
.B(n_484),
.C(n_493),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_573),
.B(n_537),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_661),
.B(n_537),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_597),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_687),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_563),
.A2(n_272),
.B1(n_308),
.B2(n_358),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_613),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_645),
.B(n_205),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_609),
.B(n_480),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_593),
.A2(n_538),
.B(n_533),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_587),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_613),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_597),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_616),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_632),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_650),
.B(n_272),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_596),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_650),
.B(n_272),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_614),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_526),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_205),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_600),
.B(n_214),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_632),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_614),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_599),
.B(n_526),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_611),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_600),
.B(n_214),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_671),
.B(n_272),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_557),
.B(n_526),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_694),
.B(n_541),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_663),
.A2(n_275),
.B1(n_379),
.B2(n_296),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_603),
.B(n_526),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_571),
.A2(n_310),
.B1(n_285),
.B2(n_312),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_604),
.B(n_526),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_596),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_638),
.B(n_526),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_620),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_684),
.B(n_486),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_600),
.B(n_217),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_578),
.A2(n_338),
.B1(n_210),
.B2(n_212),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_693),
.B(n_575),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_656),
.B(n_217),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_671),
.B(n_308),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_575),
.B(n_486),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_575),
.B(n_493),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_560),
.B(n_493),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_679),
.B(n_218),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_563),
.A2(n_501),
.B(n_506),
.C(n_505),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_567),
.B(n_501),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_671),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_631),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_569),
.B(n_501),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_651),
.A2(n_322),
.B1(n_298),
.B2(n_370),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_623),
.B(n_506),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_595),
.B(n_218),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_580),
.B(n_220),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_565),
.B(n_506),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_565),
.B(n_508),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_608),
.B(n_308),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_617),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_673),
.B(n_221),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_651),
.B(n_541),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_685),
.B(n_198),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_570),
.B(n_508),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_570),
.B(n_508),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_707),
.B(n_221),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_572),
.B(n_513),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_641),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_572),
.B(n_513),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_564),
.B(n_544),
.C(n_541),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_617),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_558),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_574),
.B(n_513),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_608),
.B(n_308),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_564),
.B(n_546),
.C(n_544),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_707),
.B(n_546),
.C(n_544),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_580),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_694),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_608),
.B(n_308),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_666),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_648),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_558),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_668),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_622),
.A2(n_338),
.B1(n_213),
.B2(n_376),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_699),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_610),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_700),
.A2(n_231),
.B1(n_203),
.B2(n_206),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_574),
.A2(n_547),
.B(n_546),
.C(n_530),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_619),
.B(n_694),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_668),
.B(n_514),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_670),
.Y(n_840)
);

NAND2x1p5_ASAP7_75t_L g841 ( 
.A(n_654),
.B(n_215),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_608),
.B(n_358),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_561),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_670),
.B(n_514),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_674),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_561),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_625),
.B(n_225),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_674),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_704),
.B(n_547),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_608),
.B(n_358),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_657),
.A2(n_547),
.B(n_530),
.C(n_524),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_703),
.B(n_358),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_601),
.A2(n_213),
.B(n_199),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_673),
.A2(n_356),
.B1(n_225),
.B2(n_228),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_676),
.B(n_514),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_605),
.B(n_545),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_676),
.B(n_519),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_616),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_681),
.Y(n_859)
);

NAND2x1_ASAP7_75t_L g860 ( 
.A(n_654),
.B(n_505),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_594),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_691),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_566),
.B(n_228),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_559),
.B(n_533),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_682),
.B(n_358),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_229),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_621),
.B(n_229),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_705),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_705),
.B(n_629),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_654),
.B(n_220),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_665),
.B(n_220),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_629),
.B(n_519),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_658),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_624),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_629),
.B(n_519),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_810),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_817),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_750),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_730),
.B(n_580),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_743),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_768),
.A2(n_669),
.B(n_677),
.C(n_672),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_768),
.A2(n_616),
.B(n_690),
.C(n_680),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_817),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_838),
.A2(n_616),
.B(n_665),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_711),
.B(n_811),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_750),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_730),
.B(n_580),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_761),
.A2(n_692),
.B(n_665),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_750),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_735),
.A2(n_753),
.B1(n_874),
.B2(n_712),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_750),
.B(n_799),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_755),
.B(n_606),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_862),
.B(n_698),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_755),
.B(n_606),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_719),
.B(n_606),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_837),
.A2(n_615),
.B(n_701),
.C(n_696),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_735),
.A2(n_686),
.B1(n_692),
.B2(n_658),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_716),
.A2(n_606),
.B1(n_692),
.B2(n_637),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_732),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_721),
.B(n_606),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_761),
.A2(n_649),
.B(n_644),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_716),
.B(n_606),
.Y(n_903)
);

CKINVDCx10_ASAP7_75t_R g904 ( 
.A(n_749),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_793),
.A2(n_794),
.B(n_799),
.Y(n_905)
);

BUFx2_ASAP7_75t_SL g906 ( 
.A(n_835),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_799),
.B(n_858),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_L g908 ( 
.A1(n_739),
.A2(n_219),
.B(n_199),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_799),
.A2(n_649),
.B(n_644),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_789),
.A2(n_646),
.B(n_635),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_764),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_827),
.B(n_661),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_778),
.B(n_661),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_837),
.A2(n_706),
.B(n_624),
.C(n_701),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_762),
.B(n_770),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_710),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_717),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_791),
.B(n_658),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_797),
.A2(n_646),
.B(n_635),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_733),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_791),
.B(n_658),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_751),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_858),
.A2(n_649),
.B(n_644),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_851),
.A2(n_706),
.B(n_633),
.C(n_696),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_858),
.B(n_577),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_764),
.B(n_661),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_713),
.B(n_667),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_858),
.A2(n_592),
.B(n_577),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_737),
.A2(n_592),
.B(n_577),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_728),
.B(n_667),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_783),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_796),
.B(n_753),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_769),
.B(n_775),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_796),
.B(n_633),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_760),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_830),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_708),
.B(n_577),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_865),
.A2(n_646),
.B(n_635),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_733),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_740),
.A2(n_592),
.B(n_577),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_733),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_773),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_865),
.A2(n_234),
.B(n_230),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_733),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_774),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_758),
.B(n_667),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_826),
.B(n_647),
.Y(n_947)
);

NOR2x1p5_ASAP7_75t_L g948 ( 
.A(n_748),
.B(n_219),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_741),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_752),
.B(n_667),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_829),
.B(n_639),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_756),
.B(n_592),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_832),
.B(n_652),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_741),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_840),
.B(n_652),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_815),
.B(n_583),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_845),
.B(n_659),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_795),
.A2(n_592),
.B(n_647),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_815),
.A2(n_227),
.B(n_226),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_785),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_834),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_798),
.A2(n_647),
.B(n_678),
.Y(n_962)
);

INVx11_ASAP7_75t_L g963 ( 
.A(n_726),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_848),
.B(n_659),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_859),
.B(n_688),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_801),
.A2(n_697),
.B(n_678),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_741),
.B(n_688),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_790),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_866),
.B(n_689),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_869),
.B(n_689),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_800),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_769),
.B(n_591),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_729),
.B(n_591),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_741),
.B(n_841),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_775),
.B(n_640),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_803),
.A2(n_697),
.B(n_678),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_864),
.B(n_678),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_757),
.A2(n_655),
.B(n_653),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_709),
.B(n_678),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_833),
.B(n_588),
.C(n_335),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_778),
.B(n_720),
.Y(n_982)
);

AO21x1_ASAP7_75t_L g983 ( 
.A1(n_738),
.A2(n_263),
.B(n_240),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_874),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_806),
.A2(n_697),
.B(n_655),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_826),
.Y(n_986)
);

AO22x1_ASAP7_75t_L g987 ( 
.A1(n_804),
.A2(n_226),
.B1(n_376),
.B2(n_374),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_852),
.A2(n_655),
.B(n_653),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_807),
.A2(n_814),
.B(n_813),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_816),
.A2(n_697),
.B(n_662),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_787),
.B(n_640),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_697),
.B(n_653),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_727),
.B(n_662),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_787),
.B(n_662),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_822),
.A2(n_683),
.B(n_589),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_749),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_734),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_833),
.B(n_227),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_868),
.B(n_847),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_734),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_731),
.B(n_683),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_870),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_767),
.B(n_683),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_772),
.B(n_702),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_849),
.B(n_576),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_722),
.B(n_533),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_841),
.A2(n_586),
.B(n_581),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_715),
.B(n_533),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_875),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_L g1010 ( 
.A(n_726),
.B(n_626),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_742),
.A2(n_702),
.B1(n_626),
.B2(n_220),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_736),
.B(n_576),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_821),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_825),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_804),
.B(n_861),
.C(n_765),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_860),
.A2(n_598),
.B(n_589),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_852),
.A2(n_598),
.B(n_586),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_871),
.A2(n_585),
.B(n_581),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_839),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_872),
.A2(n_585),
.B(n_485),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_867),
.A2(n_702),
.B1(n_626),
.B2(n_268),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_831),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_868),
.A2(n_281),
.B(n_346),
.C(n_366),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_747),
.A2(n_626),
.B(n_702),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_873),
.A2(n_505),
.B(n_512),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_867),
.B(n_702),
.Y(n_1026)
);

AOI33xp33_ASAP7_75t_L g1027 ( 
.A1(n_788),
.A2(n_530),
.A3(n_524),
.B1(n_521),
.B2(n_545),
.B3(n_538),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_763),
.A2(n_497),
.B(n_485),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_853),
.A2(n_232),
.B(n_328),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_736),
.B(n_220),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_843),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_745),
.B(n_354),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_847),
.A2(n_325),
.B(n_283),
.C(n_314),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_863),
.B(n_702),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_763),
.A2(n_626),
.B(n_369),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_749),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_846),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_844),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_863),
.B(n_626),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_819),
.A2(n_333),
.B(n_540),
.C(n_538),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_745),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_786),
.B(n_538),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_824),
.A2(n_335),
.B1(n_364),
.B2(n_356),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_765),
.A2(n_485),
.B(n_497),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_776),
.A2(n_485),
.B(n_497),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_776),
.A2(n_497),
.B(n_505),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_856),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_R g1048 ( 
.A(n_856),
.B(n_232),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_792),
.A2(n_505),
.B(n_540),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_810),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_746),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_792),
.A2(n_545),
.B(n_540),
.C(n_521),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_742),
.A2(n_354),
.B1(n_328),
.B2(n_336),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_724),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_725),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_855),
.B(n_540),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_754),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_802),
.A2(n_286),
.B(n_336),
.Y(n_1058)
);

BUFx2_ASAP7_75t_SL g1059 ( 
.A(n_746),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_714),
.A2(n_505),
.B(n_545),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_723),
.A2(n_805),
.B(n_876),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_779),
.A2(n_348),
.B1(n_350),
.B2(n_329),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_777),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_812),
.A2(n_340),
.B1(n_364),
.B2(n_367),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_788),
.B(n_286),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_906),
.B(n_780),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_975),
.A2(n_784),
.B(n_782),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_881),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_984),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_922),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_989),
.A2(n_857),
.B(n_808),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_877),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_999),
.A2(n_781),
.B(n_854),
.C(n_836),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1019),
.B(n_759),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_905),
.A2(n_850),
.B(n_842),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_879),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1038),
.B(n_766),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_932),
.A2(n_850),
.B(n_842),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_935),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_942),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_984),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1025),
.A2(n_771),
.B(n_809),
.Y(n_1082)
);

AOI222xp33_ASAP7_75t_L g1083 ( 
.A1(n_991),
.A2(n_744),
.B1(n_742),
.B2(n_351),
.C1(n_355),
.C2(n_347),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_900),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_933),
.B(n_956),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_931),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_991),
.B(n_820),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_986),
.B(n_726),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_726),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_945),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_911),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_961),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_891),
.A2(n_374),
.B1(n_339),
.B2(n_347),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_894),
.B(n_351),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_894),
.B(n_355),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_911),
.B(n_365),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_891),
.A2(n_1053),
.B1(n_1014),
.B2(n_1002),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_968),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_960),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_885),
.A2(n_823),
.B(n_808),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_882),
.B(n_365),
.Y(n_1101)
);

AND2x6_ASAP7_75t_SL g1102 ( 
.A(n_998),
.B(n_1065),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1061),
.A2(n_823),
.B(n_828),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1015),
.A2(n_828),
.B(n_329),
.C(n_350),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_879),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1002),
.B(n_726),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_998),
.B(n_373),
.C(n_344),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_934),
.B(n_520),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_913),
.B(n_521),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_982),
.B(n_520),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_981),
.A2(n_354),
.B1(n_368),
.B2(n_340),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1014),
.A2(n_343),
.B(n_367),
.C(n_344),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_971),
.B(n_520),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_972),
.B(n_524),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_878),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_883),
.A2(n_918),
.B(n_921),
.C(n_1033),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_927),
.A2(n_343),
.B(n_371),
.C(n_348),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1009),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_931),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_879),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_884),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_936),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1023),
.A2(n_527),
.B(n_523),
.C(n_520),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1065),
.A2(n_373),
.B1(n_371),
.B2(n_370),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_915),
.B(n_362),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1053),
.A2(n_898),
.B1(n_1047),
.B2(n_888),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_976),
.B(n_1050),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_879),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1013),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1047),
.B(n_362),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_913),
.B(n_912),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_893),
.A2(n_527),
.B(n_523),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_915),
.B(n_12),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_996),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_959),
.A2(n_908),
.B(n_1058),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_951),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_981),
.A2(n_527),
.B(n_523),
.C(n_512),
.Y(n_1137)
);

NAND2x1_ASAP7_75t_L g1138 ( 
.A(n_887),
.B(n_890),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1063),
.B(n_523),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_887),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_895),
.A2(n_527),
.B(n_510),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_903),
.A2(n_512),
.B(n_510),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1063),
.B(n_528),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_909),
.A2(n_512),
.B(n_510),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_946),
.B(n_528),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_912),
.B(n_354),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_949),
.B(n_512),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_880),
.A2(n_528),
.B1(n_525),
.B2(n_512),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1063),
.B(n_525),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_927),
.A2(n_510),
.B(n_498),
.C(n_496),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1008),
.A2(n_1062),
.B(n_930),
.C(n_1005),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1022),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_973),
.Y(n_1153)
);

NOR2x1_ASAP7_75t_L g1154 ( 
.A(n_949),
.B(n_510),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1026),
.A2(n_354),
.B(n_528),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_887),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_953),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_930),
.B(n_950),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_944),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_897),
.A2(n_510),
.B(n_498),
.C(n_496),
.Y(n_1160)
);

AO32x2_ASAP7_75t_L g1161 ( 
.A1(n_1027),
.A2(n_13),
.A3(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1005),
.A2(n_498),
.B(n_496),
.C(n_22),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_950),
.A2(n_498),
.B(n_496),
.C(n_23),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_889),
.A2(n_489),
.B(n_498),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1031),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1063),
.B(n_528),
.Y(n_1166)
);

CKINVDCx8_ASAP7_75t_R g1167 ( 
.A(n_904),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_923),
.A2(n_489),
.B(n_498),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_926),
.B(n_354),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_946),
.B(n_20),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_994),
.B(n_528),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_955),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_910),
.A2(n_489),
.B(n_496),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_902),
.A2(n_496),
.B(n_528),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_944),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1056),
.B(n_528),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_887),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1029),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1042),
.B(n_528),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1037),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1054),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_957),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_925),
.A2(n_525),
.B(n_141),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_973),
.B(n_354),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_964),
.B(n_965),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_916),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_926),
.B(n_25),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_890),
.B(n_354),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1055),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_969),
.B(n_525),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_970),
.B(n_525),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1040),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1192)
);

BUFx4f_ASAP7_75t_SL g1193 ( 
.A(n_1036),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1057),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_925),
.A2(n_525),
.B(n_183),
.Y(n_1195)
);

AND2x2_ASAP7_75t_SL g1196 ( 
.A(n_1011),
.B(n_26),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_917),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_948),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_1198)
);

AOI33xp33_ASAP7_75t_L g1199 ( 
.A1(n_1011),
.A2(n_31),
.A3(n_32),
.B1(n_36),
.B2(n_37),
.B3(n_38),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_924),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1048),
.B(n_36),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1064),
.B(n_37),
.C(n_39),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_944),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_987),
.B(n_42),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1034),
.A2(n_1039),
.B(n_1001),
.C(n_937),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_944),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_929),
.A2(n_525),
.B(n_85),
.Y(n_1207)
);

BUFx4f_ASAP7_75t_L g1208 ( 
.A(n_986),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_914),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_966),
.A2(n_525),
.B(n_77),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_899),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_995),
.A2(n_525),
.B(n_96),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_954),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_986),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_890),
.B(n_76),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1043),
.B(n_44),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_890),
.B(n_104),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_986),
.B(n_107),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_954),
.B(n_920),
.Y(n_1219)
);

OAI22x1_ASAP7_75t_L g1220 ( 
.A1(n_892),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1000),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1000),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1012),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_977),
.A2(n_110),
.B(n_177),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_954),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1113),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1071),
.A2(n_907),
.B(n_928),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1094),
.A2(n_1006),
.B1(n_901),
.B2(n_896),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1212),
.A2(n_979),
.B(n_1017),
.Y(n_1229)
);

AO32x2_ASAP7_75t_L g1230 ( 
.A1(n_1097),
.A2(n_1041),
.A3(n_1051),
.B1(n_943),
.B2(n_983),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1185),
.A2(n_907),
.B(n_892),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1131),
.B(n_920),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1158),
.B(n_939),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1095),
.A2(n_1030),
.B(n_1032),
.C(n_978),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1085),
.A2(n_1030),
.B(n_1032),
.C(n_978),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1068),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1119),
.Y(n_1237)
);

CKINVDCx8_ASAP7_75t_R g1238 ( 
.A(n_1072),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1185),
.A2(n_962),
.B(n_958),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1109),
.B(n_1070),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1126),
.A2(n_940),
.A3(n_992),
.B(n_990),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1196),
.A2(n_997),
.B1(n_1059),
.B2(n_941),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1126),
.A2(n_985),
.A3(n_1004),
.B(n_1007),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1082),
.A2(n_1028),
.B(n_1018),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1092),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1087),
.A2(n_939),
.B1(n_941),
.B2(n_1021),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1205),
.A2(n_1010),
.B(n_993),
.Y(n_1247)
);

AOI221x1_ASAP7_75t_L g1248 ( 
.A1(n_1212),
.A2(n_1024),
.B1(n_1035),
.B2(n_919),
.C(n_988),
.Y(n_1248)
);

CKINVDCx14_ASAP7_75t_R g1249 ( 
.A(n_1153),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_1060),
.A3(n_1049),
.B(n_1003),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1086),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1067),
.A2(n_952),
.B(n_980),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1090),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1101),
.B(n_1052),
.C(n_967),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1132),
.A2(n_980),
.B(n_1020),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1208),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1151),
.A2(n_967),
.B(n_938),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1208),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1073),
.A2(n_1016),
.B(n_1046),
.C(n_1045),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1091),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1171),
.A2(n_1044),
.B(n_974),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1113),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1186),
.B(n_1051),
.Y(n_1263)
);

AO22x2_ASAP7_75t_L g1264 ( 
.A1(n_1097),
.A2(n_1012),
.B1(n_1041),
.B2(n_59),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1135),
.A2(n_997),
.B(n_963),
.C(n_947),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1174),
.A2(n_947),
.B(n_997),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1074),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1211),
.A2(n_997),
.B1(n_56),
.B2(n_62),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1100),
.A2(n_118),
.B(n_167),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1106),
.A2(n_1108),
.B(n_1103),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1141),
.A2(n_108),
.B(n_163),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1136),
.B(n_55),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1109),
.B(n_180),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1214),
.A2(n_62),
.A3(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1216),
.B(n_63),
.C(n_70),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1200),
.A2(n_151),
.A3(n_153),
.B(n_161),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1114),
.B(n_1127),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1125),
.B(n_1096),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1116),
.A2(n_1197),
.B(n_1178),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1079),
.B(n_1080),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1075),
.A2(n_1164),
.B(n_1173),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1133),
.A2(n_1107),
.B(n_1187),
.C(n_1170),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1122),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1168),
.A2(n_1144),
.B(n_1142),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1066),
.B(n_1083),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1204),
.A2(n_1202),
.B(n_1184),
.C(n_1093),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1143),
.A2(n_1149),
.B(n_1166),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1157),
.A2(n_1182),
.B1(n_1172),
.B2(n_1098),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1163),
.A2(n_1209),
.B(n_1162),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1171),
.A2(n_1110),
.B(n_1179),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1093),
.A2(n_1124),
.B1(n_1111),
.B2(n_1201),
.C(n_1198),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1110),
.A2(n_1179),
.B(n_1176),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1206),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1118),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1130),
.A2(n_1169),
.B1(n_1146),
.B2(n_1099),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1160),
.A2(n_1176),
.B(n_1191),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1143),
.A2(n_1149),
.B(n_1166),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1089),
.A2(n_1117),
.B(n_1192),
.C(n_1112),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1190),
.A2(n_1191),
.B(n_1139),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1069),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1129),
.Y(n_1301)
);

AO32x2_ASAP7_75t_L g1302 ( 
.A1(n_1214),
.A2(n_1148),
.A3(n_1161),
.B1(n_1102),
.B2(n_1199),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1081),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1223),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1105),
.A2(n_1128),
.B(n_1207),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1152),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1134),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1105),
.A2(n_1128),
.B(n_1210),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1148),
.A2(n_1150),
.A3(n_1220),
.B(n_1224),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_SL g1311 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1188),
.C(n_1138),
.Y(n_1311)
);

AO32x2_ASAP7_75t_L g1312 ( 
.A1(n_1161),
.A2(n_1155),
.A3(n_1078),
.B1(n_1137),
.B2(n_1145),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1121),
.A2(n_1115),
.B(n_1189),
.C(n_1165),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1105),
.A2(n_1128),
.B(n_1225),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1161),
.A2(n_1088),
.B(n_1218),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1180),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1105),
.A2(n_1128),
.B(n_1225),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1193),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1181),
.A2(n_1194),
.B1(n_1222),
.B2(n_1221),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1225),
.A2(n_1078),
.B(n_1195),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1203),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1183),
.A2(n_1123),
.B(n_1213),
.C(n_1147),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1225),
.A2(n_1076),
.B(n_1155),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1218),
.B(n_1159),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1159),
.B(n_1175),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1219),
.A2(n_1175),
.B(n_1120),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1154),
.A2(n_1120),
.B(n_1140),
.C(n_1156),
.Y(n_1327)
);

CKINVDCx16_ASAP7_75t_R g1328 ( 
.A(n_1167),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1088),
.A2(n_1219),
.A3(n_1140),
.B(n_1156),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1088),
.A2(n_1120),
.B(n_1140),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1156),
.A2(n_1177),
.B(n_1088),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1177),
.A2(n_999),
.B1(n_891),
.B2(n_932),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1177),
.Y(n_1333)
);

AO32x2_ASAP7_75t_L g1334 ( 
.A1(n_1097),
.A2(n_1126),
.A3(n_1214),
.B1(n_1093),
.B2(n_712),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1087),
.B(n_999),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_L g1336 ( 
.A(n_1094),
.B(n_768),
.C(n_999),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1087),
.B(n_999),
.Y(n_1337)
);

AOI221x1_ASAP7_75t_L g1338 ( 
.A1(n_1126),
.A2(n_1212),
.B1(n_1097),
.B2(n_981),
.C(n_768),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1167),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1122),
.B(n_556),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1131),
.B(n_1109),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1158),
.B(n_862),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1068),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1092),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1208),
.B(n_1105),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1092),
.B(n_906),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1126),
.A2(n_1104),
.A3(n_1097),
.B(n_943),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1167),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1122),
.B(n_556),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1071),
.A2(n_975),
.B(n_750),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1126),
.A2(n_1104),
.A3(n_1097),
.B(n_943),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1151),
.A2(n_999),
.B(n_932),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1068),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1073),
.A2(n_883),
.B(n_932),
.C(n_1033),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1092),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1119),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1092),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1071),
.A2(n_975),
.B(n_750),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1094),
.A2(n_999),
.B(n_1095),
.C(n_768),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1071),
.A2(n_975),
.B(n_750),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1212),
.A2(n_1155),
.B(n_932),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1087),
.B(n_999),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1092),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1084),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1167),
.B(n_556),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1084),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1092),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1084),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1087),
.B(n_999),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1158),
.B(n_862),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1071),
.A2(n_975),
.B(n_750),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1082),
.A2(n_1025),
.B(n_1132),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1151),
.A2(n_999),
.B(n_932),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1087),
.B(n_999),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1082),
.A2(n_1025),
.B(n_1132),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1087),
.B(n_999),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1087),
.B(n_999),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1071),
.A2(n_975),
.B(n_750),
.Y(n_1378)
);

BUFx5_ASAP7_75t_L g1379 ( 
.A(n_1088),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1113),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_SL g1381 ( 
.A1(n_1073),
.A2(n_883),
.B(n_932),
.C(n_1033),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1087),
.B(n_886),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1072),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1113),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1212),
.A2(n_1082),
.B(n_1171),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1113),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1073),
.A2(n_883),
.B(n_932),
.C(n_1033),
.Y(n_1387)
);

INVx3_ASAP7_75t_SL g1388 ( 
.A(n_1072),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1126),
.A2(n_1104),
.A3(n_1097),
.B(n_943),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1340),
.Y(n_1390)
);

INVx6_ASAP7_75t_L g1391 ( 
.A(n_1293),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1339),
.Y(n_1392)
);

BUFx4_ASAP7_75t_SL g1393 ( 
.A(n_1318),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1336),
.A2(n_1268),
.B1(n_1275),
.B2(n_1369),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1278),
.A2(n_1285),
.B1(n_1291),
.B2(n_1342),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1370),
.A2(n_1279),
.B1(n_1382),
.B2(n_1277),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1348),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1383),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1236),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1333),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1343),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1345),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1356),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1264),
.A2(n_1373),
.B1(n_1352),
.B2(n_1377),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1264),
.A2(n_1376),
.B1(n_1337),
.B2(n_1335),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1359),
.A2(n_1282),
.B1(n_1374),
.B2(n_1362),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1267),
.B(n_1304),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1353),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1328),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1341),
.A2(n_1233),
.B1(n_1289),
.B2(n_1240),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_SL g1411 ( 
.A(n_1367),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1365),
.A2(n_1332),
.B1(n_1274),
.B2(n_1334),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_SL g1413 ( 
.A(n_1293),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1294),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1364),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1341),
.A2(n_1240),
.B1(n_1272),
.B2(n_1232),
.Y(n_1416)
);

BUFx10_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1366),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1238),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1388),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1346),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1242),
.A2(n_1295),
.B1(n_1288),
.B2(n_1251),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1346),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1273),
.A2(n_1249),
.B1(n_1283),
.B2(n_1232),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1349),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1338),
.A2(n_1248),
.B1(n_1267),
.B2(n_1368),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1280),
.A2(n_1273),
.B1(n_1308),
.B2(n_1254),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1274),
.A2(n_1334),
.B1(n_1229),
.B2(n_1257),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1330),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1280),
.A2(n_1300),
.B1(n_1228),
.B2(n_1305),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1274),
.A2(n_1334),
.B1(n_1229),
.B2(n_1286),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1301),
.A2(n_1307),
.B1(n_1316),
.B2(n_1237),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1260),
.A2(n_1303),
.B1(n_1324),
.B2(n_1386),
.Y(n_1433)
);

CKINVDCx11_ASAP7_75t_R g1434 ( 
.A(n_1245),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1344),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1357),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1226),
.A2(n_1380),
.B1(n_1386),
.B2(n_1262),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1302),
.A2(n_1315),
.B1(n_1361),
.B2(n_1387),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1226),
.A2(n_1262),
.B1(n_1384),
.B2(n_1380),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1321),
.Y(n_1440)
);

INVx6_ASAP7_75t_L g1441 ( 
.A(n_1325),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1256),
.Y(n_1442)
);

AO22x1_ASAP7_75t_L g1443 ( 
.A1(n_1258),
.A2(n_1355),
.B1(n_1363),
.B2(n_1384),
.Y(n_1443)
);

INVx3_ASAP7_75t_SL g1444 ( 
.A(n_1258),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1326),
.Y(n_1445)
);

BUFx8_ASAP7_75t_SL g1446 ( 
.A(n_1263),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1298),
.A2(n_1354),
.B1(n_1381),
.B2(n_1246),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_1276),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1319),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1313),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1379),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1361),
.A2(n_1269),
.B1(n_1231),
.B2(n_1247),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1302),
.A2(n_1290),
.B1(n_1299),
.B2(n_1292),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1302),
.A2(n_1270),
.B1(n_1296),
.B2(n_1378),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1296),
.A2(n_1297),
.B1(n_1252),
.B2(n_1239),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_1371),
.B1(n_1360),
.B2(n_1358),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1265),
.A2(n_1327),
.B1(n_1322),
.B2(n_1234),
.Y(n_1457)
);

BUFx12f_ASAP7_75t_L g1458 ( 
.A(n_1311),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1329),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1235),
.A2(n_1331),
.B1(n_1323),
.B2(n_1309),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1385),
.A2(n_1261),
.B1(n_1271),
.B2(n_1227),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1329),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1276),
.Y(n_1463)
);

BUFx2_ASAP7_75t_R g1464 ( 
.A(n_1379),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1379),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1379),
.Y(n_1466)
);

INVx6_ASAP7_75t_L g1467 ( 
.A(n_1314),
.Y(n_1467)
);

BUFx4_ASAP7_75t_SL g1468 ( 
.A(n_1317),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1306),
.A2(n_1320),
.B1(n_1259),
.B2(n_1385),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1347),
.A2(n_1389),
.B1(n_1351),
.B2(n_1281),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1261),
.A2(n_1351),
.B1(n_1347),
.B2(n_1389),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1266),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1284),
.A2(n_1255),
.B(n_1375),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1312),
.A2(n_1230),
.B1(n_1310),
.B2(n_1372),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1244),
.A2(n_1310),
.B1(n_1230),
.B2(n_1312),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1230),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1312),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1310),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1241),
.A2(n_991),
.B1(n_999),
.B2(n_1336),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1241),
.A2(n_991),
.B1(n_999),
.B2(n_1336),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1243),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1243),
.A2(n_1359),
.B1(n_991),
.B2(n_1282),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1250),
.Y(n_1484)
);

BUFx8_ASAP7_75t_SL g1485 ( 
.A(n_1250),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1339),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1383),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1253),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1333),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1236),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1253),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1293),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1293),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1253),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1340),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1278),
.A2(n_991),
.B1(n_972),
.B2(n_976),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1339),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1287),
.Y(n_1498)
);

BUFx8_ASAP7_75t_L g1499 ( 
.A(n_1293),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1339),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1293),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1293),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1340),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1293),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1278),
.A2(n_1196),
.B1(n_991),
.B2(n_529),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1293),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1382),
.B(n_1342),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1253),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1339),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1236),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1256),
.B(n_1225),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1359),
.A2(n_991),
.B1(n_1282),
.B2(n_1342),
.Y(n_1518)
);

CKINVDCx6p67_ASAP7_75t_R g1519 ( 
.A(n_1339),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1339),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1382),
.B(n_1342),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1345),
.Y(n_1522)
);

BUFx12f_ASAP7_75t_L g1523 ( 
.A(n_1339),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1359),
.A2(n_991),
.B1(n_1282),
.B2(n_1342),
.Y(n_1524)
);

BUFx10_ASAP7_75t_L g1525 ( 
.A(n_1383),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1278),
.A2(n_1196),
.B1(n_991),
.B2(n_529),
.Y(n_1526)
);

INVx5_ASAP7_75t_L g1527 ( 
.A(n_1256),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1253),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1336),
.A2(n_991),
.B1(n_999),
.B2(n_1278),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1336),
.A2(n_739),
.B1(n_1268),
.B2(n_529),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1459),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1429),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1462),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1403),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1473),
.A2(n_1460),
.B(n_1463),
.Y(n_1536)
);

AND2x6_ASAP7_75t_L g1537 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1441),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1441),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1399),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1469),
.A2(n_1455),
.B(n_1461),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1406),
.B(n_1518),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1403),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1429),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1484),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1431),
.B(n_1412),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1524),
.A2(n_1509),
.B1(n_1526),
.B2(n_1531),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1429),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1414),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1415),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1477),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1485),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1509),
.A2(n_1526),
.B1(n_1531),
.B2(n_1483),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1418),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1412),
.B(n_1428),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1428),
.B(n_1405),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1477),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1471),
.B(n_1477),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1461),
.A2(n_1452),
.B(n_1472),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1475),
.A2(n_1450),
.B(n_1404),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1390),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1458),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1430),
.A2(n_1481),
.B(n_1480),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1471),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1395),
.B(n_1512),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1448),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1425),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1426),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1441),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1495),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1449),
.A2(n_1396),
.B1(n_1528),
.B2(n_1502),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1426),
.Y(n_1575)
);

BUFx2_ASAP7_75t_SL g1576 ( 
.A(n_1413),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1448),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1478),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1470),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1470),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1451),
.B(n_1445),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1410),
.A2(n_1407),
.B(n_1439),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1521),
.B(n_1504),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1465),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1437),
.A2(n_1427),
.B(n_1416),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1453),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1422),
.A2(n_1514),
.B(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1474),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1488),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1474),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1421),
.A2(n_1423),
.B1(n_1489),
.B2(n_1400),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1486),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1491),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1401),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1494),
.Y(n_1595)
);

AO21x1_ASAP7_75t_L g1596 ( 
.A1(n_1394),
.A2(n_1454),
.B(n_1456),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1496),
.B(n_1408),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1454),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1405),
.B(n_1438),
.Y(n_1599)
);

AO31x2_ASAP7_75t_L g1600 ( 
.A1(n_1438),
.A2(n_1451),
.A3(n_1456),
.B(n_1440),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1419),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1433),
.B(n_1530),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1505),
.B(n_1507),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1490),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1467),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1508),
.A2(n_1513),
.B1(n_1511),
.B2(n_1424),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1467),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1467),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1394),
.B(n_1432),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1443),
.Y(n_1610)
);

AO21x1_ASAP7_75t_L g1611 ( 
.A1(n_1402),
.A2(n_1522),
.B(n_1517),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1527),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1466),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1468),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1464),
.A2(n_1527),
.B(n_1436),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_SL g1616 ( 
.A(n_1409),
.B(n_1435),
.C(n_1398),
.Y(n_1616)
);

NAND2x1_ASAP7_75t_L g1617 ( 
.A(n_1402),
.B(n_1522),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1442),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1442),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1400),
.A2(n_1489),
.B1(n_1487),
.B2(n_1516),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1444),
.A2(n_1413),
.B(n_1500),
.Y(n_1621)
);

AO21x2_ASAP7_75t_L g1622 ( 
.A1(n_1446),
.A2(n_1391),
.B(n_1510),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1400),
.B(n_1489),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1492),
.Y(n_1624)
);

NAND2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1400),
.B(n_1489),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1492),
.A2(n_1510),
.B(n_1506),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1501),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1501),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1501),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1417),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1503),
.Y(n_1631)
);

NAND2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1503),
.B(n_1510),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1392),
.B(n_1497),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1487),
.B(n_1417),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1493),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1493),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1499),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1499),
.A2(n_1411),
.B(n_1525),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1525),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1420),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1578),
.B(n_1519),
.Y(n_1641)
);

BUFx12f_ASAP7_75t_L g1642 ( 
.A(n_1592),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1578),
.B(n_1434),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1549),
.A2(n_1397),
.B1(n_1393),
.B2(n_1411),
.C(n_1515),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1546),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1555),
.A2(n_1393),
.B1(n_1520),
.B2(n_1523),
.C(n_1542),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1609),
.A2(n_1585),
.B(n_1574),
.C(n_1566),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1541),
.A2(n_1562),
.B(n_1571),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1584),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1547),
.B(n_1570),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1601),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1547),
.B(n_1573),
.Y(n_1653)
);

BUFx12f_ASAP7_75t_L g1654 ( 
.A(n_1633),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1560),
.A2(n_1606),
.B1(n_1548),
.B2(n_1599),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1597),
.B(n_1583),
.C(n_1603),
.D(n_1575),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_SL g1657 ( 
.A1(n_1599),
.A2(n_1603),
.B1(n_1560),
.B2(n_1602),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1586),
.B(n_1548),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1596),
.B(n_1560),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1589),
.B(n_1595),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1541),
.A2(n_1562),
.B(n_1596),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1585),
.A2(n_1566),
.B(n_1602),
.C(n_1582),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1614),
.B(n_1540),
.Y(n_1663)
);

AO32x2_ASAP7_75t_L g1664 ( 
.A1(n_1538),
.A2(n_1572),
.A3(n_1539),
.B1(n_1612),
.B2(n_1588),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1564),
.B(n_1558),
.C(n_1591),
.D(n_1610),
.Y(n_1666)
);

BUFx4f_ASAP7_75t_SL g1667 ( 
.A(n_1633),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1552),
.B(n_1556),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1610),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1581),
.A2(n_1608),
.B(n_1607),
.Y(n_1672)
);

BUFx2_ASAP7_75t_R g1673 ( 
.A(n_1622),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1582),
.A2(n_1587),
.B(n_1563),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1554),
.A2(n_1614),
.B1(n_1639),
.B2(n_1558),
.C(n_1535),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1557),
.B(n_1598),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1594),
.B(n_1616),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1543),
.B(n_1553),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1546),
.Y(n_1679)
);

AND2x2_ASAP7_75t_SL g1680 ( 
.A(n_1554),
.B(n_1615),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1533),
.B(n_1544),
.Y(n_1681)
);

AND2x2_ASAP7_75t_SL g1682 ( 
.A(n_1615),
.B(n_1621),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1620),
.A2(n_1639),
.B(n_1604),
.C(n_1608),
.Y(n_1683)
);

AO32x2_ASAP7_75t_L g1684 ( 
.A1(n_1612),
.A2(n_1588),
.A3(n_1590),
.B1(n_1557),
.B2(n_1559),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_SL g1685 ( 
.A1(n_1615),
.A2(n_1621),
.B(n_1622),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_SL g1686 ( 
.A1(n_1617),
.A2(n_1635),
.B(n_1640),
.C(n_1613),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1563),
.A2(n_1567),
.B(n_1536),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1618),
.B(n_1619),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_SL g1689 ( 
.A(n_1622),
.B(n_1577),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1567),
.B(n_1579),
.Y(n_1690)
);

AO32x2_ASAP7_75t_L g1691 ( 
.A1(n_1624),
.A2(n_1561),
.A3(n_1580),
.B1(n_1579),
.B2(n_1600),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1569),
.B(n_1577),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1625),
.A2(n_1640),
.B1(n_1565),
.B2(n_1621),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1625),
.A2(n_1640),
.B1(n_1576),
.B2(n_1605),
.C(n_1593),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1625),
.A2(n_1576),
.B1(n_1580),
.B2(n_1636),
.C(n_1637),
.Y(n_1695)
);

AND2x4_ASAP7_75t_SL g1696 ( 
.A(n_1671),
.B(n_1533),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1681),
.B(n_1550),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1649),
.B(n_1600),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1682),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1655),
.A2(n_1537),
.B1(n_1623),
.B2(n_1621),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1649),
.B(n_1600),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1691),
.B(n_1600),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1670),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1691),
.B(n_1600),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1645),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1651),
.B(n_1561),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1691),
.B(n_1600),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1647),
.A2(n_1537),
.B1(n_1623),
.B2(n_1633),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1645),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1661),
.B(n_1545),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1679),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1653),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1661),
.B(n_1687),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1679),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.B(n_1626),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1671),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1671),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1660),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1668),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1655),
.A2(n_1537),
.B1(n_1623),
.B2(n_1581),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1687),
.B(n_1532),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1664),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1664),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1664),
.B(n_1534),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1674),
.B(n_1534),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1688),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1690),
.B(n_1569),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1705),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1722),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1713),
.B(n_1654),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1703),
.B(n_1676),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1696),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1722),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1706),
.B(n_1690),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1703),
.B(n_1658),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1700),
.A2(n_1648),
.B(n_1662),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1706),
.B(n_1678),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1700),
.A2(n_1693),
.B(n_1686),
.C(n_1695),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1699),
.A2(n_1659),
.B1(n_1657),
.B2(n_1656),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1712),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1712),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1725),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1721),
.A2(n_1659),
.B(n_1657),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1715),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1713),
.B(n_1650),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1719),
.B(n_1680),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1684),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1725),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1715),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1717),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1696),
.B(n_1689),
.Y(n_1754)
);

INVx4_ASAP7_75t_SL g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1727),
.B(n_1684),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1710),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1727),
.B(n_1684),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1721),
.A2(n_1659),
.B1(n_1647),
.B2(n_1646),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1708),
.A2(n_1666),
.B1(n_1646),
.B2(n_1675),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1717),
.B(n_1692),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1711),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1702),
.A2(n_1667),
.B1(n_1675),
.B2(n_1695),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1728),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1697),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1711),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1710),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1708),
.A2(n_1673),
.B1(n_1667),
.B2(n_1694),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1765),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1677),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1738),
.A2(n_1714),
.B(n_1701),
.Y(n_1775)
);

NAND2x1_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1716),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1778)
);

AND2x2_ASAP7_75t_SL g1779 ( 
.A(n_1742),
.B(n_1702),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1765),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1765),
.Y(n_1781)
);

AND2x2_ASAP7_75t_SL g1782 ( 
.A(n_1760),
.B(n_1702),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1769),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1732),
.B(n_1737),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1757),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1755),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1755),
.B(n_1723),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1745),
.B(n_1717),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1757),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1770),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1745),
.B(n_1718),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1650),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1759),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1732),
.B(n_1724),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1759),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1770),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1769),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1729),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1729),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1756),
.B(n_1704),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1730),
.B(n_1724),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1737),
.B(n_1726),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1733),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1756),
.B(n_1704),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1730),
.B(n_1707),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1758),
.B(n_1707),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1801),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1794),
.B(n_1739),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1794),
.B(n_1739),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1761),
.Y(n_1815)
);

NAND4xp75_ASAP7_75t_L g1816 ( 
.A(n_1782),
.B(n_1738),
.C(n_1644),
.D(n_1760),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1801),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1793),
.Y(n_1819)
);

CKINVDCx16_ASAP7_75t_R g1820 ( 
.A(n_1773),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1797),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1801),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1793),
.B(n_1736),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1784),
.B(n_1761),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1804),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1784),
.B(n_1740),
.Y(n_1827)
);

NAND2x1_ASAP7_75t_L g1828 ( 
.A(n_1774),
.B(n_1753),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1802),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1802),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1802),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1806),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1805),
.B(n_1740),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1782),
.B(n_1762),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1775),
.B(n_1693),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1806),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1806),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1805),
.B(n_1735),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1786),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1786),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_R g1843 ( 
.A(n_1773),
.B(n_1623),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1786),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1785),
.B(n_1735),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1775),
.B(n_1768),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1775),
.B(n_1774),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1790),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1775),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1776),
.A2(n_1741),
.B(n_1771),
.C(n_1746),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1790),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1785),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1776),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1810),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1785),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1820),
.B(n_1779),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1816),
.B(n_1643),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1818),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1826),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1832),
.B(n_1795),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1822),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1848),
.B(n_1774),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1829),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1823),
.B(n_1795),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1816),
.B(n_1633),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1836),
.A2(n_1779),
.B1(n_1763),
.B2(n_1746),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1848),
.B(n_1777),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1835),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1827),
.B(n_1790),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1830),
.Y(n_1871)
);

NAND4xp25_ASAP7_75t_L g1872 ( 
.A(n_1851),
.B(n_1741),
.C(n_1644),
.D(n_1766),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1819),
.A2(n_1779),
.B1(n_1766),
.B2(n_1771),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1811),
.B(n_1777),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1831),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1811),
.B(n_1777),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1814),
.B(n_1778),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1827),
.B(n_1791),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1826),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1814),
.B(n_1778),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1817),
.B(n_1778),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1854),
.Y(n_1882)
);

NAND4xp25_ASAP7_75t_L g1883 ( 
.A(n_1843),
.B(n_1683),
.C(n_1663),
.D(n_1694),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1833),
.Y(n_1885)
);

XNOR2xp5_ASAP7_75t_L g1886 ( 
.A(n_1828),
.B(n_1652),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1817),
.B(n_1788),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1847),
.B(n_1788),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1837),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1837),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1872),
.A2(n_1779),
.B1(n_1850),
.B2(n_1821),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1867),
.A2(n_1853),
.B(n_1847),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1855),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1867),
.A2(n_1776),
.B1(n_1843),
.B2(n_1815),
.C(n_1825),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1859),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1869),
.B(n_1825),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1874),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1873),
.A2(n_1673),
.B1(n_1716),
.B2(n_1734),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1866),
.A2(n_1812),
.B1(n_1813),
.B2(n_1788),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1834),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1857),
.A2(n_1846),
.B1(n_1701),
.B2(n_1698),
.C1(n_1796),
.C2(n_1792),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1874),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1862),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1858),
.B(n_1815),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1877),
.B(n_1789),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1883),
.A2(n_1753),
.B1(n_1665),
.B2(n_1669),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1866),
.A2(n_1846),
.B1(n_1839),
.B2(n_1849),
.C(n_1852),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1864),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1858),
.A2(n_1683),
.B(n_1641),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1882),
.B(n_1789),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1874),
.B(n_1841),
.Y(n_1912)
);

AOI21xp33_ASAP7_75t_L g1913 ( 
.A1(n_1856),
.A2(n_1844),
.B(n_1842),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1886),
.B(n_1642),
.Y(n_1914)
);

OAI222xp33_ASAP7_75t_L g1915 ( 
.A1(n_1861),
.A2(n_1840),
.B1(n_1845),
.B2(n_1734),
.C1(n_1789),
.C2(n_1796),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1871),
.Y(n_1916)
);

OAI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1865),
.A2(n_1734),
.B1(n_1845),
.B2(n_1840),
.C(n_1748),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1894),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1893),
.A2(n_1891),
.B1(n_1890),
.B2(n_1860),
.C(n_1879),
.Y(n_1919)
);

OAI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1892),
.A2(n_1880),
.B(n_1889),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1892),
.A2(n_1876),
.B1(n_1881),
.B2(n_1887),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1908),
.A2(n_1889),
.B1(n_1891),
.B2(n_1890),
.C(n_1860),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1914),
.B(n_1876),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1914),
.B(n_1876),
.Y(n_1924)
);

AOI222xp33_ASAP7_75t_L g1925 ( 
.A1(n_1905),
.A2(n_1868),
.B1(n_1863),
.B2(n_1888),
.C1(n_1885),
.C2(n_1875),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1896),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1910),
.B(n_1881),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1904),
.Y(n_1928)
);

AND2x2_ASAP7_75t_SL g1929 ( 
.A(n_1897),
.B(n_1637),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1909),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1898),
.B(n_1879),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1916),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1912),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1903),
.B(n_1880),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1898),
.B(n_1901),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1912),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1912),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1911),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1937),
.B(n_1900),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1935),
.B(n_1906),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1920),
.A2(n_1907),
.B1(n_1899),
.B2(n_1895),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1923),
.B(n_1917),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1934),
.B(n_1881),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1931),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1938),
.B(n_1936),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1933),
.B(n_1907),
.Y(n_1946)
);

NAND5xp2_ASAP7_75t_L g1947 ( 
.A(n_1923),
.B(n_1902),
.C(n_1913),
.D(n_1863),
.E(n_1868),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1924),
.B(n_1915),
.Y(n_1948)
);

AOI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1947),
.A2(n_1919),
.B1(n_1921),
.B2(n_1922),
.C(n_1927),
.Y(n_1949)
);

NAND4xp25_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1924),
.C(n_1927),
.D(n_1925),
.Y(n_1950)
);

OAI31xp33_ASAP7_75t_L g1951 ( 
.A1(n_1948),
.A2(n_1933),
.A3(n_1932),
.B(n_1930),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1941),
.A2(n_1929),
.B1(n_1928),
.B2(n_1926),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1944),
.B(n_1918),
.C(n_1929),
.Y(n_1953)
);

OAI21xp33_ASAP7_75t_L g1954 ( 
.A1(n_1939),
.A2(n_1887),
.B(n_1878),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1940),
.B(n_1887),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1943),
.B(n_1870),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1946),
.A2(n_1638),
.B(n_1636),
.C(n_1884),
.Y(n_1957)
);

OAI211xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1949),
.A2(n_1945),
.B(n_1663),
.C(n_1791),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1953),
.Y(n_1959)
);

O2A1O1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1950),
.A2(n_1798),
.B(n_1804),
.C(n_1792),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_SL g1961 ( 
.A1(n_1954),
.A2(n_1798),
.B1(n_1799),
.B2(n_1796),
.C(n_1792),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1951),
.A2(n_1638),
.B(n_1798),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1959),
.A2(n_1952),
.B(n_1962),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1958),
.A2(n_1955),
.B1(n_1956),
.B2(n_1957),
.Y(n_1964)
);

AOI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1960),
.A2(n_1799),
.B1(n_1701),
.B2(n_1698),
.C(n_1752),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1961),
.A2(n_1754),
.B(n_1799),
.Y(n_1966)
);

AOI221x1_ASAP7_75t_L g1967 ( 
.A1(n_1958),
.A2(n_1752),
.B1(n_1744),
.B2(n_1743),
.C(n_1747),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1959),
.A2(n_1632),
.B1(n_1624),
.B2(n_1754),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1964),
.A2(n_1764),
.B1(n_1754),
.B2(n_1669),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1963),
.B(n_1808),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1967),
.Y(n_1971)
);

XOR2xp5_ASAP7_75t_L g1972 ( 
.A(n_1968),
.B(n_1627),
.Y(n_1972)
);

NAND4xp75_ASAP7_75t_L g1973 ( 
.A(n_1965),
.B(n_1750),
.C(n_1611),
.D(n_1626),
.Y(n_1973)
);

OAI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1969),
.A2(n_1966),
.B1(n_1632),
.B2(n_1630),
.C(n_1617),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1971),
.B(n_1669),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1970),
.A2(n_1631),
.B(n_1629),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1974),
.A2(n_1972),
.B1(n_1973),
.B2(n_1781),
.Y(n_1977)
);

OAI22x1_ASAP7_75t_L g1978 ( 
.A1(n_1977),
.A2(n_1975),
.B1(n_1976),
.B2(n_1632),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1978),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1978),
.B(n_1803),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1980),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1980),
.Y(n_1982)
);

AO21x2_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1979),
.B(n_1781),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1981),
.B1(n_1630),
.B2(n_1780),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1809),
.B(n_1807),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1985),
.Y(n_1986)
);

OAI221xp5_ASAP7_75t_R g1987 ( 
.A1(n_1986),
.A2(n_1800),
.B1(n_1783),
.B2(n_1780),
.C(n_1772),
.Y(n_1987)
);

AOI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1630),
.B(n_1613),
.C(n_1628),
.Y(n_1988)
);


endmodule