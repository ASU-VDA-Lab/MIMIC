module fake_jpeg_31686_n_219 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_40),
.B1(n_26),
.B2(n_22),
.Y(n_66)
);

BUFx2_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_43),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_13),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_6),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_16),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_88),
.B1(n_92),
.B2(n_27),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_80),
.B1(n_84),
.B2(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_74),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_19),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_23),
.B(n_34),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_83),
.Y(n_98)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_32),
.B1(n_35),
.B2(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_89),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_32),
.B1(n_33),
.B2(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_28),
.B1(n_33),
.B2(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_45),
.B1(n_47),
.B2(n_36),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_108),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_44),
.B1(n_46),
.B2(n_39),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_42),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_115),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_8),
.B1(n_27),
.B2(n_91),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_8),
.B1(n_27),
.B2(n_81),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_113),
.B(n_60),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_90),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_82),
.B1(n_76),
.B2(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_92),
.B(n_70),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_65),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_62),
.A2(n_79),
.B1(n_70),
.B2(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_146),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_122),
.B(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_61),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_140),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_118),
.C(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_101),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_146),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_168),
.B1(n_148),
.B2(n_127),
.C(n_134),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_124),
.C(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_149),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_166),
.B(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_116),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_169),
.B(n_133),
.Y(n_174)
);

AOI22x1_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_122),
.B1(n_96),
.B2(n_119),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_126),
.B1(n_142),
.B2(n_125),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_96),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_102),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_139),
.B(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_171),
.B1(n_179),
.B2(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_164),
.A2(n_133),
.B1(n_166),
.B2(n_162),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_174),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_183),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_144),
.B1(n_142),
.B2(n_127),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_172),
.B(n_177),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_150),
.B1(n_151),
.B2(n_169),
.C(n_157),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_158),
.C(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.C(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_167),
.C(n_165),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_193),
.B1(n_170),
.B2(n_178),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_152),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_174),
.C(n_180),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_173),
.C(n_175),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_192),
.B(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_195),
.B1(n_186),
.B2(n_175),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_208),
.B1(n_197),
.B2(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_194),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_197),
.Y(n_209)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_211),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_204),
.B(n_203),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_212),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_120),
.A3(n_136),
.B1(n_145),
.B2(n_159),
.C1(n_180),
.C2(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_136),
.C(n_145),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_217),
.B1(n_136),
.B2(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_214),
.Y(n_219)
);


endmodule