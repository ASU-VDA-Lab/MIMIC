module fake_jpeg_27840_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_15),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_52),
.Y(n_74)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_13),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_0),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_78),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_30),
.B1(n_22),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_67),
.B1(n_75),
.B2(n_3),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_23),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_73),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_89),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_27),
.B(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_22),
.B1(n_33),
.B2(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_50),
.B1(n_43),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_101),
.B1(n_90),
.B2(n_66),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_53),
.B1(n_47),
.B2(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_9),
.B1(n_10),
.B2(n_87),
.Y(n_139)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_108),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_46),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_102),
.B(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_47),
.B1(n_46),
.B2(n_3),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_12),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_110),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_110)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_12),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_118),
.Y(n_125)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_118),
.B1(n_99),
.B2(n_92),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_90),
.B1(n_67),
.B2(n_63),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_133),
.B1(n_138),
.B2(n_139),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_136),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_144),
.B(n_98),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_84),
.B1(n_80),
.B2(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_71),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_71),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_100),
.C(n_97),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

NOR2x1_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_100),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_163),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_101),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_156),
.B(n_161),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_93),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_112),
.B(n_98),
.C(n_97),
.D(n_115),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_164),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_109),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_145),
.B1(n_148),
.B2(n_140),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_138),
.B1(n_139),
.B2(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_123),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_150),
.C(n_172),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_145),
.B(n_132),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_123),
.B(n_127),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_155),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_158),
.C(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_186),
.C(n_180),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_154),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_204),
.Y(n_209)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_157),
.A3(n_152),
.B1(n_155),
.B2(n_159),
.C1(n_170),
.C2(n_166),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_162),
.B1(n_151),
.B2(n_153),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_178),
.B1(n_179),
.B2(n_192),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_213),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_182),
.B1(n_177),
.B2(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_218),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_219),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_189),
.B1(n_178),
.B2(n_186),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_189),
.A3(n_184),
.B1(n_176),
.B2(n_173),
.C1(n_180),
.C2(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_204),
.C(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_197),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_226),
.B1(n_214),
.B2(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_205),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_174),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_215),
.B1(n_216),
.B2(n_176),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_236),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_215),
.B1(n_135),
.B2(n_126),
.Y(n_234)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_223),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_217),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_236),
.Y(n_242)
);

AOI21x1_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_238),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_245),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_234),
.B(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_135),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_125),
.B(n_95),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_250),
.B(n_111),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_220),
.Y(n_253)
);


endmodule