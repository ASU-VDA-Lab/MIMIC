module fake_jpeg_19847_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_54),
.Y(n_61)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_42),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_15),
.B(n_30),
.C(n_29),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_34),
.B2(n_38),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_47),
.B1(n_22),
.B2(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_79),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_67),
.B(n_59),
.C(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_14),
.B1(n_28),
.B2(n_27),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_16),
.CI(n_25),
.CON(n_85),
.SN(n_85)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_3),
.C(n_4),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_4),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_72),
.B1(n_70),
.B2(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_84),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_92),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_96),
.C(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_83),
.B(n_91),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_85),
.Y(n_103)
);

OAI321xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_85),
.A3(n_89),
.B1(n_87),
.B2(n_6),
.C(n_7),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_11),
.B(n_12),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);


endmodule