module fake_jpeg_7373_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_26),
.B1(n_30),
.B2(n_41),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_41),
.B1(n_39),
.B2(n_20),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_83),
.B1(n_63),
.B2(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_65),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_70),
.B1(n_74),
.B2(n_19),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_69),
.Y(n_102)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_57),
.B1(n_48),
.B2(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_82),
.C(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_76),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_25),
.B1(n_29),
.B2(n_16),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_87),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_33),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_100),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_104),
.B1(n_19),
.B2(n_23),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_113),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

AND2x4_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_37),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_35),
.B(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_75),
.B1(n_76),
.B2(n_73),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_120),
.B(n_37),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_124),
.B(n_130),
.Y(n_154)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_126),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_113),
.B1(n_101),
.B2(n_94),
.Y(n_157)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_82),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_38),
.B1(n_35),
.B2(n_64),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_135),
.B1(n_142),
.B2(n_29),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_0),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_103),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_140),
.B(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_137),
.Y(n_158)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_31),
.B1(n_23),
.B2(n_90),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_75),
.C(n_59),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_147),
.C(n_36),
.Y(n_156)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_31),
.B1(n_90),
.B2(n_17),
.Y(n_142)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_44),
.C(n_37),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_92),
.B1(n_93),
.B2(n_106),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_149),
.A2(n_178),
.B1(n_71),
.B2(n_2),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_112),
.B(n_118),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_151),
.A2(n_152),
.B(n_164),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_25),
.B(n_16),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_159),
.C(n_163),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_56),
.C(n_55),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_113),
.B1(n_95),
.B2(n_32),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_161),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_95),
.B1(n_32),
.B2(n_27),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_136),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_21),
.B(n_32),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_27),
.B(n_24),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_165),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_22),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_37),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_27),
.B(n_24),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_145),
.B1(n_137),
.B2(n_126),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_51),
.B1(n_52),
.B2(n_22),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_180),
.B1(n_122),
.B2(n_138),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_179),
.Y(n_183)
);

NOR2x1_ASAP7_75t_R g192 ( 
.A(n_174),
.B(n_130),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_27),
.B1(n_24),
.B2(n_84),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_37),
.B1(n_24),
.B2(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_55),
.B1(n_71),
.B2(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_121),
.B1(n_148),
.B2(n_131),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_154),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_130),
.C(n_14),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_152),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_165),
.B(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_212),
.B1(n_150),
.B2(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_1),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_77),
.Y(n_202)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_77),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_207),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_9),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_151),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_216),
.C(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_156),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_150),
.B(n_171),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_195),
.B1(n_194),
.B2(n_188),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_154),
.CI(n_174),
.CON(n_222),
.SN(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_231),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_188),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_164),
.B1(n_155),
.B2(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

OR2x6_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_209),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_232),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_159),
.B(n_163),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_203),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_168),
.B1(n_71),
.B2(n_1),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_189),
.B1(n_184),
.B2(n_4),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_71),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_200),
.C(n_187),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_210),
.B1(n_208),
.B2(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_208),
.B1(n_210),
.B2(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_243),
.B(n_249),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_200),
.C(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_239),
.C(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_221),
.B1(n_217),
.B2(n_218),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_201),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_237),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_257),
.B1(n_237),
.B2(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_189),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_230),
.B1(n_216),
.B2(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_271),
.C(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_261),
.C(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_229),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_234),
.B(n_215),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_252),
.B(n_247),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_235),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_251),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_216),
.C(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_247),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_243),
.B(n_253),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_240),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_279),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_245),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_271),
.C(n_266),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_9),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_291),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_263),
.C(n_267),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_293),
.B(n_274),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_9),
.B(n_3),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_15),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_2),
.C(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_8),
.C(n_13),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_278),
.B1(n_10),
.B2(n_12),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_306),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_8),
.B(n_10),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_305),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_304),
.A3(n_301),
.B1(n_290),
.B2(n_298),
.C1(n_296),
.C2(n_288),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_309),
.B(n_312),
.C(n_313),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_317),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_295),
.B1(n_14),
.B2(n_15),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_13),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);

AOI221xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_295),
.B1(n_14),
.B2(n_15),
.C(n_13),
.Y(n_322)
);


endmodule