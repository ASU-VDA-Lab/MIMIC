module fake_netlist_6_3149_n_1626 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1626);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1626;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_1575;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_1380;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_1333;
wire n_1558;
wire n_699;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_619;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_645;
wire n_1381;
wire n_916;
wire n_608;
wire n_630;
wire n_792;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1075;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_928;
wire n_1214;
wire n_835;
wire n_850;
wire n_690;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_1339;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1220;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1223;
wire n_1286;
wire n_1053;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_914;
wire n_759;
wire n_1625;
wire n_1453;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1079;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_1407;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_833;
wire n_1567;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_652;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_1325;
wire n_1002;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1191;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_1028;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1450;
wire n_868;
wire n_859;
wire n_735;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1578;
wire n_1006;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_94),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_505),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_24),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_239),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_305),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_243),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_551),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_345),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_275),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_313),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_383),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_563),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_50),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_392),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_539),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_537),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_212),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_252),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_456),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_370),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_511),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_36),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_270),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_434),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_181),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_502),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_454),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_565),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_426),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_574),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_512),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_229),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_444),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_211),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_264),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_301),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_506),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_197),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_139),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_199),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_396),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_302),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_417),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_57),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_564),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_127),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_266),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_373),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_471),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_411),
.Y(n_634)
);

BUFx5_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_500),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_406),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_325),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_157),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_518),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_382),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_249),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_405),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_507),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_409),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_91),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_458),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_466),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_101),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_305),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_351),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_179),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_378),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_478),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_524),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_383),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_126),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_485),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_10),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_465),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_391),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_387),
.Y(n_663)
);

BUFx4f_ASAP7_75t_SL g664 ( 
.A(n_267),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_371),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_151),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_132),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_412),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_352),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_401),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_75),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_60),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_183),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_252),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_46),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_337),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_253),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_72),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_508),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_254),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_170),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_191),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_277),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_256),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_395),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_215),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_562),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_381),
.Y(n_688)
);

CKINVDCx16_ASAP7_75t_R g689 ( 
.A(n_251),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_513),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_90),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_158),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_573),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_545),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_250),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_528),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_331),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_318),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_498),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_404),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_346),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_194),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_149),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_159),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_355),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_365),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_397),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g708 ( 
.A(n_541),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_146),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_82),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_270),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_418),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_48),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_41),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_101),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_309),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_425),
.Y(n_717)
);

CKINVDCx14_ASAP7_75t_R g718 ( 
.A(n_245),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_481),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_376),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_152),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_398),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_297),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_372),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_107),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_141),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_212),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_255),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_566),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_570),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_366),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_363),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_66),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_561),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_523),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_150),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_350),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_448),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_399),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_569),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_169),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_94),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_455),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_529),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_248),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_567),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_472),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_217),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_420),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_374),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_153),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_510),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_390),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_287),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_400),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_390),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_216),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_380),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_42),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_560),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_558),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_242),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_415),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_138),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_95),
.Y(n_765)
);

BUFx5_ASAP7_75t_L g766 ( 
.A(n_542),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_496),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_200),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_393),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_401),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_46),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_344),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_385),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_394),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_5),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_553),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_304),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_277),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_388),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_575),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_83),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_306),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_451),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_416),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_375),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_389),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_286),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_527),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_473),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_533),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_384),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_530),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_501),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_324),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_319),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_487),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_461),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_97),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_503),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_370),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_317),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_379),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_176),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_142),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_403),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_216),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_201),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_186),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_196),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_149),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_198),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_556),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_267),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_240),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_338),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_540),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_269),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_371),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_288),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_460),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_443),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_433),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_298),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_21),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_81),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_328),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_407),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_185),
.Y(n_828)
);

BUFx2_ASAP7_75t_SL g829 ( 
.A(n_435),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_285),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_88),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_402),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_377),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_224),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_386),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_571),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_445),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_568),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_588),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_588),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_588),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_696),
.B(n_780),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_628),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_631),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_586),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_639),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_591),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_594),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_654),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_654),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_805),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_805),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_803),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_593),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_603),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_602),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_595),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_700),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_614),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_0),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_600),
.Y(n_861)
);

INVxp33_ASAP7_75t_SL g862 ( 
.A(n_579),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_598),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_605),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_718),
.B(n_2),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_608),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_757),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_689),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_585),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_635),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_609),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_610),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_743),
.B(n_2),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_592),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_612),
.Y(n_875)
);

CKINVDCx16_ASAP7_75t_R g876 ( 
.A(n_708),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_613),
.Y(n_877)
);

INVxp67_ASAP7_75t_SL g878 ( 
.A(n_648),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_635),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_584),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_607),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_635),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_635),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_840),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_841),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_843),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_855),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_868),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_855),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_880),
.Y(n_891)
);

XOR2xp5_ASAP7_75t_L g892 ( 
.A(n_848),
.B(n_620),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_876),
.B(n_607),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_845),
.B(n_719),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_844),
.Y(n_895)
);

AND2x6_ASAP7_75t_L g896 ( 
.A(n_870),
.B(n_611),
.Y(n_896)
);

BUFx8_ASAP7_75t_L g897 ( 
.A(n_881),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_846),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_847),
.B(n_735),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_857),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_849),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_863),
.B(n_767),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_850),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_851),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_852),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_842),
.A2(n_715),
.B1(n_619),
.B2(n_581),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

XOR2xp5_ASAP7_75t_L g908 ( 
.A(n_861),
.B(n_632),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_864),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_SL g910 ( 
.A(n_860),
.B(n_653),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_869),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_866),
.B(n_744),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_871),
.B(n_747),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_862),
.B(n_837),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_865),
.B(n_837),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_872),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_859),
.B(n_812),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_874),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_854),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_867),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_875),
.B(n_601),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_580),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_911),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_890),
.B(n_878),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_912),
.B(n_856),
.Y(n_925)
);

CKINVDCx8_ASAP7_75t_R g926 ( 
.A(n_900),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_887),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_913),
.B(n_877),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_887),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_916),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_919),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_918),
.B(n_611),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_894),
.B(n_873),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_909),
.B(n_690),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_917),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_899),
.B(n_879),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_902),
.B(n_915),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_914),
.B(n_853),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_893),
.B(n_645),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_891),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_889),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_885),
.A2(n_883),
.B(n_882),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_903),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_896),
.B(n_699),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_886),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_904),
.Y(n_946)
);

AND2x6_ASAP7_75t_L g947 ( 
.A(n_907),
.B(n_611),
.Y(n_947)
);

NOR2x1p5_ASAP7_75t_L g948 ( 
.A(n_920),
.B(n_582),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_906),
.B(n_587),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_896),
.B(n_746),
.Y(n_950)
);

AND2x6_ASAP7_75t_L g951 ( 
.A(n_884),
.B(n_668),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_910),
.B(n_717),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_895),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_897),
.B(n_734),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_898),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_901),
.B(n_761),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_905),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_892),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_908),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_908),
.Y(n_960)
);

AND2x2_ASAP7_75t_SL g961 ( 
.A(n_919),
.B(n_617),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_921),
.B(n_776),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_900),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_939),
.A2(n_789),
.B1(n_797),
.B2(n_784),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_942),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_949),
.A2(n_673),
.B1(n_698),
.B2(n_663),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_930),
.B(n_829),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_952),
.A2(n_748),
.B1(n_779),
.B2(n_728),
.Y(n_968)
);

AO22x2_ASAP7_75t_L g969 ( 
.A1(n_960),
.A2(n_806),
.B1(n_817),
.B2(n_802),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_L g970 ( 
.A1(n_938),
.A2(n_625),
.B(n_621),
.Y(n_970)
);

NAND2xp33_ASAP7_75t_L g971 ( 
.A(n_962),
.B(n_627),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_940),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_961),
.B(n_821),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_941),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_928),
.B(n_925),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_937),
.A2(n_633),
.B1(n_634),
.B2(n_629),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_953),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_927),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_957),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_926),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_936),
.A2(n_799),
.B1(n_738),
.B2(n_616),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_924),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_943),
.B(n_626),
.Y(n_983)
);

AO22x2_ASAP7_75t_L g984 ( 
.A1(n_959),
.A2(n_824),
.B1(n_678),
.B2(n_683),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_955),
.Y(n_985)
);

AO22x2_ASAP7_75t_L g986 ( 
.A1(n_958),
.A2(n_716),
.B1(n_725),
.B2(n_674),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_929),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_946),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_935),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_956),
.B(n_664),
.Y(n_990)
);

NOR2xp67_ASAP7_75t_L g991 ( 
.A(n_944),
.B(n_640),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_950),
.B(n_624),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_934),
.A2(n_835),
.B1(n_638),
.B2(n_652),
.C(n_651),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_922),
.B(n_583),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_945),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_946),
.B(n_636),
.Y(n_997)
);

AO22x2_ASAP7_75t_L g998 ( 
.A1(n_954),
.A2(n_705),
.B1(n_714),
.B2(n_692),
.Y(n_998)
);

NOR2x1_ASAP7_75t_L g999 ( 
.A(n_963),
.B(n_646),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_947),
.Y(n_1000)
);

OR2x2_ASAP7_75t_SL g1001 ( 
.A(n_947),
.B(n_622),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_932),
.B(n_661),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_932),
.A2(n_641),
.B1(n_655),
.B2(n_649),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_951),
.Y(n_1004)
);

OAI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_933),
.A2(n_665),
.B1(n_684),
.B2(n_670),
.C(n_660),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_L g1006 ( 
.A(n_933),
.B(n_656),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_942),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_942),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_931),
.B(n_637),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_926),
.Y(n_1010)
);

AO22x2_ASAP7_75t_L g1011 ( 
.A1(n_949),
.A2(n_685),
.B1(n_770),
.B2(n_739),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_931),
.B(n_686),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_942),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_934),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_942),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_923),
.Y(n_1016)
);

OAI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_933),
.A2(n_765),
.B1(n_768),
.B2(n_758),
.C(n_724),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_940),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_923),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_923),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_923),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_931),
.B(n_686),
.Y(n_1022)
);

AND2x6_ASAP7_75t_L g1023 ( 
.A(n_939),
.B(n_740),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_1014),
.B(n_659),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_982),
.B(n_783),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_1018),
.B(n_777),
.Y(n_1026)
);

AND2x2_ASAP7_75t_SL g1027 ( 
.A(n_964),
.B(n_1009),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_994),
.B(n_658),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_974),
.B(n_687),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1012),
.B(n_693),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_1022),
.B(n_694),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_788),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1023),
.B(n_790),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_1010),
.B(n_680),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_1016),
.B(n_712),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_816),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_973),
.B(n_729),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_990),
.B(n_995),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_996),
.B(n_730),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1006),
.B(n_820),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_977),
.B(n_749),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_979),
.B(n_752),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_976),
.B(n_760),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_991),
.B(n_763),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_972),
.B(n_985),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_989),
.B(n_793),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_1004),
.B(n_774),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_992),
.B(n_838),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_999),
.B(n_796),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_978),
.B(n_822),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_971),
.B(n_836),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_997),
.B(n_785),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_987),
.B(n_791),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_966),
.B(n_755),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_988),
.B(n_800),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_970),
.B(n_679),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1003),
.B(n_679),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_981),
.B(n_792),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_983),
.B(n_792),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1000),
.B(n_807),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1002),
.B(n_792),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_968),
.B(n_808),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_965),
.B(n_766),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_1007),
.B(n_809),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1008),
.B(n_766),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1013),
.B(n_814),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1011),
.B(n_786),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1015),
.B(n_828),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_SL g1070 ( 
.A(n_993),
.B(n_833),
.Y(n_1070)
);

NAND2xp33_ASAP7_75t_SL g1071 ( 
.A(n_998),
.B(n_589),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_1001),
.B(n_590),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_967),
.B(n_596),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_SL g1074 ( 
.A(n_967),
.B(n_597),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_984),
.B(n_818),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1005),
.B(n_819),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1017),
.B(n_599),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_986),
.B(n_604),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_969),
.B(n_606),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_975),
.B(n_615),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_994),
.B(n_618),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_975),
.B(n_623),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_SL g1083 ( 
.A(n_994),
.B(n_630),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_994),
.B(n_642),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_975),
.B(n_643),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_SL g1086 ( 
.A(n_994),
.B(n_644),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_975),
.B(n_647),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_975),
.B(n_650),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_975),
.B(n_657),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_994),
.B(n_662),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_975),
.B(n_666),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_975),
.B(n_667),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_975),
.B(n_669),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_975),
.B(n_671),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_975),
.B(n_672),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_975),
.B(n_675),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_975),
.B(n_676),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_L g1098 ( 
.A(n_1023),
.B(n_677),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_975),
.B(n_681),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_975),
.B(n_682),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_975),
.B(n_688),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_975),
.B(n_691),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_SL g1103 ( 
.A(n_994),
.B(n_697),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_975),
.B(n_701),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_SL g1105 ( 
.A(n_994),
.B(n_702),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_975),
.B(n_703),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_975),
.B(n_704),
.Y(n_1107)
);

XOR2xp5_ASAP7_75t_L g1108 ( 
.A(n_980),
.B(n_408),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_975),
.B(n_706),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1094),
.B(n_1100),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1027),
.A2(n_709),
.B1(n_710),
.B2(n_707),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1064),
.A2(n_723),
.B(n_720),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1101),
.B(n_711),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1066),
.A2(n_823),
.B(n_804),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1070),
.A2(n_834),
.B(n_832),
.C(n_713),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_1039),
.B(n_410),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1046),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_1065),
.A2(n_1),
.B(n_3),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1080),
.B(n_721),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1067),
.A2(n_726),
.B(n_727),
.C(n_722),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1034),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1061),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1036),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1069),
.A2(n_732),
.B1(n_733),
.B2(n_731),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1028),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1037),
.A2(n_414),
.B(n_413),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1082),
.B(n_736),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_1038),
.B(n_737),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1025),
.A2(n_421),
.B(n_419),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1041),
.A2(n_423),
.B(n_422),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1032),
.A2(n_427),
.A3(n_428),
.B(n_424),
.Y(n_1131)
);

AND2x6_ASAP7_75t_L g1132 ( 
.A(n_1075),
.B(n_429),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1109),
.A2(n_742),
.B(n_745),
.C(n_741),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_SL g1134 ( 
.A(n_1030),
.B(n_753),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1033),
.A2(n_431),
.A3(n_432),
.B(n_430),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1085),
.B(n_750),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1087),
.B(n_751),
.Y(n_1137)
);

INVx8_ASAP7_75t_L g1138 ( 
.A(n_1026),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1049),
.A2(n_437),
.B(n_436),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_1075),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1024),
.B(n_754),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1088),
.B(n_756),
.Y(n_1142)
);

AOI221x1_ASAP7_75t_L g1143 ( 
.A1(n_1063),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.C(n_7),
.Y(n_1143)
);

NAND3x1_ASAP7_75t_L g1144 ( 
.A(n_1068),
.B(n_762),
.C(n_759),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_1052),
.A2(n_439),
.B(n_438),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1089),
.B(n_764),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1079),
.A2(n_441),
.A3(n_442),
.B(n_440),
.Y(n_1147)
);

BUFx10_ASAP7_75t_L g1148 ( 
.A(n_1076),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1076),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1051),
.A2(n_447),
.B(n_446),
.Y(n_1150)
);

AO31x2_ASAP7_75t_L g1151 ( 
.A1(n_1058),
.A2(n_450),
.A3(n_452),
.B(n_449),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_SL g1152 ( 
.A(n_1055),
.B(n_830),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1071),
.A2(n_7),
.A3(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1091),
.A2(n_771),
.B1(n_772),
.B2(n_769),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1108),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_1053),
.B(n_775),
.C(n_773),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1092),
.B(n_778),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1093),
.A2(n_782),
.B1(n_787),
.B2(n_781),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1095),
.A2(n_795),
.B(n_794),
.Y(n_1159)
);

AO32x2_ASAP7_75t_L g1160 ( 
.A1(n_1048),
.A2(n_11),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1096),
.B(n_798),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1097),
.B(n_801),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1060),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_L g1164 ( 
.A(n_1107),
.B(n_815),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1042),
.A2(n_459),
.B(n_457),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1043),
.A2(n_463),
.B(n_462),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1106),
.A2(n_811),
.B1(n_813),
.B2(n_810),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1029),
.B(n_467),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1040),
.B(n_468),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1099),
.B(n_825),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1057),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1054),
.B(n_827),
.C(n_826),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1035),
.A2(n_470),
.B(n_469),
.Y(n_1173)
);

CKINVDCx14_ASAP7_75t_R g1174 ( 
.A(n_1073),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1102),
.B(n_831),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1098),
.A2(n_577),
.A3(n_578),
.B(n_576),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1112),
.A2(n_1062),
.B(n_1059),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_1110),
.A2(n_1044),
.B(n_1104),
.C(n_1050),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1138),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1113),
.B(n_1031),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1155),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1150),
.A2(n_1045),
.B(n_1047),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1117),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1117),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1123),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1140),
.Y(n_1186)
);

AO32x2_ASAP7_75t_L g1187 ( 
.A1(n_1154),
.A2(n_1056),
.A3(n_1078),
.B1(n_1072),
.B2(n_1074),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1170),
.A2(n_1077),
.B1(n_1083),
.B2(n_1081),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1122),
.A2(n_1121),
.B1(n_1172),
.B2(n_1149),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1165),
.A2(n_1086),
.B(n_1084),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1129),
.A2(n_1103),
.B(n_1090),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1152),
.A2(n_1105),
.B1(n_12),
.B2(n_9),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1166),
.A2(n_475),
.B(n_474),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1139),
.A2(n_477),
.B(n_476),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1173),
.A2(n_480),
.B(n_479),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1114),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1171),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1115),
.A2(n_483),
.B(n_482),
.Y(n_1198)
);

AOI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1124),
.A2(n_486),
.B1(n_488),
.B2(n_484),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1159),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1163),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1118),
.A2(n_490),
.A3(n_491),
.B(n_489),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1145),
.A2(n_493),
.B(n_492),
.Y(n_1203)
);

OR3x4_ASAP7_75t_SL g1204 ( 
.A(n_1144),
.B(n_15),
.C(n_16),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1175),
.B(n_17),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1126),
.A2(n_495),
.B(n_494),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1130),
.A2(n_499),
.B(n_497),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1119),
.A2(n_18),
.B(n_19),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1138),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1148),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1125),
.B(n_20),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1132),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1168),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1127),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1116),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_1174),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1153),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_1158),
.A2(n_30),
.A3(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1141),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1169),
.B(n_504),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1164),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1153),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1120),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1128),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_SL g1225 ( 
.A(n_1156),
.B(n_509),
.Y(n_1225)
);

OAI221xp5_ASAP7_75t_L g1226 ( 
.A1(n_1111),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1176),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1160),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1132),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1167),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1136),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1137),
.B(n_1142),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1161),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1157),
.A2(n_515),
.B(n_514),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1143),
.A2(n_517),
.B(n_516),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1147),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1133),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1134),
.B(n_43),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1131),
.A2(n_520),
.B(n_519),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1147),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1135),
.A2(n_522),
.B(n_521),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1135),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1110),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_1174),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1123),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1138),
.B(n_525),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_SL g1248 ( 
.A(n_1152),
.B(n_48),
.C(n_49),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1185),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1241),
.A2(n_532),
.B(n_531),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1246),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1201),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1179),
.B(n_1183),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1197),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1243),
.A2(n_535),
.B(n_534),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1237),
.A2(n_538),
.B(n_536),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1216),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1196),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1184),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1209),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_R g1261 ( 
.A(n_1181),
.B(n_1231),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1234),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1210),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1227),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1217),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1222),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1186),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1220),
.B(n_51),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1242),
.A2(n_544),
.B(n_543),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1245),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1228),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1247),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1213),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1218),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1207),
.A2(n_547),
.B(n_546),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1218),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1206),
.A2(n_549),
.B(n_548),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1212),
.B(n_550),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1205),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1187),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1236),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1244),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1238),
.Y(n_1283)
);

OAI222xp33_ASAP7_75t_L g1284 ( 
.A1(n_1226),
.A2(n_54),
.B1(n_56),
.B2(n_52),
.C1(n_53),
.C2(n_55),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1214),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1224),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1180),
.B(n_52),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1229),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_SL g1289 ( 
.A(n_1211),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1232),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1215),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1219),
.B(n_552),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1191),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1223),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1233),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1202),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1202),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1178),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1239),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1235),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1261),
.B(n_1248),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1272),
.B(n_1189),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1249),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_R g1304 ( 
.A(n_1257),
.B(n_1188),
.Y(n_1304)
);

XNOR2xp5_ASAP7_75t_L g1305 ( 
.A(n_1270),
.B(n_1192),
.Y(n_1305)
);

CKINVDCx8_ASAP7_75t_R g1306 ( 
.A(n_1263),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1286),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1290),
.B(n_1208),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1251),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1259),
.B(n_1190),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1279),
.B(n_1221),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1299),
.B(n_1198),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_R g1313 ( 
.A(n_1289),
.B(n_1288),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1252),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_R g1315 ( 
.A(n_1278),
.B(n_1253),
.Y(n_1315)
);

NAND2xp33_ASAP7_75t_R g1316 ( 
.A(n_1287),
.B(n_1177),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1254),
.B(n_1200),
.Y(n_1317)
);

NAND2xp33_ASAP7_75t_R g1318 ( 
.A(n_1268),
.B(n_1240),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_1267),
.B(n_1194),
.Y(n_1319)
);

OR2x4_ASAP7_75t_L g1320 ( 
.A(n_1292),
.B(n_1204),
.Y(n_1320)
);

XNOR2xp5_ASAP7_75t_L g1321 ( 
.A(n_1273),
.B(n_1199),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1260),
.B(n_1225),
.Y(n_1322)
);

NAND2xp33_ASAP7_75t_R g1323 ( 
.A(n_1269),
.B(n_1193),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1295),
.B(n_1230),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1265),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_R g1326 ( 
.A(n_1269),
.B(n_1195),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1258),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1266),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1285),
.B(n_1203),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1291),
.B(n_1182),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_R g1331 ( 
.A(n_1256),
.B(n_1280),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1303),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1313),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1309),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1325),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1301),
.B(n_1294),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_SL g1337 ( 
.A(n_1312),
.B(n_1329),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1314),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1327),
.B(n_1282),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1328),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1311),
.B(n_1283),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1310),
.B(n_1271),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1302),
.B(n_1298),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1330),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1317),
.B(n_1274),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1307),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1322),
.B(n_1262),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1324),
.B(n_1321),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1306),
.B(n_1284),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1331),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1319),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1320),
.B(n_1276),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_1296),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1305),
.B(n_1297),
.Y(n_1354)
);

NOR2x1_ASAP7_75t_L g1355 ( 
.A(n_1316),
.B(n_1255),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1318),
.B(n_1293),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1323),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1326),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1315),
.B(n_1281),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1308),
.B(n_1264),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1310),
.B(n_1300),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1333),
.Y(n_1362)
);

AND2x2_ASAP7_75t_SL g1363 ( 
.A(n_1351),
.B(n_1250),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1346),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1335),
.Y(n_1365)
);

AOI33xp33_ASAP7_75t_L g1366 ( 
.A1(n_1348),
.A2(n_56),
.A3(n_58),
.B1(n_53),
.B2(n_55),
.B3(n_57),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1334),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1338),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1358),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1342),
.B(n_1275),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1342),
.B(n_1277),
.Y(n_1371)
);

XNOR2xp5_ASAP7_75t_L g1372 ( 
.A(n_1354),
.B(n_59),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1357),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

OAI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1352),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_62),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1360),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1356),
.B(n_1345),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1359),
.B(n_63),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1337),
.B(n_64),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1341),
.B(n_65),
.Y(n_1380)
);

NOR2xp67_ASAP7_75t_L g1381 ( 
.A(n_1350),
.B(n_1344),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1361),
.B(n_66),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1361),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1347),
.Y(n_1384)
);

OAI31xp33_ASAP7_75t_L g1385 ( 
.A1(n_1353),
.A2(n_1343),
.A3(n_1355),
.B(n_69),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1336),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1349),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1339),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1340),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1332),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1336),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1340),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1340),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1362),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1373),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1377),
.B(n_77),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1376),
.B(n_78),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1367),
.Y(n_1399)
);

INVx3_ASAP7_75t_R g1400 ( 
.A(n_1378),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1388),
.B(n_79),
.Y(n_1401)
);

AND2x2_ASAP7_75t_SL g1402 ( 
.A(n_1366),
.B(n_79),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1390),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1383),
.B(n_80),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1393),
.B(n_1394),
.Y(n_1405)
);

NOR2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1379),
.B(n_80),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1381),
.B(n_81),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1368),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1391),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1382),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1370),
.B(n_84),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1371),
.B(n_1363),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1380),
.B(n_85),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1372),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1385),
.B(n_86),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1375),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_86),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1387),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1392),
.B(n_87),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1374),
.B(n_89),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1376),
.B(n_89),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1365),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1369),
.B(n_91),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1377),
.B(n_92),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1389),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1364),
.Y(n_1426)
);

NAND2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1384),
.B(n_554),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1377),
.B(n_93),
.Y(n_1428)
);

AO221x2_ASAP7_75t_L g1429 ( 
.A1(n_1416),
.A2(n_98),
.B1(n_100),
.B2(n_97),
.C(n_99),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1400),
.B(n_96),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_R g1431 ( 
.A(n_1402),
.B(n_100),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1415),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1426),
.Y(n_1433)
);

NAND2xp33_ASAP7_75t_SL g1434 ( 
.A(n_1406),
.B(n_106),
.Y(n_1434)
);

AO221x2_ASAP7_75t_L g1435 ( 
.A1(n_1401),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.C(n_111),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1418),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1405),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1417),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1412),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1414),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1410),
.Y(n_1441)
);

AO221x2_ASAP7_75t_L g1442 ( 
.A1(n_1398),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1407),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1403),
.B(n_124),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_125),
.Y(n_1445)
);

AO221x2_ASAP7_75t_L g1446 ( 
.A1(n_1421),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_1446)
);

NOR4xp25_ASAP7_75t_SL g1447 ( 
.A(n_1399),
.B(n_130),
.C(n_128),
.D(n_129),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1422),
.B(n_133),
.Y(n_1448)
);

OAI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1419),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1411),
.B(n_137),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1420),
.B(n_137),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1397),
.B(n_140),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1424),
.B(n_141),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1408),
.B(n_143),
.Y(n_1454)
);

NOR4xp25_ASAP7_75t_SL g1455 ( 
.A(n_1409),
.B(n_147),
.C(n_144),
.D(n_145),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1423),
.B(n_148),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1428),
.B(n_150),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1404),
.Y(n_1458)
);

AO221x2_ASAP7_75t_L g1459 ( 
.A1(n_1427),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.C(n_156),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1395),
.Y(n_1460)
);

AO221x2_ASAP7_75t_L g1461 ( 
.A1(n_1416),
.A2(n_162),
.B1(n_164),
.B2(n_161),
.C(n_163),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1425),
.B(n_160),
.Y(n_1462)
);

AO221x2_ASAP7_75t_L g1463 ( 
.A1(n_1416),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.C(n_168),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1396),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1425),
.B(n_171),
.Y(n_1465)
);

AO221x2_ASAP7_75t_L g1466 ( 
.A1(n_1416),
.A2(n_173),
.B1(n_175),
.B2(n_172),
.C(n_174),
.Y(n_1466)
);

AO221x2_ASAP7_75t_L g1467 ( 
.A1(n_1416),
.A2(n_179),
.B1(n_181),
.B2(n_178),
.C(n_180),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1416),
.A2(n_180),
.B1(n_177),
.B2(n_178),
.C(n_182),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_SL g1469 ( 
.A(n_1400),
.B(n_184),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1400),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1396),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1430),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1432),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1433),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1464),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1471),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1458),
.B(n_192),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1469),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_193),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1460),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1454),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1434),
.B(n_195),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1463),
.A2(n_1429),
.B1(n_1466),
.B2(n_1461),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1448),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1467),
.A2(n_1459),
.B1(n_1435),
.B2(n_1446),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1444),
.B(n_202),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_203),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1462),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1465),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_204),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1456),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1459),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1445),
.B(n_206),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1442),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_208),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1449),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1450),
.B(n_1439),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1436),
.A2(n_1438),
.B1(n_1440),
.B2(n_1468),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_213),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_214),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1470),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1443),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1464),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1443),
.B(n_218),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_L g1506 ( 
.A1(n_1431),
.A2(n_219),
.B(n_220),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1437),
.B(n_221),
.Y(n_1507)
);

AOI222xp33_ASAP7_75t_L g1508 ( 
.A1(n_1432),
.A2(n_224),
.B1(n_226),
.B2(n_222),
.C1(n_223),
.C2(n_225),
.Y(n_1508)
);

NAND3x1_ASAP7_75t_L g1509 ( 
.A(n_1452),
.B(n_225),
.C(n_227),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1437),
.B(n_228),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1437),
.B(n_230),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1470),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1470),
.B(n_232),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1494),
.B(n_234),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1509),
.A2(n_235),
.B(n_236),
.Y(n_1515)
);

OAI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1498),
.A2(n_1485),
.B1(n_1506),
.B2(n_1483),
.C(n_1478),
.Y(n_1516)
);

NAND2xp33_ASAP7_75t_L g1517 ( 
.A(n_1472),
.B(n_236),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1508),
.A2(n_238),
.B(n_237),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1502),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1503),
.B(n_241),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1513),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1496),
.C(n_1492),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_244),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1482),
.A2(n_246),
.B(n_247),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1476),
.Y(n_1526)
);

OAI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1512),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1488),
.B(n_260),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1501),
.Y(n_1530)
);

AOI32xp33_ASAP7_75t_L g1531 ( 
.A1(n_1497),
.A2(n_263),
.A3(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1489),
.B(n_261),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1481),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1484),
.B(n_265),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1474),
.B(n_268),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1477),
.B(n_271),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_L g1537 ( 
.A1(n_1500),
.A2(n_272),
.B(n_273),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1480),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1479),
.B(n_274),
.Y(n_1539)
);

AOI222xp33_ASAP7_75t_L g1540 ( 
.A1(n_1522),
.A2(n_1499),
.B1(n_1495),
.B2(n_1493),
.C1(n_1487),
.C2(n_1490),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1505),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1530),
.B(n_1486),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1519),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1516),
.A2(n_1507),
.B1(n_1511),
.B2(n_1510),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1538),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1524),
.B(n_276),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1517),
.A2(n_278),
.B(n_279),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1535),
.Y(n_1549)
);

NAND2x1_ASAP7_75t_L g1550 ( 
.A(n_1533),
.B(n_280),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1514),
.B(n_281),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_282),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1515),
.B(n_283),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_284),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1549),
.B(n_1531),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1545),
.B(n_1539),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1550),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1547),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1552),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1543),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1546),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1537),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1541),
.Y(n_1563)
);

INVxp33_ASAP7_75t_L g1564 ( 
.A(n_1542),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1544),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1554),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1553),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1548),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1551),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1562),
.B(n_1527),
.C(n_1518),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1564),
.A2(n_1525),
.B(n_1523),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1568),
.A2(n_1532),
.B(n_1529),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1555),
.B(n_285),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_SL g1575 ( 
.A(n_1565),
.B(n_289),
.C(n_290),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1556),
.B(n_291),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1558),
.B(n_292),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1567),
.A2(n_293),
.B(n_294),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_SL g1579 ( 
.A(n_1563),
.B(n_295),
.C(n_296),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1561),
.B(n_298),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1559),
.B(n_299),
.C(n_300),
.Y(n_1581)
);

NOR2xp67_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_303),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1569),
.A2(n_307),
.B(n_308),
.Y(n_1583)
);

OAI211xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1566),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1579),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1582),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1571),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1570),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_323),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1571),
.Y(n_1589)
);

O2A1O1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1575),
.A2(n_329),
.B(n_326),
.C(n_327),
.Y(n_1590)
);

AOI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1578),
.A2(n_330),
.B(n_331),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1574),
.B(n_330),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1576),
.B(n_332),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1573),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1572),
.B(n_333),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1583),
.A2(n_341),
.B1(n_343),
.B2(n_339),
.C1(n_340),
.C2(n_342),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1577),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1580),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1581),
.B(n_346),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1584),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1589),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1587),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1586),
.Y(n_1603)
);

NOR3xp33_ASAP7_75t_L g1604 ( 
.A(n_1595),
.B(n_351),
.C(n_353),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1597),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1597),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1598),
.B(n_1597),
.Y(n_1607)
);

NOR2x1_ASAP7_75t_L g1608 ( 
.A(n_1588),
.B(n_354),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1602),
.B(n_1594),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_R g1610 ( 
.A(n_1607),
.B(n_1593),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_R g1611 ( 
.A(n_1601),
.B(n_1591),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_R g1612 ( 
.A(n_1605),
.B(n_1599),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1603),
.B(n_1592),
.Y(n_1613)
);

NAND2x1_ASAP7_75t_SL g1614 ( 
.A(n_1608),
.B(n_1585),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1606),
.B(n_1590),
.Y(n_1615)
);

INVxp33_ASAP7_75t_SL g1616 ( 
.A(n_1610),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1616),
.A2(n_1609),
.B(n_1615),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1613),
.B(n_1614),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1618),
.A2(n_1611),
.B1(n_1612),
.B2(n_1604),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1619),
.A2(n_1596),
.B1(n_1600),
.B2(n_358),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1619),
.B(n_356),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1620),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1621),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1622),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1623),
.B1(n_365),
.B2(n_362),
.C(n_364),
.Y(n_1625)
);

AOI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_1626)
);


endmodule