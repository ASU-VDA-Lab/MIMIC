module fake_jpeg_749_n_226 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_36),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_44),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_60),
.Y(n_83)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_18),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_67),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_35),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_96),
.B1(n_107),
.B2(n_24),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_65),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_98),
.B1(n_20),
.B2(n_49),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_21),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_41),
.B1(n_59),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_28),
.B(n_27),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_125),
.B1(n_135),
.B2(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_18),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_115),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_136)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_63),
.B(n_65),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_80),
.B(n_102),
.C(n_69),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_15),
.B1(n_6),
.B2(n_8),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_5),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_132),
.Y(n_153)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_76),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_8),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_11),
.B1(n_15),
.B2(n_91),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_11),
.B1(n_77),
.B2(n_84),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_106),
.B1(n_90),
.B2(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_151),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_153),
.B(n_151),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_129),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_116),
.C(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_156),
.C(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_97),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_93),
.B(n_95),
.C(n_69),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_126),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_93),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_118),
.B1(n_131),
.B2(n_113),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_89),
.B1(n_117),
.B2(n_126),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_162),
.B1(n_152),
.B2(n_155),
.Y(n_179)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_114),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_167),
.C(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_158),
.B1(n_153),
.B2(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_140),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_143),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_128),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_139),
.B(n_153),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_153),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_188),
.B(n_174),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_166),
.B1(n_185),
.B2(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_141),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_138),
.C(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_174),
.C(n_171),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.C(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_168),
.C(n_175),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_159),
.B1(n_169),
.B2(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_146),
.C(n_157),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_146),
.C(n_169),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_184),
.C(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_196),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_200),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_195),
.C(n_207),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_211),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.C(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_208),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_218),
.B1(n_212),
.B2(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_207),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_179),
.B(n_183),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_137),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_225),
.Y(n_226)
);


endmodule