module real_jpeg_2392_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_33),
.B1(n_37),
.B2(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_27),
.C(n_28),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_23),
.B1(n_40),
.B2(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_28),
.B1(n_40),
.B2(n_50),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_3),
.B(n_49),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_58),
.C(n_62),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_3),
.B(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_76),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_37),
.C(n_77),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_64),
.Y(n_172)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_23),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_28),
.B1(n_38),
.B2(n_50),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_33),
.B1(n_37),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_128),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_210),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_189),
.B(n_209),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_108),
.B(n_131),
.C(n_132),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_17),
.B(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_68),
.B2(n_69),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_18),
.B(n_71),
.C(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_41),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_20),
.B(n_43),
.C(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_46),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_28),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_30),
.A2(n_31),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_31),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_31),
.B(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_31),
.B(n_130),
.C(n_172),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_32),
.B(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_33),
.A2(n_37),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_37),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_39),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_53),
.B2(n_67),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_42),
.A2(n_43),
.B1(n_90),
.B2(n_101),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_42),
.B(n_90),
.C(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_52),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_105),
.C(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_53),
.A2(n_67),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_53),
.A2(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_53),
.B(n_228),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_64),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_66),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_60),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22x1_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_62),
.B(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_88),
.B2(n_89),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_82),
.B2(n_83),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_72),
.A2(n_73),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_72),
.B(n_166),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_72),
.A2(n_73),
.B1(n_90),
.B2(n_101),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_72),
.B(n_90),
.C(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_75),
.B(n_80),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_74),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_76),
.A2(n_207),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_80),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_86),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_87),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_86),
.B(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.C(n_93),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_92),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_94),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_93),
.B(n_116),
.C(n_121),
.Y(n_192)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_95),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_104),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_106),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_133),
.C(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_114),
.C(n_123),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_125),
.B(n_129),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_127),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_130),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_129),
.A2(n_130),
.B1(n_144),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_139),
.C(n_144),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_151),
.B(n_188),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_138),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_182),
.B(n_187),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_176),
.B(n_181),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_168),
.B(n_175),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_162),
.B(n_167),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B(n_161),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_174),
.Y(n_175)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_186),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_191),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_194),
.C(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_208),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_208),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_233),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_232),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_226),
.B2(n_227),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);


endmodule