module fake_jpeg_20567_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_90),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_69),
.B(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_69),
.B1(n_57),
.B2(n_51),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_57),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_114),
.Y(n_135)
);

OA22x2_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_73),
.B1(n_55),
.B2(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_60),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_122),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_59),
.B1(n_48),
.B2(n_72),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_123),
.B1(n_109),
.B2(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_64),
.B1(n_71),
.B2(n_52),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_27),
.B(n_40),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_24),
.B(n_45),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_56),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_138),
.B(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_2),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_49),
.C(n_75),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_139),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_46),
.B1(n_68),
.B2(n_5),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_148),
.B1(n_136),
.B2(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_127),
.B1(n_8),
.B2(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_8),
.B1(n_13),
.B2(n_16),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_152),
.C(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_147),
.C(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_144),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_18),
.B(n_21),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_22),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_25),
.C(n_28),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_36),
.B(n_39),
.Y(n_165)
);


endmodule