module fake_jpeg_13864_n_496 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_496);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_496;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_59),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_60),
.B(n_110),
.Y(n_158)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_64),
.B(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_12),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_72),
.B(n_85),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_19),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_105),
.Y(n_131)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g172 ( 
.A(n_81),
.Y(n_172)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_12),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_31),
.A2(n_10),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_87),
.B(n_0),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_89),
.Y(n_154)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_46),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_36),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_44),
.B1(n_39),
.B2(n_47),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_31),
.B(n_8),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_108),
.Y(n_148)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_41),
.B(n_0),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_114),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_116),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_28),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_115),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_119),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_50),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_8),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_53),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_42),
.B1(n_23),
.B2(n_49),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_121),
.A2(n_133),
.B1(n_137),
.B2(n_174),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_43),
.B1(n_35),
.B2(n_56),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_166),
.B1(n_168),
.B2(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_49),
.B1(n_50),
.B2(n_27),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_35),
.B1(n_36),
.B2(n_27),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_131),
.Y(n_200)
);

NAND2xp67_ASAP7_75t_SL g218 ( 
.A(n_147),
.B(n_126),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_182),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_76),
.B(n_1),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_167),
.C(n_170),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_53),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_88),
.B(n_25),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_164),
.B(n_169),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_71),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_61),
.A2(n_46),
.B(n_3),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_68),
.A2(n_39),
.B1(n_57),
.B2(n_29),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_68),
.B(n_57),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_29),
.C(n_18),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_179),
.B1(n_181),
.B2(n_191),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_88),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_69),
.B1(n_67),
.B2(n_66),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_4),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_177),
.B(n_178),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_4),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_73),
.A2(n_6),
.B1(n_7),
.B2(n_46),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_74),
.A2(n_79),
.B1(n_95),
.B2(n_83),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_80),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_100),
.A2(n_109),
.B1(n_93),
.B2(n_92),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_123),
.B1(n_156),
.B2(n_126),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_91),
.A2(n_98),
.B1(n_99),
.B2(n_89),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_89),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_191),
.C(n_187),
.Y(n_225)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_196),
.B(n_197),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_143),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_199),
.B(n_200),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_143),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_205),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_186),
.B(n_146),
.C(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_207),
.B(n_217),
.Y(n_302)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_137),
.A2(n_193),
.B1(n_147),
.B2(n_162),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_210),
.A2(n_251),
.B1(n_231),
.B2(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_148),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_218),
.A2(n_252),
.B1(n_239),
.B2(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_221),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_130),
.B(n_176),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_231),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_227),
.Y(n_271)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_159),
.B(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_242),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_229),
.A2(n_214),
.B(n_218),
.C(n_225),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_163),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_188),
.C(n_183),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_237),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_235),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_183),
.A2(n_130),
.B1(n_139),
.B2(n_154),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_234),
.A2(n_255),
.B1(n_256),
.B2(n_259),
.Y(n_275)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_166),
.B(n_127),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_172),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_241),
.Y(n_292)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_149),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_244),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_139),
.B(n_172),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_151),
.B(n_124),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_247),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_151),
.B(n_173),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_124),
.B(n_128),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_248),
.B(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_208),
.Y(n_309)
);

BUFx16f_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_135),
.A2(n_153),
.B1(n_189),
.B2(n_184),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_152),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_153),
.A2(n_152),
.B1(n_157),
.B2(n_175),
.Y(n_256)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_157),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_175),
.B(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_198),
.Y(n_273)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_266),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_273),
.A2(n_290),
.B(n_288),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_204),
.A2(n_247),
.B1(n_209),
.B2(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_279),
.B1(n_289),
.B2(n_298),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_301),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_204),
.A2(n_209),
.B1(n_237),
.B2(n_228),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_198),
.A2(n_211),
.B1(n_202),
.B2(n_213),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_287),
.B1(n_205),
.B2(n_240),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_215),
.A2(n_219),
.B1(n_216),
.B2(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_200),
.B(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_299),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_253),
.B1(n_255),
.B2(n_212),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_197),
.B(n_206),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_250),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_223),
.B(n_226),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_270),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_207),
.B(n_230),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_268),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_195),
.B(n_227),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_273),
.A2(n_249),
.B1(n_222),
.B2(n_236),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_315),
.B1(n_319),
.B2(n_336),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_323),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_279),
.A2(n_245),
.B1(n_235),
.B2(n_254),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_317),
.A2(n_269),
.B1(n_281),
.B2(n_284),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_272),
.A2(n_203),
.B1(n_250),
.B2(n_296),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_289),
.B1(n_266),
.B2(n_308),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_337),
.B1(n_281),
.B2(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_263),
.B(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_325),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_265),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_263),
.B(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_282),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_334),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_290),
.B(n_271),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_338),
.B(n_327),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_285),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_266),
.C(n_293),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_335),
.C(n_342),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_303),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_299),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_266),
.A2(n_275),
.B1(n_304),
.B2(n_309),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_266),
.A2(n_298),
.B1(n_303),
.B2(n_270),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_274),
.Y(n_368)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_339),
.A2(n_340),
.B1(n_344),
.B2(n_332),
.Y(n_367)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_260),
.B(n_283),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_306),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_343),
.Y(n_363)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_301),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_345),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_269),
.A2(n_278),
.B1(n_285),
.B2(n_284),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_274),
.B1(n_291),
.B2(n_277),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_360),
.Y(n_386)
);

XOR2x2_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_305),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_314),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_368),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_356),
.A2(n_315),
.B1(n_314),
.B2(n_334),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_346),
.A2(n_294),
.B(n_281),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_357),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_346),
.A2(n_300),
.B(n_295),
.C(n_262),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_329),
.B(n_347),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_294),
.B(n_300),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_262),
.B(n_261),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_366),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_378),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_311),
.A2(n_277),
.B1(n_261),
.B2(n_286),
.Y(n_369)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_262),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_371),
.B(n_313),
.Y(n_402)
);

CKINVDCx9p33_ASAP7_75t_R g372 ( 
.A(n_312),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_372),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_261),
.C(n_286),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_319),
.C(n_324),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_286),
.B(n_337),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_402),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_393),
.B1(n_365),
.B2(n_363),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_335),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_385),
.C(n_389),
.Y(n_406)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_322),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_388),
.B(n_394),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_310),
.C(n_336),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_390),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_310),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_401),
.C(n_403),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_356),
.A2(n_317),
.B1(n_343),
.B2(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_370),
.B(n_325),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_398),
.Y(n_405)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_377),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_329),
.C(n_316),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_321),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_392),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_403),
.B(n_370),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_391),
.B(n_365),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_421),
.Y(n_438)
);

HAxp5_ASAP7_75t_SL g410 ( 
.A(n_395),
.B(n_372),
.CON(n_410),
.SN(n_410)
);

NOR3xp33_ASAP7_75t_SL g439 ( 
.A(n_410),
.B(n_387),
.C(n_364),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_412),
.B1(n_390),
.B2(n_359),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_393),
.A2(n_349),
.B1(n_363),
.B2(n_378),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_386),
.B1(n_396),
.B2(n_399),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_371),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_379),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_355),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_349),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_419),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_360),
.C(n_353),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_423),
.C(n_395),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_387),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_364),
.C(n_374),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_376),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_405),
.Y(n_428)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_428),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_386),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_429),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_385),
.C(n_358),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_432),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_417),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_440),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_437),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_SL g436 ( 
.A(n_425),
.B(n_368),
.C(n_396),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_436),
.B(n_411),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_425),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_352),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_352),
.C(n_368),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_415),
.C(n_408),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_415),
.Y(n_453)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_443),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_446),
.B(n_433),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_424),
.B1(n_421),
.B2(n_380),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_361),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_453),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_423),
.C(n_416),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_456),
.C(n_457),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_416),
.C(n_413),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_407),
.C(n_422),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_419),
.C(n_414),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_449),
.B(n_438),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_460),
.B(n_404),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_448),
.A2(n_431),
.B1(n_426),
.B2(n_429),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_463),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_427),
.B1(n_432),
.B2(n_422),
.Y(n_463)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_464),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_453),
.C(n_454),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_466),
.B(n_467),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_447),
.C(n_455),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_446),
.A2(n_439),
.B(n_357),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_468),
.A2(n_359),
.B(n_456),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_474),
.Y(n_481)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_340),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_409),
.B1(n_414),
.B2(n_380),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_477),
.B(n_409),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_466),
.Y(n_478)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_478),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_476),
.B(n_467),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_480),
.A2(n_483),
.B(n_465),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_472),
.Y(n_486)
);

A2O1A1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_465),
.B(n_435),
.C(n_459),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_485),
.A2(n_487),
.B(n_488),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_486),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_459),
.C(n_469),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_447),
.C(n_475),
.Y(n_488)
);

AOI322xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_479),
.A3(n_377),
.B1(n_375),
.B2(n_351),
.C1(n_326),
.C2(n_330),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_490),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_491),
.A2(n_348),
.B(n_344),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_492),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_493),
.Y(n_496)
);


endmodule