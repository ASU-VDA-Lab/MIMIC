module fake_jpeg_20708_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_20),
.A2(n_14),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_75),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_60),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_67),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_72),
.B(n_86),
.Y(n_108)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_74),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_12),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_0),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_85),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_90),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_23),
.B1(n_35),
.B2(n_17),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_97),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_17),
.B1(n_38),
.B2(n_28),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_23),
.B1(n_35),
.B2(n_17),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_123),
.B1(n_130),
.B2(n_138),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_35),
.B1(n_29),
.B2(n_43),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_44),
.A2(n_29),
.B1(n_24),
.B2(n_38),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_65),
.A2(n_27),
.B1(n_28),
.B2(n_19),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_27),
.B1(n_15),
.B2(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_129),
.Y(n_158)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_51),
.A2(n_19),
.B1(n_36),
.B2(n_32),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_33),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_66),
.A2(n_33),
.B1(n_41),
.B2(n_36),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_76),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_50),
.B(n_33),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_5),
.B(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_53),
.B1(n_63),
.B2(n_60),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_48),
.B1(n_45),
.B2(n_78),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_141),
.B1(n_143),
.B2(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_153),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_84),
.B1(n_78),
.B2(n_62),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_62),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_149),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_36),
.B1(n_32),
.B2(n_41),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_146),
.Y(n_200)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_145),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_36),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_151),
.Y(n_187)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_32),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_108),
.A2(n_68),
.B1(n_32),
.B2(n_40),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_152),
.A2(n_88),
.B1(n_107),
.B2(n_117),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_109),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_40),
.B1(n_2),
.B2(n_4),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_1),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_160),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_4),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_89),
.B1(n_131),
.B2(n_88),
.Y(n_207)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

OR2x2_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_4),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_169),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_106),
.B1(n_121),
.B2(n_167),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_91),
.B(n_7),
.Y(n_173)
);

CKINVDCx6p67_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_181),
.B1(n_105),
.B2(n_100),
.Y(n_204)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_91),
.B(n_8),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_8),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OR2x4_ASAP7_75t_L g180 ( 
.A(n_92),
.B(n_10),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_93),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_100),
.A2(n_10),
.B1(n_105),
.B2(n_113),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_103),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_89),
.B(n_114),
.C(n_113),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_103),
.C(n_102),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_93),
.B(n_94),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_205),
.B(n_145),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_142),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_131),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_196),
.B(n_186),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_121),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_207),
.B1(n_161),
.B2(n_148),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_136),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_156),
.B(n_95),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_141),
.B1(n_154),
.B2(n_162),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_174),
.B1(n_166),
.B2(n_168),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_218),
.B1(n_174),
.B2(n_157),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_154),
.A2(n_107),
.B1(n_135),
.B2(n_106),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_165),
.B(n_178),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_152),
.B(n_180),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_222),
.A2(n_224),
.B(n_228),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_221),
.B(n_212),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_146),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_231),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_144),
.B(n_176),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_247),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_185),
.B(n_153),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_232),
.A2(n_248),
.B(n_250),
.Y(n_280)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_251),
.B1(n_184),
.B2(n_189),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_155),
.Y(n_240)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_157),
.B1(n_163),
.B2(n_174),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_249),
.B1(n_199),
.B2(n_195),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_155),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_204),
.B1(n_191),
.B2(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_168),
.B(n_166),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_168),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_254),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_198),
.B(n_194),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_201),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_257),
.B(n_250),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_200),
.B(n_218),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_261),
.A2(n_278),
.B1(n_243),
.B2(n_227),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_191),
.B1(n_202),
.B2(n_192),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_271),
.B1(n_273),
.B2(n_246),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_200),
.B(n_220),
.C(n_206),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_270),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_187),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_277),
.C(n_253),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_224),
.A2(n_216),
.B(n_197),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_268),
.Y(n_305)
);

NAND2x1p5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_197),
.Y(n_269)
);

XNOR2x2_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_228),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_216),
.B(n_197),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_206),
.B1(n_199),
.B2(n_193),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_193),
.B(n_189),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_243),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

HB1xp67_ASAP7_75t_SL g284 ( 
.A(n_269),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_269),
.C(n_262),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_270),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_248),
.C(n_252),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_291),
.C(n_292),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_293),
.B1(n_303),
.B2(n_261),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_298),
.B(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_255),
.B(n_231),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_296),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_248),
.C(n_233),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_248),
.C(n_233),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_245),
.B1(n_240),
.B2(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_249),
.C(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.C(n_257),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_247),
.C(n_244),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_239),
.B1(n_241),
.B2(n_236),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_239),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_307),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_272),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_319),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_276),
.B1(n_271),
.B2(n_275),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_318),
.B1(n_287),
.B2(n_303),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_264),
.B(n_294),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_317),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_280),
.C(n_276),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_323),
.C(n_302),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_297),
.A2(n_258),
.B1(n_268),
.B2(n_273),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_290),
.A2(n_259),
.B1(n_265),
.B2(n_263),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_326),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_280),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_264),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_292),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_229),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_260),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_306),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_329),
.A2(n_343),
.B(n_344),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_336),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_331),
.A2(n_345),
.B1(n_322),
.B2(n_327),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_294),
.B1(n_299),
.B2(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_332),
.A2(n_346),
.B1(n_318),
.B2(n_311),
.Y(n_348)
);

BUFx12_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_289),
.A3(n_283),
.B1(n_305),
.B2(n_296),
.C1(n_295),
.C2(n_288),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_324),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_236),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_298),
.C(n_256),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_314),
.C(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

INVx13_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_260),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_348),
.B(n_349),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_331),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_353),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_316),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_323),
.B1(n_307),
.B2(n_313),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_335),
.B1(n_338),
.B2(n_343),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_317),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_358),
.B(n_298),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_313),
.C(n_256),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_336),
.C(n_341),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_357),
.A2(n_329),
.B(n_335),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_362),
.A2(n_369),
.B1(n_370),
.B2(n_352),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_363),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_364),
.B(n_371),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_359),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_366),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_356),
.B(n_332),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_360),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_367),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_355),
.A2(n_344),
.B(n_334),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_362),
.A2(n_354),
.B(n_350),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_374),
.A2(n_358),
.B1(n_368),
.B2(n_345),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_353),
.B(n_334),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_L g381 ( 
.A1(n_378),
.A2(n_370),
.B(n_347),
.Y(n_381)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_334),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_368),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_369),
.A2(n_349),
.B1(n_345),
.B2(n_266),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_380),
.B(n_347),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_381),
.A2(n_383),
.B(n_385),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_382),
.B(n_377),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_373),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_376),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_387),
.A2(n_388),
.B(n_389),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_375),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_374),
.C(n_379),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_393),
.C(n_234),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_387),
.A2(n_384),
.B1(n_372),
.B2(n_266),
.Y(n_393)
);

AOI321xp33_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_272),
.A3(n_234),
.B1(n_237),
.B2(n_230),
.C(n_189),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_395),
.C(n_391),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_237),
.Y(n_397)
);


endmodule