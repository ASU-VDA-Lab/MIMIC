module fake_jpeg_10289_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_40),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_20),
.CON(n_62),
.SN(n_62)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_47),
.B1(n_27),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_30),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_34),
.B1(n_37),
.B2(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_22),
.B1(n_20),
.B2(n_33),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_38),
.B1(n_43),
.B2(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_32),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_18),
.B1(n_32),
.B2(n_26),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_38),
.B(n_27),
.C(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_78),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_26),
.Y(n_67)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_91),
.A3(n_68),
.B1(n_81),
.B2(n_85),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_26),
.A3(n_61),
.B1(n_30),
.B2(n_31),
.Y(n_105)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_43),
.B1(n_34),
.B2(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_66),
.B1(n_88),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_59),
.B1(n_46),
.B2(n_30),
.Y(n_119)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_43),
.B1(n_34),
.B2(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_51),
.B1(n_46),
.B2(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_89),
.B1(n_48),
.B2(n_45),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_40),
.C(n_42),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_42),
.C(n_37),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_56),
.B(n_47),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_18),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_75),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_121),
.B2(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_109),
.B(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_51),
.B1(n_89),
.B2(n_71),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_122),
.B(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_84),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_59),
.B1(n_46),
.B2(n_65),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_79),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_48),
.B1(n_23),
.B2(n_29),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_29),
.B1(n_19),
.B2(n_14),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_127),
.B1(n_137),
.B2(n_140),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_135),
.B1(n_107),
.B2(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_90),
.B1(n_80),
.B2(n_72),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_87),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_141),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_148),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_86),
.B1(n_83),
.B2(n_70),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_87),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_83),
.B1(n_29),
.B2(n_64),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_142),
.B1(n_154),
.B2(n_98),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_63),
.B1(n_37),
.B2(n_19),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_76),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_37),
.B1(n_13),
.B2(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_141),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_37),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_37),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_2),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_2),
.C(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_13),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_154)
);

BUFx12f_ASAP7_75t_SL g155 ( 
.A(n_144),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_158),
.B(n_164),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_161),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_109),
.B1(n_122),
.B2(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_167),
.B1(n_168),
.B2(n_125),
.Y(n_198)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_112),
.B1(n_104),
.B2(n_97),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_104),
.B(n_97),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_149),
.B(n_151),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_98),
.B1(n_99),
.B2(n_110),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_124),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_174),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_124),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_131),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_11),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_11),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_185)
);

OAI22x1_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_154),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_10),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_200),
.Y(n_234)
);

NAND2x1_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_145),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_212),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_214),
.B(n_185),
.C(n_186),
.Y(n_220)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_215),
.B1(n_159),
.B2(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_153),
.B1(n_150),
.B2(n_126),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_158),
.B1(n_177),
.B2(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_207),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_178),
.C(n_176),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_222),
.C(n_223),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_178),
.C(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_166),
.C(n_164),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_232),
.B1(n_235),
.B2(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_214),
.B1(n_201),
.B2(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_157),
.B1(n_163),
.B2(n_161),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_233),
.B1(n_202),
.B2(n_200),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_180),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_240),
.C(n_216),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_156),
.B1(n_174),
.B2(n_157),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_198),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_189),
.A2(n_170),
.B1(n_4),
.B2(n_5),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_196),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_6),
.C(n_7),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_244),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_203),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_253),
.C(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_233),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_196),
.B(n_205),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_227),
.B(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_212),
.C(n_209),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_259),
.A2(n_230),
.B(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_245),
.C(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_264),
.C(n_275),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_236),
.C(n_219),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_271),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_260),
.B(n_208),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_223),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_244),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_220),
.B(n_225),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_229),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_289),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_208),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_286),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_246),
.C(n_190),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_191),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_235),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_274),
.B1(n_250),
.B2(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_288),
.A2(n_240),
.B1(n_275),
.B2(n_208),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_236),
.B1(n_267),
.B2(n_276),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_12),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_261),
.B(n_263),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_199),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_296),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_284),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_191),
.B(n_199),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_289),
.C(n_269),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_305),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_6),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_293),
.Y(n_310)
);

AOI31xp67_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_290),
.A3(n_298),
.B(n_296),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_304),
.B(n_305),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_292),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_312),
.B(n_302),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_316),
.A3(n_314),
.B1(n_9),
.B2(n_8),
.C(n_7),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_8),
.B(n_9),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_9),
.Y(n_320)
);


endmodule