module fake_jpeg_11787_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_2),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_69),
.B1(n_52),
.B2(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_49),
.B1(n_63),
.B2(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_55),
.B1(n_66),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_49),
.B1(n_55),
.B2(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_87),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_48),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_67),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_63),
.C(n_5),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_84),
.B1(n_82),
.B2(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_105),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_112),
.B1(n_4),
.B2(n_10),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_113),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_58),
.B1(n_57),
.B2(n_56),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_11),
.B(n_12),
.Y(n_122)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_64),
.B1(n_7),
.B2(n_9),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_4),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_125),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_30),
.C(n_40),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_17),
.C(n_21),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_39),
.B1(n_28),
.B2(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_127),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_12),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_13),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_14),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_16),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.C(n_141),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_22),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_143),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_119),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_24),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_146),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_27),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_34),
.C(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_116),
.B(n_117),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_150),
.C(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_155),
.C(n_137),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_140),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_160),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_153),
.C(n_154),
.Y(n_163)
);

HAxp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_146),
.CON(n_164),
.SN(n_164)
);


endmodule