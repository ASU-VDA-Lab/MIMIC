module fake_jpeg_6152_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_36),
.C(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_57),
.B1(n_35),
.B2(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_60),
.B1(n_30),
.B2(n_20),
.Y(n_82)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_41),
.C(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_36),
.B1(n_33),
.B2(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_65),
.B1(n_74),
.B2(n_85),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_76),
.B(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_78),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_25),
.B1(n_41),
.B2(n_26),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_82),
.B1(n_45),
.B2(n_50),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_60),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_27),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_77),
.C(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_41),
.B1(n_20),
.B2(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_29),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_58),
.C(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_28),
.B1(n_31),
.B2(n_4),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_51),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_69),
.B1(n_76),
.B2(n_62),
.C(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_71),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_105),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_45),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_106),
.B1(n_46),
.B2(n_50),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_47),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_58),
.B1(n_55),
.B2(n_54),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_75),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_90),
.B(n_95),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_73),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_125),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_63),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_120),
.B(n_94),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_84),
.B(n_64),
.Y(n_118)
);

XNOR2x2_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_42),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_R g120 ( 
.A(n_91),
.B(n_83),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_78),
.B(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_130),
.B(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_127),
.B1(n_98),
.B2(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_81),
.B1(n_54),
.B2(n_46),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_42),
.B1(n_40),
.B2(n_54),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_108),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_75),
.B(n_40),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_40),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_102),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_42),
.B1(n_40),
.B2(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_93),
.B1(n_87),
.B2(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_144),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_90),
.B(n_88),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_134),
.C(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_113),
.B1(n_117),
.B2(n_135),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_1),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_127),
.B(n_118),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_3),
.B(n_4),
.Y(n_155)
);

AOI22x1_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_135),
.B1(n_114),
.B2(n_133),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_131),
.B1(n_124),
.B2(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_42),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_15),
.B1(n_14),
.B2(n_8),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_167),
.C(n_172),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_122),
.C(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_178),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_145),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_131),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_119),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_157),
.C(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_174),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_141),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_202),
.B(n_175),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_195),
.C(n_199),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_148),
.B1(n_150),
.B2(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_197),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_150),
.B1(n_176),
.B2(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_173),
.B1(n_183),
.B2(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_152),
.B(n_155),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_170),
.B(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_160),
.B1(n_136),
.B2(n_111),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_12),
.C(n_6),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_5),
.C(n_6),
.Y(n_211)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_216),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_166),
.C(n_8),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_224),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_190),
.B1(n_199),
.B2(n_185),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_188),
.C(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_193),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_192),
.B(n_214),
.Y(n_231)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_234),
.B(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_201),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_210),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_211),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_195),
.B(n_184),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_221),
.C(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.C(n_223),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_218),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_239),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_230),
.B(n_221),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_222),
.C(n_227),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_241),
.Y(n_251)
);

AOI321xp33_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_252),
.A3(n_249),
.B1(n_11),
.B2(n_12),
.C(n_10),
.Y(n_253)
);

OAI31xp33_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_5),
.A3(n_9),
.B(n_10),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_12),
.B(n_10),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_11),
.Y(n_255)
);


endmodule