module fake_jpeg_1549_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_56),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_41),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_53),
.B1(n_39),
.B2(n_38),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_52),
.B1(n_51),
.B2(n_58),
.Y(n_77)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_46),
.B1(n_40),
.B2(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_69),
.B1(n_52),
.B2(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_40),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_48),
.B1(n_39),
.B2(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_5),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_84),
.C(n_1),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_69),
.B(n_61),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_36),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_90),
.B1(n_98),
.B2(n_12),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_64),
.B1(n_66),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_101),
.B1(n_81),
.B2(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_95),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_49),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_1),
.B(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_11),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_10),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_9),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_35),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_112),
.B(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_113),
.B1(n_94),
.B2(n_14),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_10),
.Y(n_111)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_14),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_34),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_15),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_93),
.C(n_94),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_94),
.C(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_114),
.B1(n_18),
.B2(n_19),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_16),
.Y(n_130)
);

OAI322xp33_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_17),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_26),
.C2(n_27),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_108),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_117),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_138),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_125),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_133),
.C(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_122),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_129),
.B(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_139),
.C(n_123),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_29),
.B(n_30),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_31),
.Y(n_153)
);


endmodule