module real_aes_1726_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_0), .B(n_148), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_1), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_2), .A2(n_142), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_3), .B(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_4), .B(n_159), .Y(n_187) );
INVx1_ASAP7_75t_L g147 ( .A(n_5), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_6), .B(n_159), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_7), .B(n_183), .Y(n_556) );
INVx1_ASAP7_75t_L g473 ( .A(n_8), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_9), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_10), .Y(n_489) );
NAND2xp33_ASAP7_75t_L g259 ( .A(n_11), .B(n_157), .Y(n_259) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
AOI221x1_ASAP7_75t_L g141 ( .A1(n_13), .A2(n_25), .B1(n_142), .B2(n_148), .C(n_155), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_15), .B(n_148), .Y(n_255) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_16), .A2(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g564 ( .A(n_17), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_18), .B(n_137), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_19), .B(n_159), .Y(n_241) );
AO21x1_ASAP7_75t_L g181 ( .A1(n_20), .A2(n_148), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g119 ( .A(n_21), .Y(n_119) );
NOR2xp33_ASAP7_75t_SL g784 ( .A(n_21), .B(n_120), .Y(n_784) );
INVx1_ASAP7_75t_L g562 ( .A(n_22), .Y(n_562) );
INVx1_ASAP7_75t_SL g527 ( .A(n_23), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_24), .B(n_149), .Y(n_548) );
NAND2x1_ASAP7_75t_L g169 ( .A(n_26), .B(n_159), .Y(n_169) );
AOI33xp33_ASAP7_75t_L g501 ( .A1(n_27), .A2(n_54), .A3(n_455), .B1(n_460), .B2(n_502), .B3(n_503), .Y(n_501) );
NAND2x1_ASAP7_75t_L g215 ( .A(n_28), .B(n_157), .Y(n_215) );
INVx1_ASAP7_75t_L g482 ( .A(n_29), .Y(n_482) );
OR2x2_ASAP7_75t_L g140 ( .A(n_30), .B(n_87), .Y(n_140) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_30), .A2(n_87), .B(n_139), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_31), .B(n_463), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_32), .B(n_157), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_33), .A2(n_92), .B1(n_761), .B2(n_762), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_33), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_34), .B(n_159), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_35), .B(n_157), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_36), .A2(n_142), .B(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g143 ( .A(n_37), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g154 ( .A(n_37), .B(n_147), .Y(n_154) );
INVx1_ASAP7_75t_L g454 ( .A(n_37), .Y(n_454) );
OR2x6_ASAP7_75t_L g117 ( .A(n_38), .B(n_118), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g785 ( .A(n_38), .B(n_115), .C(n_786), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_39), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_40), .A2(n_51), .B1(n_775), .B2(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_40), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_41), .B(n_148), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_42), .B(n_463), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_43), .A2(n_174), .B1(n_183), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_44), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_45), .B(n_149), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_46), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_47), .B(n_157), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_48), .B(n_253), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_49), .B(n_149), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_50), .A2(n_142), .B(n_214), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_51), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_52), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_53), .B(n_157), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_55), .B(n_149), .Y(n_513) );
INVx1_ASAP7_75t_L g146 ( .A(n_56), .Y(n_146) );
INVx1_ASAP7_75t_L g151 ( .A(n_56), .Y(n_151) );
AND2x2_ASAP7_75t_L g514 ( .A(n_57), .B(n_137), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_58), .A2(n_75), .B1(n_452), .B2(n_463), .C(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_59), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_60), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_61), .B(n_174), .Y(n_491) );
AOI21xp5_ASAP7_75t_SL g451 ( .A1(n_62), .A2(n_452), .B(n_457), .Y(n_451) );
INVxp33_ASAP7_75t_L g789 ( .A(n_63), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_64), .A2(n_142), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g559 ( .A(n_65), .Y(n_559) );
AO21x1_ASAP7_75t_L g184 ( .A1(n_66), .A2(n_142), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_67), .B(n_148), .Y(n_205) );
INVx1_ASAP7_75t_L g512 ( .A(n_68), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_69), .B(n_148), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_70), .A2(n_452), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g198 ( .A(n_71), .B(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g144 ( .A(n_72), .Y(n_144) );
INVx1_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
AND2x2_ASAP7_75t_L g219 ( .A(n_73), .B(n_173), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_74), .B(n_463), .Y(n_504) );
AND2x2_ASAP7_75t_L g529 ( .A(n_76), .B(n_173), .Y(n_529) );
INVx1_ASAP7_75t_L g560 ( .A(n_77), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_78), .A2(n_452), .B(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_79), .A2(n_760), .B1(n_764), .B2(n_767), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_80), .A2(n_452), .B(n_496), .C(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
AND2x2_ASAP7_75t_L g203 ( .A(n_82), .B(n_173), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_83), .B(n_148), .Y(n_243) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_84), .B(n_173), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_85), .A2(n_452), .B1(n_499), .B2(n_500), .Y(n_498) );
AND2x2_ASAP7_75t_L g182 ( .A(n_86), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g176 ( .A(n_88), .B(n_173), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_89), .B(n_157), .Y(n_242) );
INVx1_ASAP7_75t_L g458 ( .A(n_90), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_91), .B(n_159), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_92), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_93), .B(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_94), .A2(n_142), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g505 ( .A(n_95), .B(n_173), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_96), .B(n_159), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_97), .A2(n_480), .B(n_481), .C(n_484), .Y(n_479) );
BUFx2_ASAP7_75t_L g107 ( .A(n_98), .Y(n_107) );
BUFx2_ASAP7_75t_SL g771 ( .A(n_98), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_99), .A2(n_142), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_100), .B(n_149), .Y(n_461) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_779), .B(n_788), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_122), .B(n_769), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_109), .A2(n_773), .B(n_778), .Y(n_772) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_121), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_113), .Y(n_778) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g128 ( .A(n_115), .B(n_117), .Y(n_128) );
OR2x6_ASAP7_75t_SL g439 ( .A(n_115), .B(n_116), .Y(n_439) );
OR2x2_ASAP7_75t_L g768 ( .A(n_115), .B(n_117), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_760), .B(n_763), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B1(n_437), .B2(n_440), .Y(n_124) );
CKINVDCx11_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
CKINVDCx6p67_ASAP7_75t_R g766 ( .A(n_126), .Y(n_766) );
INVx3_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_129), .A2(n_130), .B1(n_774), .B2(n_777), .Y(n_773) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_130), .A2(n_441), .B1(n_765), .B2(n_766), .Y(n_764) );
NAND4xp75_ASAP7_75t_L g130 ( .A(n_131), .B(n_347), .C(n_387), .D(n_416), .Y(n_130) );
NOR2x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_309), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_266), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_199), .B(n_220), .Y(n_133) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_162), .Y(n_134) );
AND2x4_ASAP7_75t_L g265 ( .A(n_135), .B(n_225), .Y(n_265) );
INVx1_ASAP7_75t_SL g318 ( .A(n_135), .Y(n_318) );
AOI21xp33_ASAP7_75t_L g353 ( .A1(n_135), .A2(n_354), .B(n_357), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_SL g357 ( .A1(n_135), .A2(n_358), .B(n_359), .C(n_360), .Y(n_357) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_135), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_135), .B(n_359), .Y(n_420) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g223 ( .A(n_136), .Y(n_223) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_136), .Y(n_297) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_161), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_137), .A2(n_205), .B(n_206), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_137), .Y(n_218) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_137), .A2(n_141), .B(n_161), .Y(n_307) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g183 ( .A(n_139), .B(n_140), .Y(n_183) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx3_ASAP7_75t_L g466 ( .A(n_143), .Y(n_466) );
AND2x6_ASAP7_75t_L g157 ( .A(n_144), .B(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g456 ( .A(n_144), .Y(n_456) );
AND2x4_ASAP7_75t_L g452 ( .A(n_145), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x4_ASAP7_75t_L g159 ( .A(n_146), .B(n_152), .Y(n_159) );
INVx2_ASAP7_75t_L g460 ( .A(n_146), .Y(n_460) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_147), .Y(n_465) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_154), .Y(n_148) );
INVx1_ASAP7_75t_L g483 ( .A(n_149), .Y(n_483) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx5_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_154), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_160), .Y(n_155) );
INVxp67_ASAP7_75t_L g563 ( .A(n_157), .Y(n_563) );
INVxp67_ASAP7_75t_L g565 ( .A(n_159), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_160), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_160), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_160), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_160), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_160), .A2(n_258), .B(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_160), .A2(n_458), .B(n_459), .C(n_461), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_160), .A2(n_459), .B(n_473), .C(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g499 ( .A(n_160), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_160), .A2(n_459), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g526 ( .A1(n_160), .A2(n_459), .B(n_527), .C(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_160), .A2(n_548), .B(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_160), .B(n_183), .Y(n_566) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_177), .Y(n_162) );
AND2x2_ASAP7_75t_L g289 ( .A(n_163), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g370 ( .A(n_163), .B(n_225), .Y(n_370) );
INVx1_ASAP7_75t_L g430 ( .A(n_163), .Y(n_430) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g274 ( .A(n_164), .B(n_190), .Y(n_274) );
AND2x2_ASAP7_75t_L g399 ( .A(n_164), .B(n_191), .Y(n_399) );
AND2x2_ASAP7_75t_L g404 ( .A(n_164), .B(n_364), .Y(n_404) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVxp67_ASAP7_75t_L g280 ( .A(n_165), .Y(n_280) );
BUFx3_ASAP7_75t_L g313 ( .A(n_165), .Y(n_313) );
AND2x2_ASAP7_75t_L g359 ( .A(n_165), .B(n_191), .Y(n_359) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_172), .B(n_176), .Y(n_165) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_166), .A2(n_172), .B(n_176), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B(n_198), .Y(n_191) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_172), .A2(n_192), .B(n_198), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_172), .A2(n_173), .B1(n_479), .B2(n_485), .Y(n_478) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_172), .A2(n_508), .B(n_514), .Y(n_507) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_172), .A2(n_508), .B(n_514), .Y(n_572) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_174), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
AND2x2_ASAP7_75t_L g344 ( .A(n_177), .B(n_222), .Y(n_344) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_190), .Y(n_177) );
AND2x4_ASAP7_75t_L g225 ( .A(n_178), .B(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g336 ( .A(n_178), .B(n_320), .Y(n_336) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_178), .B(n_307), .Y(n_379) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g315 ( .A(n_179), .Y(n_315) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g276 ( .A(n_180), .Y(n_276) );
OAI21x1_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_184), .B(n_188), .Y(n_180) );
INVx1_ASAP7_75t_L g189 ( .A(n_182), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_183), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_SL g237 ( .A(n_183), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_183), .A2(n_255), .B(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_183), .A2(n_451), .B(n_462), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_190), .B(n_276), .Y(n_279) );
AND2x2_ASAP7_75t_L g364 ( .A(n_190), .B(n_307), .Y(n_364) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g361 ( .A(n_191), .B(n_223), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_191), .B(n_307), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_193), .B(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_199), .B(n_270), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_199), .A2(n_393), .B1(n_394), .B2(n_395), .C(n_397), .Y(n_392) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI332xp33_ASAP7_75t_L g426 ( .A1(n_200), .A2(n_286), .A3(n_293), .B1(n_352), .B2(n_427), .B3(n_428), .C1(n_429), .C2(n_431), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_201), .B(n_210), .Y(n_200) );
AND2x2_ASAP7_75t_L g231 ( .A(n_201), .B(n_211), .Y(n_231) );
AND2x2_ASAP7_75t_L g248 ( .A(n_201), .B(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g261 ( .A(n_201), .Y(n_261) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_201), .B(n_262), .Y(n_321) );
INVx5_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2x1_ASAP7_75t_SL g283 ( .A(n_202), .B(n_249), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_202), .B(n_210), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_202), .B(n_211), .Y(n_294) );
BUFx2_ASAP7_75t_L g329 ( .A(n_202), .Y(n_329) );
AND2x2_ASAP7_75t_L g384 ( .A(n_202), .B(n_252), .Y(n_384) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
OR2x2_ASAP7_75t_L g251 ( .A(n_210), .B(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g262 ( .A(n_210), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g302 ( .A(n_210), .Y(n_302) );
AND2x2_ASAP7_75t_L g372 ( .A(n_210), .B(n_271), .Y(n_372) );
AND2x2_ASAP7_75t_L g385 ( .A(n_210), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_210), .B(n_386), .Y(n_403) );
INVx4_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_218), .A2(n_523), .B(n_529), .Y(n_522) );
OAI32xp33_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_227), .A3(n_232), .B1(n_246), .B2(n_264), .Y(n_220) );
INVx2_ASAP7_75t_L g330 ( .A(n_221), .Y(n_330) );
OR2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g341 ( .A(n_222), .Y(n_341) );
BUFx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g275 ( .A(n_223), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g408 ( .A(n_223), .B(n_313), .Y(n_408) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g320 ( .A(n_226), .Y(n_320) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g308 ( .A(n_229), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_229), .B(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_SL g319 ( .A(n_230), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g396 ( .A(n_230), .Y(n_396) );
AND2x2_ASAP7_75t_L g414 ( .A(n_230), .B(n_276), .Y(n_414) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp67_ASAP7_75t_SL g358 ( .A(n_233), .B(n_287), .Y(n_358) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_234), .B(n_269), .Y(n_356) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g432 ( .A(n_235), .B(n_302), .Y(n_432) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
INVx2_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_237), .B(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_260), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_247), .B(n_306), .Y(n_391) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND3x2_ASAP7_75t_L g346 ( .A(n_248), .B(n_293), .C(n_302), .Y(n_346) );
AND2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_249), .B(n_252), .Y(n_327) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g281 ( .A(n_251), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
INVx1_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
BUFx3_ASAP7_75t_L g293 ( .A(n_252), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_252), .B(n_304), .Y(n_303) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_253), .A2(n_471), .B(n_475), .Y(n_470) );
INVx2_ASAP7_75t_SL g496 ( .A(n_253), .Y(n_496) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x4_ASAP7_75t_L g312 ( .A(n_261), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_261), .B(n_271), .Y(n_355) );
AND2x2_ASAP7_75t_L g311 ( .A(n_262), .B(n_286), .Y(n_311) );
INVx2_ASAP7_75t_L g338 ( .A(n_262), .Y(n_338) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AOI211xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_272), .B(n_277), .C(n_298), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_267), .A2(n_394), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_270), .B(n_329), .Y(n_328) );
AOI211xp5_ASAP7_75t_SL g348 ( .A1(n_270), .A2(n_349), .B(n_353), .C(n_362), .Y(n_348) );
AND2x2_ASAP7_75t_L g334 ( .A(n_271), .B(n_294), .Y(n_334) );
OR2x2_ASAP7_75t_L g337 ( .A(n_271), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_274), .B(n_379), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_275), .B(n_320), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_275), .A2(n_301), .B1(n_381), .B2(n_384), .C(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g306 ( .A(n_276), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g352 ( .A(n_276), .B(n_307), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_281), .B1(n_284), .B2(n_288), .C(n_291), .Y(n_277) );
AND2x2_ASAP7_75t_L g423 ( .A(n_278), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g290 ( .A(n_279), .Y(n_290) );
INVx1_ASAP7_75t_L g376 ( .A(n_280), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_281), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g295 ( .A(n_283), .B(n_286), .Y(n_295) );
AND2x2_ASAP7_75t_L g371 ( .A(n_283), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_290), .B(n_297), .Y(n_296) );
OAI21xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_295), .B(n_296), .Y(n_291) );
INVx1_ASAP7_75t_L g415 ( .A(n_292), .Y(n_415) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g394 ( .A(n_293), .B(n_321), .Y(n_394) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_294), .B(n_303), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_305), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_333), .B1(n_336), .B2(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g405 ( .A(n_299), .Y(n_405) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
INVx1_ASAP7_75t_L g386 ( .A(n_304), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_306), .B(n_376), .Y(n_427) );
AND2x2_ASAP7_75t_L g395 ( .A(n_307), .B(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_308), .A2(n_389), .B(n_392), .C(n_400), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_331), .Y(n_309) );
AOI322xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .A3(n_314), .B1(n_316), .B2(n_321), .C1(n_322), .C2(n_330), .Y(n_310) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_312), .Y(n_428) );
AND2x2_ASAP7_75t_L g378 ( .A(n_313), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g412 ( .A(n_313), .Y(n_412) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_315), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_315), .B(n_361), .Y(n_369) );
AND2x2_ASAP7_75t_L g393 ( .A(n_315), .B(n_359), .Y(n_393) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g365 ( .A(n_319), .Y(n_365) );
NAND2xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_SL g368 ( .A1(n_324), .A2(n_369), .B1(n_370), .B2(n_371), .C(n_373), .Y(n_368) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g435 ( .A(n_327), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_335), .C(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g410 ( .A(n_334), .Y(n_410) );
INVx1_ASAP7_75t_L g342 ( .A(n_336), .Y(n_342) );
OR2x2_ASAP7_75t_L g429 ( .A(n_336), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g425 ( .A(n_337), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .B(n_345), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_341), .B(n_359), .Y(n_436) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_368), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_351), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
OR2x2_ASAP7_75t_L g402 ( .A(n_355), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI21xp33_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_365), .B(n_366), .Y(n_362) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AOI31xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .A3(n_380), .B(n_382), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_379), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B1(n_405), .B2(n_406), .C(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_413), .B2(n_415), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_426), .C(n_433), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_418), .B(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g765 ( .A(n_438), .Y(n_765) );
CKINVDCx11_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND3x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_650), .C(n_715), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_604), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_551), .B(n_577), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_515), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_467), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_447), .A2(n_652), .B(n_663), .Y(n_651) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_447), .B(n_593), .Y(n_686) );
AND2x2_ASAP7_75t_L g701 ( .A(n_447), .B(n_702), .Y(n_701) );
OR2x6_ASAP7_75t_L g711 ( .A(n_447), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_447), .B(n_703), .Y(n_713) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g587 ( .A(n_448), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_448), .B(n_601), .Y(n_600) );
INVx4_ASAP7_75t_L g619 ( .A(n_448), .Y(n_619) );
AND2x2_ASAP7_75t_L g622 ( .A(n_448), .B(n_540), .Y(n_622) );
NOR2x1_ASAP7_75t_SL g625 ( .A(n_448), .B(n_555), .Y(n_625) );
AND2x4_ASAP7_75t_L g637 ( .A(n_448), .B(n_635), .Y(n_637) );
OR2x2_ASAP7_75t_L g647 ( .A(n_448), .B(n_522), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_448), .B(n_659), .Y(n_664) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVxp67_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
NOR2x1p5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g503 ( .A(n_455), .Y(n_503) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x6_ASAP7_75t_L g459 ( .A(n_456), .B(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g480 ( .A(n_459), .Y(n_480) );
INVx2_ASAP7_75t_L g550 ( .A(n_459), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_459), .A2(n_483), .B1(n_559), .B2(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g464 ( .A(n_460), .B(n_465), .Y(n_464) );
INVxp33_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
INVx1_ASAP7_75t_L g492 ( .A(n_463), .Y(n_492) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_466), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_467), .A2(n_593), .B1(n_688), .B2(n_689), .Y(n_687) );
INVx1_ASAP7_75t_SL g731 ( .A(n_467), .Y(n_731) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_493), .Y(n_467) );
INVx2_ASAP7_75t_L g662 ( .A(n_468), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_468), .B(n_608), .Y(n_734) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_476), .Y(n_468) );
BUFx3_ASAP7_75t_L g580 ( .A(n_469), .Y(n_580) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g573 ( .A(n_470), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_470), .B(n_495), .Y(n_595) );
AND2x4_ASAP7_75t_L g612 ( .A(n_470), .B(n_613), .Y(n_612) );
INVxp67_ASAP7_75t_L g628 ( .A(n_470), .Y(n_628) );
INVx2_ASAP7_75t_L g685 ( .A(n_470), .Y(n_685) );
AND2x2_ASAP7_75t_L g603 ( .A(n_476), .B(n_569), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g649 ( .A(n_476), .B(n_572), .Y(n_649) );
AND2x2_ASAP7_75t_L g668 ( .A(n_476), .B(n_572), .Y(n_668) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g532 ( .A(n_477), .Y(n_532) );
INVx1_ASAP7_75t_L g611 ( .A(n_477), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_477), .B(n_507), .Y(n_630) );
AND2x4_ASAP7_75t_L g684 ( .A(n_477), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g643 ( .A(n_493), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_493), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
AND2x2_ASAP7_75t_L g627 ( .A(n_494), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g667 ( .A(n_494), .Y(n_667) );
AND2x2_ASAP7_75t_L g672 ( .A(n_494), .B(n_572), .Y(n_672) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_495), .B(n_507), .Y(n_534) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_505), .Y(n_495) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_496), .A2(n_497), .B(n_505), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_498), .B(n_504), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g608 ( .A(n_506), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_506), .B(n_580), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_506), .B(n_532), .Y(n_747) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_507), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
OAI21xp33_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_530), .B(n_535), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_518), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g585 ( .A(n_519), .Y(n_585) );
AND2x2_ASAP7_75t_L g599 ( .A(n_519), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g699 ( .A(n_519), .B(n_617), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_519), .B(n_746), .C(n_747), .Y(n_745) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_522), .B(n_555), .Y(n_598) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
AND2x2_ASAP7_75t_L g654 ( .A(n_522), .B(n_554), .Y(n_654) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_522), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_522), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g736 ( .A(n_530), .Y(n_736) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_531), .B(n_607), .Y(n_708) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g570 ( .A(n_532), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI211x1_ASAP7_75t_L g604 ( .A1(n_536), .A2(n_605), .B(n_614), .C(n_631), .Y(n_604) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_537), .B(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g657 ( .A(n_537), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g593 ( .A(n_539), .B(n_554), .Y(n_593) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g553 ( .A(n_540), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_540), .Y(n_618) );
INVx1_ASAP7_75t_L g635 ( .A(n_540), .Y(n_635) );
AND2x2_ASAP7_75t_L g703 ( .A(n_540), .B(n_555), .Y(n_703) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .C(n_545), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_567), .B(n_574), .Y(n_551) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_552), .B(n_619), .Y(n_722) );
INVx2_ASAP7_75t_L g754 ( .A(n_552), .Y(n_754) );
INVx4_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g586 ( .A(n_553), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g659 ( .A(n_554), .Y(n_659) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_566), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
OR2x2_ASAP7_75t_L g661 ( .A(n_568), .B(n_662), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g683 ( .A(n_568), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g583 ( .A(n_569), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g613 ( .A(n_569), .Y(n_613) );
INVx1_ASAP7_75t_L g737 ( .A(n_570), .Y(n_737) );
AND2x2_ASAP7_75t_L g602 ( .A(n_571), .B(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g584 ( .A(n_572), .Y(n_584) );
INVxp33_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g641 ( .A(n_576), .B(n_634), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_588), .C(n_596), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g665 ( .A(n_579), .B(n_666), .Y(n_665) );
NOR2xp67_ASAP7_75t_SL g670 ( .A(n_579), .B(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_580), .B(n_667), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_586), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
AND2x2_ASAP7_75t_L g714 ( .A(n_583), .B(n_684), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_586), .A2(n_733), .B1(n_735), .B2(n_738), .C1(n_739), .C2(n_742), .Y(n_732) );
INVx1_ASAP7_75t_L g696 ( .A(n_587), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_592), .Y(n_623) );
AND2x4_ASAP7_75t_SL g658 ( .A(n_592), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g712 ( .A(n_593), .Y(n_712) );
AND2x2_ASAP7_75t_L g757 ( .A(n_593), .B(n_609), .Y(n_757) );
AND2x2_ASAP7_75t_L g638 ( .A(n_594), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g751 ( .A(n_595), .B(n_630), .Y(n_751) );
OAI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_602), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_597), .A2(n_617), .B(n_658), .Y(n_718) );
AND2x2_ASAP7_75t_L g742 ( .A(n_598), .B(n_619), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g752 ( .A(n_598), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g690 ( .A(n_601), .Y(n_690) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_601), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g725 ( .A(n_603), .Y(n_725) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g728 ( .A(n_608), .B(n_612), .Y(n_728) );
BUFx2_ASAP7_75t_L g616 ( .A(n_609), .Y(n_616) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g639 ( .A(n_611), .Y(n_639) );
INVx2_ASAP7_75t_L g645 ( .A(n_611), .Y(n_645) );
AND2x2_ASAP7_75t_L g681 ( .A(n_611), .B(n_672), .Y(n_681) );
AND2x4_ASAP7_75t_L g648 ( .A(n_612), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g688 ( .A(n_612), .B(n_645), .Y(n_688) );
AND2x2_ASAP7_75t_L g739 ( .A(n_612), .B(n_740), .Y(n_739) );
AOI31xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_620), .A3(n_624), .B(n_626), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g636 ( .A(n_616), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x4_ASAP7_75t_L g634 ( .A(n_619), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_622), .A2(n_674), .B1(n_705), .B2(n_708), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_622), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g759 ( .A(n_622), .B(n_675), .Y(n_759) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g674 ( .A(n_625), .B(n_675), .Y(n_674) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
AND2x2_ASAP7_75t_L g697 ( .A(n_627), .B(n_668), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_629), .Y(n_707) );
INVx2_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_640), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g730 ( .A(n_633), .Y(n_730) );
AND2x2_ASAP7_75t_L g738 ( .A(n_634), .B(n_690), .Y(n_738) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_634), .Y(n_744) );
AND2x2_ASAP7_75t_L g689 ( .A(n_637), .B(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B1(n_646), .B2(n_648), .Y(n_640) );
NOR2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_643), .A2(n_662), .B1(n_756), .B2(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g655 ( .A(n_648), .Y(n_655) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_678), .Y(n_650) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OAI21xp33_ASAP7_75t_L g656 ( .A1(n_654), .A2(n_657), .B(n_660), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_657), .A2(n_681), .B1(n_682), .B2(n_686), .Y(n_680) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_669), .B2(n_673), .Y(n_663) );
INVx1_ASAP7_75t_L g698 ( .A(n_666), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g678 ( .A(n_679), .B(n_691), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_687), .Y(n_679) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
NAND2xp33_ASAP7_75t_SL g733 ( .A(n_683), .B(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g706 ( .A(n_684), .Y(n_706) );
INVx3_ASAP7_75t_L g720 ( .A(n_688), .Y(n_720) );
INVxp67_ASAP7_75t_L g749 ( .A(n_689), .Y(n_749) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_700), .C(n_704), .D(n_709), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_L g702 ( .A(n_694), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g750 ( .A(n_698), .Y(n_750) );
NAND2xp33_ASAP7_75t_SL g705 ( .A(n_706), .B(n_707), .Y(n_705) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B(n_714), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND3x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_732), .C(n_743), .Y(n_715) );
AOI221x1_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_721), .B2(n_723), .C(n_729), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_727), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_748), .C(n_755), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_748) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g777 ( .A(n_774), .Y(n_777) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
INVx3_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g791 ( .A(n_782), .Y(n_791) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_SL g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
endmodule