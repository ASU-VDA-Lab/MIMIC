module fake_jpeg_32054_n_293 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_52),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_2),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_26),
.B1(n_34),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_66),
.B1(n_67),
.B2(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_64),
.Y(n_93)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_38),
.B1(n_22),
.B2(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_26),
.B1(n_34),
.B2(n_22),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_38),
.B1(n_20),
.B2(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_23),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_29),
.C(n_38),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_70),
.C(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_36),
.B1(n_20),
.B2(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_75),
.B1(n_81),
.B2(n_86),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_36),
.B1(n_20),
.B2(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_46),
.B1(n_40),
.B2(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_36),
.B1(n_30),
.B2(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_37),
.B1(n_35),
.B2(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_24),
.B1(n_23),
.B2(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_27),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_33),
.C(n_30),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_124),
.C(n_5),
.Y(n_156)
);

NOR4xp25_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_103),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_107),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_109),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_37),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_32),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_33),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_32),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_18),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_18),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_17),
.Y(n_120)
);

INVxp33_ASAP7_75t_SL g122 ( 
.A(n_81),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_125),
.B1(n_59),
.B2(n_91),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_24),
.C(n_23),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_86),
.B1(n_79),
.B2(n_82),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_137),
.B1(n_140),
.B2(n_144),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_118),
.B1(n_97),
.B2(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_149),
.B1(n_121),
.B2(n_126),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_87),
.A3(n_74),
.B1(n_58),
.B2(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_135),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_113),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_127),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_79),
.B1(n_63),
.B2(n_59),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_16),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_14),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_93),
.A2(n_83),
.B1(n_65),
.B2(n_88),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_9),
.B(n_10),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_148),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_124),
.B1(n_111),
.B2(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_74),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_137),
.B1(n_128),
.B2(n_132),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_115),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_11),
.Y(n_183)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_8),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_95),
.C(n_106),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_167),
.C(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_172),
.B1(n_175),
.B2(n_179),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_164),
.B(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_95),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_126),
.C(n_117),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_178),
.B(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_113),
.B1(n_117),
.B2(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_113),
.B1(n_117),
.B2(n_13),
.Y(n_175)
);

AO21x1_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_113),
.B(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_10),
.B1(n_11),
.B2(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_11),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_132),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_135),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_156),
.B(n_154),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_168),
.B(n_182),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_179),
.C(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_144),
.C(n_140),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_202),
.C(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_136),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_131),
.C(n_152),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_151),
.C(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_141),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_138),
.B1(n_157),
.B2(n_172),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_213),
.B(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_162),
.B1(n_169),
.B2(n_166),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_229),
.B1(n_188),
.B2(n_190),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_174),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_228),
.C(n_210),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

FAx1_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_178),
.CI(n_183),
.CON(n_221),
.SN(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_188),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_231),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_194),
.C(n_203),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_166),
.B1(n_163),
.B2(n_180),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_210),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_205),
.B1(n_190),
.B2(n_197),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_198),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_240),
.B(n_221),
.C(n_215),
.D(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_236),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_229),
.B1(n_217),
.B2(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_232),
.B(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_206),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_199),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_226),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_256),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_257),
.B1(n_259),
.B2(n_225),
.Y(n_266)
);

BUFx12f_ASAP7_75t_SL g255 ( 
.A(n_245),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_260),
.B(n_243),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_234),
.C(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_215),
.C(n_233),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_238),
.B(n_240),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_233),
.B(n_237),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_269),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_221),
.C(n_232),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_248),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_251),
.B1(n_259),
.B2(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_262),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_250),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_264),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_282),
.C(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_263),
.C(n_214),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_258),
.B(n_254),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_277),
.B(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_274),
.C(n_276),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_279),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_284),
.B(n_224),
.Y(n_290)
);

AOI321xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_289),
.A3(n_253),
.B1(n_201),
.B2(n_195),
.C(n_204),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_195),
.B(n_191),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_191),
.Y(n_293)
);


endmodule