module fake_netlist_1_10079_n_658 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_658);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_13), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_60), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
OR2x2_ASAP7_75t_L g90 ( .A(n_76), .B(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_6), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_63), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_62), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_37), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_56), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_21), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_85), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_48), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_47), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_78), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_20), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_83), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_53), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_11), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_33), .B(n_79), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_23), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_75), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_32), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_34), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_36), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_35), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_55), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_49), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_50), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_41), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_82), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_22), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_58), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_92), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_99), .B(n_0), .Y(n_127) );
XOR2xp5_ASAP7_75t_L g128 ( .A(n_86), .B(n_0), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_100), .A2(n_108), .B1(n_104), .B2(n_91), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_87), .B(n_1), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_87), .B(n_1), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_116), .B(n_89), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_89), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_114), .B(n_2), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_98), .B(n_30), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_101), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_101), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_112), .A2(n_31), .B(n_81), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_91), .B(n_3), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_97), .B(n_4), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
NAND3x1_ASAP7_75t_L g156 ( .A(n_136), .B(n_97), .C(n_102), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_134), .B(n_111), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_132), .A2(n_102), .B1(n_105), .B2(n_124), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_132), .B(n_105), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_132), .B(n_113), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_140), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_134), .B(n_123), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_126), .B(n_94), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_126), .B(n_96), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_129), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
AND2x6_ASAP7_75t_L g172 ( .A(n_152), .B(n_122), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g173 ( .A(n_143), .B(n_90), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_152), .B(n_90), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_143), .B(n_115), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_138), .B(n_107), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_140), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_138), .B(n_103), .Y(n_179) );
INVx4_ASAP7_75t_SL g180 ( .A(n_143), .Y(n_180) );
CKINVDCx11_ASAP7_75t_R g181 ( .A(n_129), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_139), .B(n_122), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_143), .A2(n_120), .B1(n_117), .B2(n_113), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_139), .B(n_141), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_136), .A2(n_121), .B1(n_120), .B2(n_117), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_141), .B(n_118), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_175), .A2(n_127), .B1(n_147), .B2(n_149), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_175), .A2(n_127), .B1(n_147), .B2(n_149), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_154), .B(n_153), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_175), .B(n_153), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_159), .B(n_130), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_164), .B(n_145), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_169), .B(n_145), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_179), .B(n_144), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_157), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_183), .B(n_144), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_159), .B(n_130), .Y(n_206) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_172), .B(n_143), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_170), .B(n_128), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_162), .B(n_148), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_172), .B(n_121), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_189), .B(n_140), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_158), .A2(n_140), .B1(n_148), .B2(n_150), .Y(n_212) );
AND2x6_ASAP7_75t_SL g213 ( .A(n_181), .B(n_128), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_183), .B(n_148), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_159), .B(n_148), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_161), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_154), .B(n_109), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_177), .B(n_187), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_142), .B1(n_150), .B2(n_137), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_160), .B(n_150), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_160), .B(n_159), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_172), .A2(n_137), .B1(n_131), .B2(n_125), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
OAI22xp33_ASAP7_75t_SL g229 ( .A1(n_173), .A2(n_125), .B1(n_131), .B2(n_137), .Y(n_229) );
NOR2x1p5_ASAP7_75t_L g230 ( .A(n_156), .B(n_125), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_160), .B(n_131), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_172), .B(n_135), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_167), .B(n_135), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_167), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_174), .B(n_135), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_174), .B(n_135), .Y(n_236) );
NOR2xp33_ASAP7_75t_R g237 ( .A(n_210), .B(n_176), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_207), .A2(n_154), .B(n_182), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_199), .B(n_174), .Y(n_239) );
NOR2xp33_ASAP7_75t_R g240 ( .A(n_210), .B(n_174), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_203), .B(n_188), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_199), .B(n_186), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_154), .B(n_184), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_191), .Y(n_246) );
INVx4_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_194), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_196), .A2(n_184), .B(n_182), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_190), .A2(n_156), .B1(n_184), .B2(n_182), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_205), .B(n_180), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_200), .A2(n_184), .B(n_182), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_151), .B(n_163), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_166), .B(n_168), .C(n_171), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_199), .B(n_180), .Y(n_258) );
NOR2xp33_ASAP7_75t_R g259 ( .A(n_213), .B(n_5), .Y(n_259) );
AOI21x1_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_185), .B(n_171), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_193), .A2(n_133), .B1(n_135), .B2(n_106), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_195), .B(n_192), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_198), .A2(n_133), .B1(n_135), .B2(n_151), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_201), .A2(n_185), .B(n_168), .C(n_166), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_198), .A2(n_180), .B1(n_133), .B2(n_151), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_206), .A2(n_180), .B1(n_133), .B2(n_151), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_206), .B(n_133), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_211), .A2(n_163), .B(n_39), .C(n_84), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_192), .B(n_133), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_202), .A2(n_163), .B(n_165), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_206), .B(n_5), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_227), .B(n_165), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_204), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_6), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_221), .A2(n_165), .B(n_38), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_225), .A2(n_165), .B1(n_8), .B2(n_9), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_215), .B(n_7), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_SL g284 ( .A1(n_263), .A2(n_236), .B(n_235), .C(n_231), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_255), .A2(n_234), .B(n_228), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_243), .B(n_208), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_255), .A2(n_212), .B(n_224), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_260), .A2(n_234), .B(n_228), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_259), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_252), .A2(n_217), .B(n_209), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_260), .A2(n_218), .B(n_219), .Y(n_291) );
AO32x2_ASAP7_75t_L g292 ( .A1(n_261), .A2(n_229), .A3(n_230), .B1(n_223), .B2(n_165), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_241), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_257), .B(n_230), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_273), .B(n_208), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_250), .A2(n_219), .B1(n_218), .B2(n_216), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_247), .B(n_216), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_271), .A2(n_197), .B(n_9), .C(n_10), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_244), .A2(n_197), .B(n_10), .C(n_12), .Y(n_300) );
OAI22x1_ASAP7_75t_L g301 ( .A1(n_282), .A2(n_8), .B1(n_12), .B2(n_13), .Y(n_301) );
OAI22x1_ASAP7_75t_L g302 ( .A1(n_282), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_239), .B(n_14), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_251), .B(n_15), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_253), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_238), .A2(n_52), .B(n_77), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_265), .A2(n_51), .B(n_74), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_280), .A2(n_17), .B1(n_18), .B2(n_19), .C(n_20), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_SL g310 ( .A1(n_279), .A2(n_46), .B(n_72), .C(n_70), .Y(n_310) );
OAI211xp5_ASAP7_75t_SL g311 ( .A1(n_281), .A2(n_17), .B(n_18), .C(n_19), .Y(n_311) );
CKINVDCx11_ASAP7_75t_R g312 ( .A(n_247), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_274), .A2(n_21), .B1(n_24), .B2(n_25), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_267), .A2(n_26), .B(n_27), .C(n_28), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_251), .B(n_29), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_254), .A2(n_40), .B1(n_42), .B2(n_54), .C(n_57), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_284), .A2(n_270), .B(n_266), .Y(n_318) );
CKINVDCx14_ASAP7_75t_R g319 ( .A(n_312), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_286), .A2(n_240), .B1(n_276), .B2(n_275), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_293), .A2(n_265), .B1(n_276), .B2(n_275), .Y(n_321) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_291), .A2(n_277), .B(n_254), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_287), .A2(n_285), .B(n_300), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_305), .Y(n_325) );
OR2x6_ASAP7_75t_L g326 ( .A(n_298), .B(n_277), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_295), .B(n_241), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_284), .A2(n_268), .B(n_256), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_290), .A2(n_264), .B(n_246), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_288), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_310), .A2(n_246), .B(n_248), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
AOI221x1_ASAP7_75t_SL g334 ( .A1(n_294), .A2(n_248), .B1(n_258), .B2(n_65), .C(n_66), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_296), .B(n_317), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_312), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_287), .A2(n_245), .B(n_249), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_300), .A2(n_272), .B(n_269), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_304), .B(n_242), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_306), .A2(n_242), .B(n_262), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_283), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_283), .Y(n_343) );
AO31x2_ASAP7_75t_L g344 ( .A1(n_301), .A2(n_302), .A3(n_313), .B(n_315), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_331), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_323), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_323), .B(n_292), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_325), .B(n_292), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
AO21x2_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_307), .B(n_311), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_322), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_326), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_328), .B(n_292), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_333), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_327), .B(n_303), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_345), .B(n_307), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_345), .A2(n_289), .B1(n_308), .B2(n_316), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_318), .A2(n_329), .B(n_332), .Y(n_366) );
AO21x2_ASAP7_75t_L g367 ( .A1(n_329), .A2(n_311), .B(n_310), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g372 ( .A1(n_336), .A2(n_299), .B(n_314), .C(n_237), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_332), .A2(n_297), .B(n_61), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_369), .B(n_337), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_350), .B(n_336), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_349), .B(n_324), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_350), .B(n_334), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_324), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_321), .B(n_337), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_370), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_370), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_370), .A2(n_326), .B1(n_333), .B2(n_327), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_357), .B(n_319), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_346), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_369), .B(n_333), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_360), .A2(n_334), .B1(n_320), .B2(n_338), .C(n_326), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_364), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_349), .B(n_358), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_358), .B(n_324), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_358), .B(n_324), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_347), .B(n_324), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_347), .B(n_321), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_347), .B(n_344), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_348), .B(n_344), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_348), .B(n_344), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_369), .B(n_333), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_352), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_403), .B(n_348), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_375), .B(n_360), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_381), .B(n_360), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_403), .B(n_352), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_374), .B(n_352), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_397), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_381), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_374), .B(n_353), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_388), .B(n_365), .C(n_372), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_403), .B(n_353), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_395), .B(n_371), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_410), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_410), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_376), .B(n_353), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_376), .B(n_354), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_376), .B(n_354), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_378), .B(n_354), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_374), .B(n_369), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_385), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_378), .B(n_362), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_393), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_374), .B(n_362), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_386), .B(n_362), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_395), .B(n_371), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_378), .B(n_364), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_406), .B(n_407), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_377), .B(n_344), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_377), .B(n_344), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_393), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_396), .B(n_364), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_385), .Y(n_450) );
AND2x4_ASAP7_75t_SL g451 ( .A(n_391), .B(n_359), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_406), .B(n_344), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_374), .B(n_357), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_396), .B(n_361), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_385), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_407), .B(n_359), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
NAND2x1_ASAP7_75t_L g458 ( .A(n_408), .B(n_373), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_408), .B(n_361), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_387), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_446), .B(n_401), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_399), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_417), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_415), .B(n_396), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_447), .B(n_401), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_413), .B(n_401), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_442), .B(n_392), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_398), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_420), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_420), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_425), .B(n_398), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_412), .B(n_398), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_451), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_425), .B(n_400), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_430), .B(n_400), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_411), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_421), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_411), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_423), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_412), .B(n_400), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_445), .B(n_382), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_426), .B(n_443), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_423), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_414), .B(n_382), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_451), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_430), .B(n_380), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_424), .B(n_392), .C(n_372), .D(n_384), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_452), .B(n_384), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_433), .B(n_408), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
INVx3_ASAP7_75t_SL g499 ( .A(n_451), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_441), .A2(n_359), .B1(n_409), .B2(n_391), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_431), .B(n_380), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_431), .B(n_380), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_432), .B(n_434), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_428), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_437), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_418), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_432), .B(n_380), .Y(n_509) );
NOR2xp67_ASAP7_75t_SL g510 ( .A(n_418), .B(n_373), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_434), .B(n_404), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_454), .B(n_404), .Y(n_512) );
AOI32xp33_ASAP7_75t_L g513 ( .A1(n_438), .A2(n_365), .A3(n_391), .B1(n_409), .B2(n_408), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_440), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_436), .B(n_409), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_454), .B(n_404), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_436), .B(n_409), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_439), .B(n_391), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_439), .B(n_389), .Y(n_520) );
OR2x6_ASAP7_75t_L g521 ( .A(n_458), .B(n_394), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_437), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_418), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_465), .B(n_462), .Y(n_524) );
BUFx2_ASAP7_75t_SL g525 ( .A(n_493), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_466), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_494), .B(n_463), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_494), .B(n_463), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g529 ( .A1(n_513), .A2(n_441), .B(n_438), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_469), .B(n_448), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_471), .A2(n_441), .B(n_456), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g533 ( .A(n_495), .B(n_458), .C(n_457), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_493), .B(n_435), .Y(n_534) );
NOR2xp33_ASAP7_75t_SL g535 ( .A(n_499), .B(n_441), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_504), .B(n_435), .Y(n_536) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_471), .B(n_462), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_502), .B(n_460), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_489), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_495), .B(n_460), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_467), .B(n_457), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_505), .Y(n_543) );
AOI322xp5_ASAP7_75t_SL g544 ( .A1(n_477), .A2(n_444), .A3(n_449), .B1(n_453), .B2(n_335), .C1(n_416), .C2(n_422), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_499), .A2(n_453), .B1(n_448), .B2(n_422), .Y(n_545) );
NAND2x1_ASAP7_75t_SL g546 ( .A(n_499), .B(n_444), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_473), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_474), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_474), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_435), .Y(n_551) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_511), .B(n_449), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_479), .B(n_435), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_502), .B(n_459), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_505), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_476), .B(n_419), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_514), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_467), .A2(n_339), .B(n_335), .C(n_343), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_518), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_511), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_486), .B(n_419), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_503), .B(n_459), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_479), .B(n_419), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_512), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_484), .Y(n_567) );
OAI311xp33_ASAP7_75t_L g568 ( .A1(n_513), .A2(n_461), .A3(n_419), .B1(n_338), .C1(n_343), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_468), .B(n_461), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_485), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_480), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_500), .A2(n_461), .B1(n_453), .B2(n_450), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_523), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_488), .B(n_453), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_529), .A2(n_487), .B1(n_498), .B2(n_470), .C(n_519), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_527), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_537), .A2(n_541), .B(n_529), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_546), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_526), .B(n_503), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_532), .A2(n_517), .B1(n_515), .B2(n_491), .C(n_521), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_542), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_538), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_552), .A2(n_496), .B1(n_478), .B2(n_468), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_540), .B(n_496), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_547), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_571), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_558), .A2(n_521), .B(n_508), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_545), .B(n_521), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_530), .B(n_509), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_535), .A2(n_509), .B(n_516), .C(n_512), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_559), .B(n_472), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_557), .A2(n_497), .B(n_464), .C(n_485), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_539), .B(n_472), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_524), .B(n_475), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g601 ( .A1(n_531), .A2(n_490), .B1(n_516), .B2(n_501), .C1(n_492), .C2(n_478), .Y(n_601) );
OAI211xp5_ASAP7_75t_L g602 ( .A1(n_533), .A2(n_464), .B(n_490), .C(n_492), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_554), .B(n_475), .Y(n_603) );
OAI222xp33_ASAP7_75t_L g604 ( .A1(n_544), .A2(n_521), .B1(n_510), .B2(n_501), .C1(n_464), .C2(n_520), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_545), .A2(n_521), .B1(n_416), .B2(n_422), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_535), .A2(n_461), .B1(n_373), .B2(n_506), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_553), .B(n_416), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_534), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_575), .A2(n_564), .B1(n_569), .B2(n_565), .Y(n_609) );
AOI221x1_ASAP7_75t_SL g610 ( .A1(n_588), .A2(n_572), .B1(n_562), .B2(n_574), .C(n_534), .Y(n_610) );
OAI222xp33_ASAP7_75t_L g611 ( .A1(n_593), .A2(n_573), .B1(n_560), .B2(n_510), .C1(n_556), .C2(n_561), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_578), .A2(n_536), .B(n_551), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_587), .A2(n_543), .B1(n_555), .B2(n_573), .Y(n_613) );
AOI22xp5_ASAP7_75t_SL g614 ( .A1(n_585), .A2(n_568), .B1(n_570), .B2(n_567), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_579), .A2(n_568), .B1(n_566), .B2(n_563), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_589), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_604), .A2(n_550), .B(n_416), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_602), .A2(n_422), .B1(n_459), .B2(n_506), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_608), .Y(n_620) );
AOI211xp5_ASAP7_75t_SL g621 ( .A1(n_605), .A2(n_596), .B(n_581), .C(n_592), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_588), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_596), .A2(n_459), .B(n_507), .C(n_483), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_601), .B(n_522), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_608), .A2(n_522), .B1(n_507), .B2(n_483), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_576), .A2(n_481), .B1(n_480), .B2(n_450), .C(n_455), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_598), .A2(n_481), .B(n_373), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_577), .A2(n_351), .B1(n_450), .B2(n_455), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_610), .A2(n_583), .B1(n_582), .B2(n_584), .C(n_590), .Y(n_629) );
NOR2xp33_ASAP7_75t_R g630 ( .A(n_622), .B(n_579), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_621), .A2(n_608), .B1(n_584), .B2(n_597), .C(n_595), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_611), .A2(n_606), .B(n_580), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_618), .A2(n_594), .B1(n_600), .B2(n_599), .C(n_603), .Y(n_633) );
NAND2xp33_ASAP7_75t_SL g634 ( .A(n_620), .B(n_607), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_615), .A2(n_606), .B(n_591), .C(n_351), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_611), .A2(n_591), .B(n_373), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_609), .A2(n_351), .B1(n_342), .B2(n_343), .C(n_394), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_624), .B(n_351), .Y(n_638) );
AOI322xp5_ASAP7_75t_L g639 ( .A1(n_612), .A2(n_394), .A3(n_389), .B1(n_387), .B2(n_342), .C1(n_343), .C2(n_373), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_630), .A2(n_619), .B(n_613), .C(n_623), .Y(n_640) );
AO22x1_ASAP7_75t_L g641 ( .A1(n_638), .A2(n_627), .B1(n_614), .B2(n_617), .Y(n_641) );
NAND4xp75_ASAP7_75t_L g642 ( .A(n_637), .B(n_628), .C(n_626), .D(n_616), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g643 ( .A1(n_631), .A2(n_625), .B(n_330), .C(n_340), .Y(n_643) );
NOR3x1_ASAP7_75t_L g644 ( .A(n_632), .B(n_340), .C(n_341), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g645 ( .A(n_629), .B(n_366), .C(n_330), .D(n_389), .Y(n_645) );
NOR4xp75_ASAP7_75t_SL g646 ( .A(n_644), .B(n_633), .C(n_634), .D(n_635), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_643), .Y(n_647) );
OR5x1_ASAP7_75t_L g648 ( .A(n_640), .B(n_636), .C(n_639), .D(n_68), .E(n_69), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_641), .B(n_387), .C(n_367), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_647), .B(n_642), .C(n_645), .D(n_242), .Y(n_650) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_646), .B(n_366), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_648), .B1(n_649), .B2(n_366), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_650), .A2(n_366), .B1(n_367), .B2(n_341), .Y(n_653) );
OAI22xp5_ASAP7_75t_SL g654 ( .A1(n_652), .A2(n_366), .B1(n_367), .B2(n_80), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_654), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_653), .B(n_341), .Y(n_656) );
AO21x2_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_367), .B(n_67), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_367), .B1(n_366), .B2(n_59), .Y(n_658) );
endmodule