module real_jpeg_9404_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_24),
.B1(n_62),
.B2(n_63),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_12),
.B(n_34),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_3),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_33),
.B(n_44),
.C(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_9),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_92),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_92),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_92),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_10),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_87),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_87),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_87),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_46),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_12),
.B(n_46),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_12),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_12),
.A2(n_33),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_33),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_37),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_12),
.A2(n_25),
.B1(n_27),
.B2(n_112),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_13),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_99),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_99),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_14),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_128),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_128),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_25),
.B1(n_27),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_15),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_16),
.A2(n_25),
.B1(n_27),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_16),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_17),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_147),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_147),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_17),
.A2(n_25),
.B1(n_27),
.B2(n_147),
.Y(n_279)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_74),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_23),
.A2(n_28),
.B1(n_37),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_30),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_25),
.A2(n_30),
.B(n_112),
.C(n_177),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_28),
.A2(n_37),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_29),
.A2(n_32),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_29),
.A2(n_32),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_29),
.A2(n_32),
.B1(n_210),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_29),
.A2(n_32),
.B1(n_235),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_29),
.A2(n_32),
.B1(n_253),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_29),
.A2(n_32),
.B1(n_53),
.B2(n_279),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_66),
.C(n_68),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_39),
.A2(n_40),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_51),
.C(n_57),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_306),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_43),
.A2(n_45),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_43),
.A2(n_45),
.B1(n_138),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_43),
.A2(n_45),
.B1(n_155),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_43),
.A2(n_45),
.B1(n_195),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_43),
.A2(n_45),
.B1(n_206),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_43),
.A2(n_45),
.B1(n_232),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_44),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_45),
.B(n_112),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_59),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_46),
.B(n_48),
.Y(n_142)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_47),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_51),
.A2(n_52),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_57),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_57),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_65),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_61),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_61),
.B1(n_98),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_58),
.A2(n_61),
.B1(n_125),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_58),
.A2(n_61),
.B1(n_134),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_58),
.A2(n_61),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_58),
.A2(n_61),
.B1(n_218),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_58),
.A2(n_61),
.B1(n_227),
.B2(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_61),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_62),
.B(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_65),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_66),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_70),
.A2(n_71),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_324),
.B(n_330),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_297),
.A3(n_317),
.B1(n_322),
.B2(n_323),
.C(n_333),
.Y(n_75)
);

AOI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_243),
.A3(n_285),
.B1(n_291),
.B2(n_296),
.C(n_334),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_200),
.C(n_239),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_170),
.B(n_199),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_149),
.B(n_169),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_130),
.B(n_148),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_119),
.B(n_129),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_105),
.B(n_118),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_93),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_88),
.A2(n_89),
.B1(n_146),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_109),
.B1(n_110),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_104),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_104),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_113),
.B(n_117),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_110),
.B1(n_127),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_109),
.A2(n_110),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_109),
.A2(n_110),
.B1(n_181),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_109),
.A2(n_110),
.B1(n_215),
.B2(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_109),
.A2(n_110),
.B(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_121),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.C(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.CI(n_139),
.CON(n_132),
.SN(n_132)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_162),
.B2(n_163),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_165),
.C(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_159),
.C(n_161),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_185),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_184),
.C(n_185),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_193),
.C(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_190),
.A2(n_192),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_201),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_220),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_202),
.B(n_220),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_219),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_219),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_237),
.B2(n_238),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_228),
.C(n_238),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_226),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_241),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_262),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_244),
.B(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_255),
.C(n_261),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_246),
.B1(n_255),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_251),
.C(n_254),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_257),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_278),
.B(n_281),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_258),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_283),
.B2(n_284),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_275),
.C(n_284),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_270),
.B(n_273),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_272),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_273),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_273),
.A2(n_299),
.B1(n_308),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_282),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_310),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_308),
.C(n_309),
.Y(n_298)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_301),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_306),
.C(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_312),
.C(n_316),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_304),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);


endmodule