module fake_jpeg_6398_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_3),
.B(n_0),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx4f_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

AND2x6_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_19),
.B(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_7),
.B1(n_12),
.B2(n_9),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_9),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_5),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_11),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_15),
.B(n_13),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_17),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_33),
.A3(n_27),
.B1(n_25),
.B2(n_28),
.C1(n_13),
.C2(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_27),
.C(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.C(n_21),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_27),
.B1(n_33),
.B2(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_40),
.C(n_34),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_35),
.B(n_40),
.C(n_11),
.Y(n_43)
);


endmodule