module real_aes_18419_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g910 ( .A(n_0), .Y(n_910) );
INVx1_ASAP7_75t_L g601 ( .A(n_1), .Y(n_601) );
AOI221x1_ASAP7_75t_SL g625 ( .A1(n_1), .A2(n_3), .B1(n_626), .B2(n_629), .C(n_631), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g1341 ( .A1(n_2), .A2(n_6), .B1(n_395), .B2(n_617), .Y(n_1341) );
AOI22xp33_ASAP7_75t_SL g1378 ( .A1(n_2), .A2(n_224), .B1(n_985), .B2(n_1077), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_3), .A2(n_23), .B1(n_605), .B2(n_606), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_4), .A2(n_767), .B(n_771), .C(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g793 ( .A(n_4), .Y(n_793) );
AOI221x1_ASAP7_75t_SL g921 ( .A1(n_5), .A2(n_240), .B1(n_922), .B2(n_923), .C(n_925), .Y(n_921) );
AOI21xp33_ASAP7_75t_L g982 ( .A1(n_5), .A2(n_513), .B(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_6), .A2(n_225), .B1(n_548), .B2(n_985), .Y(n_1383) );
CKINVDCx5p33_ASAP7_75t_R g1111 ( .A(n_7), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_8), .A2(n_203), .B1(n_461), .B2(n_465), .C(n_470), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_8), .A2(n_203), .B1(n_516), .B2(n_521), .Y(n_515) );
INVx1_ASAP7_75t_L g657 ( .A(n_9), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_9), .A2(n_424), .B(n_684), .C(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_10), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_10), .A2(n_28), .B1(n_385), .B2(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g457 ( .A(n_11), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_11), .A2(n_243), .B1(n_505), .B2(n_510), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_12), .A2(n_235), .B1(n_279), .B2(n_446), .C(n_448), .Y(n_445) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_12), .A2(n_64), .B1(n_132), .B2(n_371), .C1(n_534), .C2(n_535), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_13), .A2(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g643 ( .A(n_13), .Y(n_643) );
INVx1_ASAP7_75t_L g313 ( .A(n_14), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_14), .B(n_263), .Y(n_392) );
AND2x2_ASAP7_75t_L g443 ( .A(n_14), .B(n_307), .Y(n_443) );
AND2x2_ASAP7_75t_L g452 ( .A(n_14), .B(n_213), .Y(n_452) );
INVx1_ASAP7_75t_L g811 ( .A(n_15), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g851 ( .A1(n_15), .A2(n_114), .B1(n_510), .B2(n_852), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g814 ( .A1(n_16), .A2(n_241), .B1(n_461), .B2(n_465), .C(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g848 ( .A(n_16), .Y(n_848) );
INVx1_ASAP7_75t_L g892 ( .A(n_17), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_18), .A2(n_170), .B1(n_837), .B2(n_1001), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_18), .A2(n_90), .B1(n_264), .B2(n_1015), .C(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1353 ( .A(n_19), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_19), .A2(n_35), .B1(n_1365), .B2(n_1367), .Y(n_1364) );
INVx1_ASAP7_75t_L g1359 ( .A(n_20), .Y(n_1359) );
INVx1_ASAP7_75t_L g1101 ( .A(n_21), .Y(n_1101) );
INVx2_ASAP7_75t_L g1158 ( .A(n_22), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_22), .B(n_1159), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_22), .B(n_101), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_23), .A2(n_167), .B1(n_629), .B2(n_638), .C(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g864 ( .A(n_24), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_25), .A2(n_129), .B1(n_495), .B2(n_943), .Y(n_942) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_25), .A2(n_217), .B1(n_951), .B2(n_953), .C(n_955), .Y(n_950) );
AOI22xp5_ASAP7_75t_SL g1171 ( .A1(n_26), .A2(n_128), .B1(n_1163), .B2(n_1165), .Y(n_1171) );
AOI22xp5_ASAP7_75t_SL g1183 ( .A1(n_27), .A2(n_237), .B1(n_1160), .B2(n_1184), .Y(n_1183) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_28), .Y(n_342) );
INVx1_ASAP7_75t_L g868 ( .A(n_29), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_30), .A2(n_199), .B1(n_835), .B2(n_1099), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g1116 ( .A1(n_30), .A2(n_60), .B1(n_589), .B2(n_1117), .C(n_1119), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_31), .A2(n_75), .B1(n_395), .B2(n_606), .Y(n_1405) );
INVx1_ASAP7_75t_L g1431 ( .A(n_31), .Y(n_1431) );
INVx1_ASAP7_75t_L g282 ( .A(n_32), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_33), .A2(n_173), .B1(n_429), .B2(n_430), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_33), .A2(n_173), .B1(n_299), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g681 ( .A(n_34), .Y(n_681) );
INVx1_ASAP7_75t_L g1357 ( .A(n_35), .Y(n_1357) );
INVx1_ASAP7_75t_L g1041 ( .A(n_36), .Y(n_1041) );
INVx1_ASAP7_75t_L g656 ( .A(n_37), .Y(n_656) );
INVx1_ASAP7_75t_L g742 ( .A(n_38), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_39), .A2(n_166), .B1(n_1155), .B2(n_1160), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_40), .A2(n_212), .B1(n_382), .B2(n_1015), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_40), .A2(n_107), .B1(n_1073), .B2(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g863 ( .A(n_41), .Y(n_863) );
INVx1_ASAP7_75t_L g1360 ( .A(n_42), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_43), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_44), .A2(n_77), .B1(n_546), .B2(n_968), .Y(n_998) );
INVx1_ASAP7_75t_L g1032 ( .A(n_44), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_45), .A2(n_150), .B1(n_297), .B2(n_304), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_45), .A2(n_150), .B1(n_703), .B2(n_705), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_46), .A2(n_126), .B1(n_279), .B2(n_448), .C(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_46), .A2(n_78), .B1(n_835), .B2(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_47), .A2(n_97), .B1(n_1163), .B2(n_1189), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_48), .A2(n_84), .B1(n_1155), .B2(n_1163), .Y(n_1174) );
INVx1_ASAP7_75t_L g354 ( .A(n_49), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_49), .A2(n_124), .B1(n_382), .B2(n_384), .Y(n_381) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_50), .A2(n_169), .B1(n_492), .B2(n_553), .Y(n_584) );
INVx1_ASAP7_75t_L g588 ( .A(n_50), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_51), .A2(n_159), .B1(n_617), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_51), .A2(n_100), .B1(n_626), .B2(n_840), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_52), .A2(n_172), .B1(n_1163), .B2(n_1184), .Y(n_1203) );
INVx1_ASAP7_75t_L g326 ( .A(n_53), .Y(n_326) );
INVx1_ASAP7_75t_L g333 ( .A(n_53), .Y(n_333) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_54), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_54), .A2(n_235), .B1(n_546), .B2(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g726 ( .A(n_55), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_56), .A2(n_246), .B1(n_1155), .B2(n_1160), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_57), .A2(n_72), .B1(n_395), .B2(n_1117), .Y(n_1346) );
INVx1_ASAP7_75t_L g1377 ( .A(n_57), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_58), .Y(n_930) );
INVx1_ASAP7_75t_L g1415 ( .A(n_59), .Y(n_1415) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_60), .A2(n_178), .B1(n_534), .B2(n_546), .Y(n_1108) );
INVx1_ASAP7_75t_L g1140 ( .A(n_61), .Y(n_1140) );
INVx2_ASAP7_75t_L g352 ( .A(n_62), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_63), .A2(n_136), .B1(n_712), .B2(n_895), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_63), .A2(n_136), .B1(n_661), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_64), .A2(n_147), .B1(n_382), .B2(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_65), .A2(n_144), .B1(n_297), .B2(n_304), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_65), .A2(n_144), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g278 ( .A(n_66), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_67), .A2(n_69), .B1(n_1155), .B2(n_1163), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_68), .A2(n_210), .B1(n_497), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g826 ( .A(n_70), .Y(n_826) );
INVx1_ASAP7_75t_L g1349 ( .A(n_71), .Y(n_1349) );
INVxp67_ASAP7_75t_SL g1382 ( .A(n_72), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_73), .A2(n_122), .B1(n_427), .B2(n_889), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_73), .A2(n_122), .B1(n_304), .B2(n_898), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_74), .A2(n_105), .B1(n_481), .B2(n_483), .C(n_924), .Y(n_1409) );
INVxp67_ASAP7_75t_SL g1419 ( .A(n_74), .Y(n_1419) );
INVxp67_ASAP7_75t_SL g1421 ( .A(n_75), .Y(n_1421) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_76), .A2(n_378), .B(n_654), .C(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g709 ( .A(n_76), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_77), .A2(n_115), .B1(n_1014), .B2(n_1015), .C(n_1016), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_78), .Y(n_818) );
INVx1_ASAP7_75t_L g1105 ( .A(n_79), .Y(n_1105) );
INVx1_ASAP7_75t_L g550 ( .A(n_80), .Y(n_550) );
INVx1_ASAP7_75t_L g775 ( .A(n_81), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g784 ( .A1(n_81), .A2(n_591), .B(n_785), .C(n_789), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_82), .A2(n_163), .B1(n_927), .B2(n_928), .Y(n_1050) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_82), .B(n_1091), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_83), .A2(n_186), .B1(n_1160), .B2(n_1165), .Y(n_1173) );
INVx1_ASAP7_75t_L g1355 ( .A(n_85), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_86), .Y(n_1009) );
INVx1_ASAP7_75t_L g608 ( .A(n_87), .Y(n_608) );
INVx1_ASAP7_75t_L g745 ( .A(n_88), .Y(n_745) );
INVx1_ASAP7_75t_L g744 ( .A(n_89), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_90), .A2(n_117), .B1(n_626), .B2(n_840), .Y(n_1097) );
OA222x2_ASAP7_75t_L g912 ( .A1(n_91), .A2(n_200), .B1(n_217), .B2(n_913), .C1(n_915), .C2(n_919), .Y(n_912) );
INVx1_ASAP7_75t_L g966 ( .A(n_91), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g1394 ( .A1(n_92), .A2(n_1395), .B1(n_1396), .B2(n_1444), .Y(n_1394) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_92), .Y(n_1444) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_93), .A2(n_650), .B1(n_651), .B2(n_713), .Y(n_649) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_93), .Y(n_713) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_94), .A2(n_441), .B(n_444), .C(n_453), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_94), .A2(n_205), .B1(n_491), .B2(n_497), .Y(n_490) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_95), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_95), .B(n_1140), .Y(n_1156) );
XNOR2xp5_ASAP7_75t_L g438 ( .A(n_96), .B(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_98), .A2(n_149), .B1(n_1155), .B2(n_1160), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_99), .Y(n_1005) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_100), .A2(n_148), .B1(n_807), .B2(n_820), .C(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g1159 ( .A(n_101), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_101), .B(n_1158), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_102), .A2(n_189), .B1(n_264), .B2(n_385), .Y(n_1055) );
INVxp67_ASAP7_75t_SL g1071 ( .A(n_102), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_103), .A2(n_183), .B1(n_1155), .B2(n_1160), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_104), .A2(n_109), .B1(n_629), .B2(n_762), .Y(n_999) );
INVx1_ASAP7_75t_L g1035 ( .A(n_104), .Y(n_1035) );
INVx1_ASAP7_75t_L g1429 ( .A(n_105), .Y(n_1429) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_106), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g1402 ( .A1(n_107), .A2(n_180), .B1(n_448), .B2(n_924), .C(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g994 ( .A(n_108), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_108), .A2(n_221), .B1(n_274), .B2(n_473), .Y(n_1025) );
INVx1_ASAP7_75t_L g1018 ( .A(n_109), .Y(n_1018) );
INVx2_ASAP7_75t_L g351 ( .A(n_110), .Y(n_351) );
INVx1_ASAP7_75t_L g365 ( .A(n_110), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_110), .B(n_352), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_111), .A2(n_223), .B1(n_777), .B2(n_778), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_111), .A2(n_223), .B1(n_795), .B2(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g668 ( .A(n_112), .Y(n_668) );
INVx1_ASAP7_75t_L g870 ( .A(n_113), .Y(n_870) );
INVx1_ASAP7_75t_L g812 ( .A(n_114), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_115), .A2(n_152), .B1(n_546), .B2(n_845), .Y(n_1003) );
AOI22xp5_ASAP7_75t_SL g1179 ( .A1(n_116), .A2(n_242), .B1(n_1163), .B2(n_1165), .Y(n_1179) );
INVx1_ASAP7_75t_L g1121 ( .A(n_117), .Y(n_1121) );
INVx1_ASAP7_75t_L g286 ( .A(n_118), .Y(n_286) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_119), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_119), .A2(n_218), .B1(n_473), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_120), .A2(n_239), .B1(n_617), .B2(n_809), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_120), .A2(n_220), .B1(n_630), .B2(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g893 ( .A(n_121), .Y(n_893) );
OAI211xp5_ASAP7_75t_L g899 ( .A1(n_121), .A2(n_292), .B(n_378), .C(n_900), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_123), .B(n_466), .Y(n_1412) );
INVxp67_ASAP7_75t_SL g1440 ( .A(n_123), .Y(n_1440) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_124), .Y(n_321) );
INVx1_ASAP7_75t_L g677 ( .A(n_125), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_126), .A2(n_164), .B1(n_534), .B2(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1062 ( .A(n_127), .Y(n_1062) );
INVx1_ASAP7_75t_L g563 ( .A(n_128), .Y(n_563) );
INVx1_ASAP7_75t_L g967 ( .A(n_129), .Y(n_967) );
INVx1_ASAP7_75t_L g1224 ( .A(n_130), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_131), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_132), .A2(n_209), .B1(n_481), .B2(n_482), .C(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g729 ( .A(n_133), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_134), .Y(n_733) );
INVx1_ASAP7_75t_L g873 ( .A(n_135), .Y(n_873) );
INVx1_ASAP7_75t_L g1112 ( .A(n_137), .Y(n_1112) );
INVx1_ASAP7_75t_L g1411 ( .A(n_138), .Y(n_1411) );
INVx1_ASAP7_75t_L g1414 ( .A(n_139), .Y(n_1414) );
OAI322xp33_ASAP7_75t_L g1417 ( .A1(n_139), .A2(n_346), .A3(n_573), .B1(n_1418), .B2(n_1422), .C1(n_1428), .C2(n_1435), .Y(n_1417) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_140), .A2(n_179), .B1(n_1163), .B2(n_1189), .Y(n_1188) );
BUFx3_ASAP7_75t_L g324 ( .A(n_141), .Y(n_324) );
INVx1_ASAP7_75t_L g680 ( .A(n_142), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_143), .A2(n_248), .B1(n_264), .B2(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_143), .A2(n_190), .B1(n_957), .B2(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1399 ( .A(n_145), .Y(n_1399) );
INVx1_ASAP7_75t_L g1340 ( .A(n_146), .Y(n_1340) );
INVx1_ASAP7_75t_L g544 ( .A(n_147), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_148), .A2(n_159), .B1(n_762), .B2(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g327 ( .A(n_151), .Y(n_327) );
AOI211xp5_ASAP7_75t_SL g1029 ( .A1(n_152), .A2(n_1030), .B(n_1031), .C(n_1034), .Y(n_1029) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_153), .Y(n_1103) );
INVx1_ASAP7_75t_L g1134 ( .A(n_154), .Y(n_1134) );
AOI22xp5_ASAP7_75t_L g1162 ( .A1(n_154), .A2(n_211), .B1(n_1163), .B2(n_1165), .Y(n_1162) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_155), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_156), .A2(n_192), .B1(n_840), .B2(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1017 ( .A(n_156), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_157), .A2(n_193), .B1(n_885), .B2(n_1064), .C(n_1066), .Y(n_1063) );
INVx1_ASAP7_75t_L g1083 ( .A(n_157), .Y(n_1083) );
OAI22xp33_ASAP7_75t_SL g1051 ( .A1(n_158), .A2(n_204), .B1(n_935), .B2(n_1033), .Y(n_1051) );
INVx1_ASAP7_75t_L g1086 ( .A(n_158), .Y(n_1086) );
AOI21xp5_ASAP7_75t_SL g1058 ( .A1(n_160), .A2(n_483), .B(n_611), .Y(n_1058) );
INVx1_ASAP7_75t_L g1070 ( .A(n_160), .Y(n_1070) );
INVx1_ASAP7_75t_L g1053 ( .A(n_161), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_161), .A2(n_248), .B1(n_957), .B2(n_1077), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_162), .Y(n_1057) );
INVx1_ASAP7_75t_L g1085 ( .A(n_163), .Y(n_1085) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_164), .Y(n_816) );
INVx1_ASAP7_75t_L g367 ( .A(n_165), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_167), .A2(n_481), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g260 ( .A(n_168), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_169), .Y(n_595) );
INVx1_ASAP7_75t_L g1120 ( .A(n_170), .Y(n_1120) );
INVx1_ASAP7_75t_L g270 ( .A(n_171), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_174), .Y(n_991) );
INVx1_ASAP7_75t_L g1350 ( .A(n_175), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_176), .Y(n_1437) );
XOR2x2_ASAP7_75t_L g798 ( .A(n_177), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1132 ( .A(n_178), .Y(n_1132) );
INVx1_ASAP7_75t_L g1426 ( .A(n_180), .Y(n_1426) );
INVx1_ASAP7_75t_L g723 ( .A(n_181), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_182), .A2(n_215), .B1(n_227), .B2(n_497), .C1(n_566), .C2(n_571), .Y(n_565) );
INVx1_ASAP7_75t_L g1407 ( .A(n_184), .Y(n_1407) );
XOR2xp5_ASAP7_75t_L g858 ( .A(n_185), .B(n_859), .Y(n_858) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_186), .B(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_187), .A2(n_247), .B1(n_605), .B2(n_606), .Y(n_604) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_187), .Y(n_641) );
INVx1_ASAP7_75t_L g866 ( .A(n_188), .Y(n_866) );
INVxp67_ASAP7_75t_L g1075 ( .A(n_189), .Y(n_1075) );
AOI21xp33_ASAP7_75t_L g1054 ( .A1(n_190), .A2(n_611), .B(n_612), .Y(n_1054) );
INVx1_ASAP7_75t_L g774 ( .A(n_191), .Y(n_774) );
INVx1_ASAP7_75t_L g1037 ( .A(n_192), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_193), .Y(n_1088) );
INVx1_ASAP7_75t_L g355 ( .A(n_194), .Y(n_355) );
INVx1_ASAP7_75t_L g675 ( .A(n_195), .Y(n_675) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
INVx1_ASAP7_75t_L g671 ( .A(n_197), .Y(n_671) );
INVx1_ASAP7_75t_L g685 ( .A(n_198), .Y(n_685) );
INVx1_ASAP7_75t_L g1133 ( .A(n_199), .Y(n_1133) );
INVx1_ASAP7_75t_L g956 ( .A(n_200), .Y(n_956) );
INVx1_ASAP7_75t_L g336 ( .A(n_201), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_202), .Y(n_947) );
INVx1_ASAP7_75t_L g1089 ( .A(n_204), .Y(n_1089) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_206), .A2(n_216), .B1(n_661), .B2(n_663), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_206), .A2(n_216), .B1(n_711), .B2(n_712), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_207), .Y(n_582) );
INVx1_ASAP7_75t_L g738 ( .A(n_208), .Y(n_738) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_209), .Y(n_542) );
OAI211xp5_ASAP7_75t_L g801 ( .A1(n_210), .A2(n_802), .B(n_803), .C(n_810), .Y(n_801) );
INVxp67_ASAP7_75t_SL g1423 ( .A(n_212), .Y(n_1423) );
BUFx3_ASAP7_75t_L g263 ( .A(n_213), .Y(n_263) );
INVx1_ASAP7_75t_L g307 ( .A(n_213), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_214), .Y(n_437) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_218), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_219), .Y(n_934) );
INVx1_ASAP7_75t_L g926 ( .A(n_220), .Y(n_926) );
INVx1_ASAP7_75t_L g1039 ( .A(n_221), .Y(n_1039) );
INVx1_ASAP7_75t_L g683 ( .A(n_222), .Y(n_683) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_224), .Y(n_1344) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_225), .Y(n_1345) );
INVx1_ASAP7_75t_L g317 ( .A(n_226), .Y(n_317) );
INVx1_ASAP7_75t_L g364 ( .A(n_226), .Y(n_364) );
INVx2_ASAP7_75t_L g391 ( .A(n_226), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_227), .A2(n_232), .B1(n_615), .B2(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g1339 ( .A(n_228), .Y(n_1339) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_229), .A2(n_245), .B1(n_1155), .B2(n_1160), .Y(n_1170) );
INVx1_ASAP7_75t_L g874 ( .A(n_230), .Y(n_874) );
OAI211xp5_ASAP7_75t_L g890 ( .A1(n_231), .A2(n_767), .B(n_771), .C(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g901 ( .A(n_231), .Y(n_901) );
INVx1_ASAP7_75t_L g583 ( .A(n_232), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_233), .Y(n_948) );
INVx1_ASAP7_75t_L g1044 ( .A(n_234), .Y(n_1044) );
INVx1_ASAP7_75t_L g871 ( .A(n_236), .Y(n_871) );
INVx1_ASAP7_75t_L g1222 ( .A(n_238), .Y(n_1222) );
XNOR2xp5_ASAP7_75t_L g1335 ( .A(n_238), .B(n_1336), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_238), .A2(n_1391), .B1(n_1393), .B2(n_1445), .Y(n_1390) );
INVx1_ASAP7_75t_L g980 ( .A(n_239), .Y(n_980) );
INVx1_ASAP7_75t_L g979 ( .A(n_240), .Y(n_979) );
INVx1_ASAP7_75t_L g850 ( .A(n_241), .Y(n_850) );
INVx1_ASAP7_75t_L g454 ( .A(n_243), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g996 ( .A(n_244), .Y(n_996) );
INVx1_ASAP7_75t_L g632 ( .A(n_247), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_1137), .B(n_1145), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_857), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_715), .B1(n_716), .B2(n_856), .Y(n_251) );
INVx1_ASAP7_75t_L g856 ( .A(n_252), .Y(n_856) );
OA22x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_560), .B2(n_561), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
XNOR2x1_ASAP7_75t_L g254 ( .A(n_255), .B(n_438), .Y(n_254) );
XOR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_437), .Y(n_255) );
NAND3x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_318), .C(n_402), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_296), .B(n_310), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_277), .C(n_292), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B1(n_270), .B2(n_271), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_260), .A2(n_270), .B1(n_419), .B2(n_422), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g1348 ( .A1(n_261), .A2(n_271), .B1(n_1349), .B2(n_1350), .C(n_1351), .Y(n_1348) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g273 ( .A(n_262), .B(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g284 ( .A(n_262), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g790 ( .A(n_262), .B(n_285), .Y(n_790) );
BUFx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g289 ( .A(n_263), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g295 ( .A(n_263), .Y(n_295) );
AND2x4_ASAP7_75t_L g399 ( .A(n_263), .B(n_313), .Y(n_399) );
INVx3_ASAP7_75t_L g383 ( .A(n_264), .Y(n_383) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_264), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g1026 ( .A1(n_264), .A2(n_598), .B(n_996), .C(n_1027), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_L g1126 ( .A1(n_264), .A2(n_1105), .B(n_1127), .C(n_1129), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g396 ( .A(n_265), .Y(n_396) );
AND2x2_ASAP7_75t_L g456 ( .A(n_265), .B(n_443), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_265), .B(n_452), .Y(n_556) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
OR2x2_ASAP7_75t_L g377 ( .A(n_266), .B(n_269), .Y(n_377) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_266), .Y(n_597) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_267), .B(n_269), .Y(n_281) );
INVx1_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_267), .B(n_269), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_267), .B(n_309), .Y(n_308) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_267), .B(n_269), .Y(n_380) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
INVx2_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
AND2x2_ASAP7_75t_L g386 ( .A(n_269), .B(n_276), .Y(n_386) );
INVx1_ASAP7_75t_L g903 ( .A(n_271), .Y(n_903) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g664 ( .A(n_273), .Y(n_664) );
INVx8_ASAP7_75t_L g478 ( .A(n_274), .Y(n_478) );
BUFx2_ASAP7_75t_L g817 ( .A(n_274), .Y(n_817) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI222xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B1(n_282), .B2(n_283), .C1(n_286), .C2(n_287), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_278), .A2(n_282), .B1(n_286), .B2(n_405), .C1(n_410), .C2(n_413), .Y(n_404) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_280), .B(n_294), .Y(n_293) );
AND2x6_ASAP7_75t_L g451 ( .A(n_280), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_SL g464 ( .A(n_280), .B(n_443), .Y(n_464) );
BUFx3_ASAP7_75t_L g482 ( .A(n_280), .Y(n_482) );
INVx1_ASAP7_75t_L g821 ( .A(n_280), .Y(n_821) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_280), .Y(n_924) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_280), .Y(n_1030) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g788 ( .A(n_281), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_283), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_283), .A2(n_791), .B1(n_892), .B2(n_901), .Y(n_900) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g468 ( .A(n_285), .Y(n_468) );
BUFx2_ASAP7_75t_L g594 ( .A(n_285), .Y(n_594) );
INVx1_ASAP7_75t_L g945 ( .A(n_285), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_285), .A2(n_596), .B1(n_991), .B2(n_1009), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_285), .B(n_294), .Y(n_1354) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g658 ( .A(n_289), .Y(n_658) );
INVx2_ASAP7_75t_L g792 ( .A(n_289), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_290), .B(n_452), .Y(n_496) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g654 ( .A(n_293), .Y(n_654) );
AND2x2_ASAP7_75t_L g786 ( .A(n_294), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
AND2x4_ASAP7_75t_L g484 ( .A(n_295), .B(n_313), .Y(n_484) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g898 ( .A(n_298), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_298), .B(n_1144), .Y(n_1143) );
AOI22xp33_ASAP7_75t_SL g1358 ( .A1(n_298), .A2(n_305), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AND2x4_ASAP7_75t_SL g1387 ( .A(n_298), .B(n_1388), .Y(n_1387) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
OR2x6_ASAP7_75t_L g662 ( .A(n_300), .B(n_306), .Y(n_662) );
INVxp67_ASAP7_75t_L g725 ( .A(n_300), .Y(n_725) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g473 ( .A(n_301), .Y(n_473) );
BUFx4f_ASAP7_75t_L g692 ( .A(n_301), .Y(n_692) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx3_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx4_ASAP7_75t_L g783 ( .A(n_305), .Y(n_783) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g447 ( .A(n_308), .Y(n_447) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_308), .Y(n_459) );
BUFx3_ASAP7_75t_L g481 ( .A(n_308), .Y(n_481) );
BUFx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_311), .A2(n_653), .A3(n_659), .B(n_660), .Y(n_652) );
BUFx3_ASAP7_75t_L g797 ( .A(n_311), .Y(n_797) );
INVx1_ASAP7_75t_L g1361 ( .A(n_311), .Y(n_1361) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g1144 ( .A(n_312), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_312), .B(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g495 ( .A(n_315), .B(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_L g503 ( .A(n_315), .Y(n_503) );
INVx1_ASAP7_75t_L g570 ( .A(n_315), .Y(n_570) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_373), .Y(n_318) );
OAI33xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_335), .A3(n_346), .B1(n_353), .B2(n_359), .B3(n_366), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_327), .B2(n_328), .Y(n_320) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_322), .A2(n_354), .B1(n_355), .B2(n_356), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_322), .A2(n_930), .B1(n_936), .B2(n_974), .C(n_975), .Y(n_973) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x4_ASAP7_75t_L g420 ( .A(n_323), .B(n_421), .Y(n_420) );
OR2x4_ASAP7_75t_L g429 ( .A(n_323), .B(n_362), .Y(n_429) );
INVx2_ASAP7_75t_L g507 ( .A(n_323), .Y(n_507) );
BUFx4f_ASAP7_75t_L g642 ( .A(n_323), .Y(n_642) );
BUFx3_ASAP7_75t_L g753 ( .A(n_323), .Y(n_753) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_324), .Y(n_334) );
INVx2_ASAP7_75t_L g341 ( .A(n_324), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_324), .B(n_333), .Y(n_345) );
AND2x4_ASAP7_75t_L g416 ( .A(n_324), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g500 ( .A(n_325), .Y(n_500) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g340 ( .A(n_326), .Y(n_340) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_327), .A2(n_355), .B1(n_375), .B2(n_378), .C(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g684 ( .A(n_329), .Y(n_684) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g1427 ( .A(n_330), .Y(n_1427) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
BUFx2_ASAP7_75t_L g756 ( .A(n_331), .Y(n_756) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
BUFx2_ASAP7_75t_L g412 ( .A(n_332), .Y(n_412) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g417 ( .A(n_333), .Y(n_417) );
BUFx2_ASAP7_75t_L g409 ( .A(n_334), .Y(n_409) );
INVx2_ASAP7_75t_L g518 ( .A(n_334), .Y(n_518) );
AND2x4_ASAP7_75t_L g630 ( .A(n_334), .B(n_526), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_342), .B2(n_343), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_336), .A2(n_367), .B1(n_375), .B2(n_378), .C(n_381), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_337), .A2(n_343), .B1(n_1339), .B2(n_1377), .C(n_1378), .Y(n_1376) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g368 ( .A(n_338), .Y(n_368) );
AND2x4_ASAP7_75t_L g431 ( .A(n_338), .B(n_421), .Y(n_431) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_338), .Y(n_762) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_338), .Y(n_978) );
INVx2_ASAP7_75t_L g1380 ( .A(n_338), .Y(n_1380) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx8_ASAP7_75t_L g513 ( .A(n_339), .Y(n_513) );
INVx2_ASAP7_75t_L g536 ( .A(n_339), .Y(n_536) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_339), .Y(n_628) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x4_ASAP7_75t_L g499 ( .A(n_341), .B(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x6_ASAP7_75t_L g423 ( .A(n_344), .B(n_362), .Y(n_423) );
INVx1_ASAP7_75t_L g765 ( .A(n_344), .Y(n_765) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g372 ( .A(n_345), .Y(n_372) );
OAI33xp33_ASAP7_75t_L g666 ( .A1(n_346), .A2(n_537), .A3(n_667), .B1(n_674), .B2(n_678), .B3(n_682), .Y(n_666) );
OAI33xp33_ASAP7_75t_L g861 ( .A1(n_346), .A2(n_537), .A3(n_862), .B1(n_865), .B2(n_869), .B3(n_872), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g1067 ( .A1(n_346), .A2(n_1068), .B1(n_1074), .B2(n_1078), .Y(n_1067) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx4f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g528 ( .A(n_348), .Y(n_528) );
BUFx8_ASAP7_75t_L g749 ( .A(n_348), .Y(n_749) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g401 ( .A(n_349), .Y(n_401) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_349), .Y(n_436) );
OR2x2_ASAP7_75t_L g493 ( .A(n_349), .B(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g983 ( .A(n_350), .Y(n_983) );
NAND2xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_352), .Y(n_350) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_351), .Y(n_434) );
INVx1_ASAP7_75t_L g502 ( .A(n_351), .Y(n_502) );
AND3x4_ASAP7_75t_L g647 ( .A(n_351), .B(n_408), .C(n_623), .Y(n_647) );
INVx3_ASAP7_75t_L g362 ( .A(n_352), .Y(n_362) );
BUFx3_ASAP7_75t_L g408 ( .A(n_352), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_356), .A2(n_506), .B1(n_873), .B2(n_874), .Y(n_872) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g673 ( .A(n_357), .Y(n_673) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g492 ( .A(n_358), .B(n_493), .Y(n_492) );
INVx4_ASAP7_75t_L g636 ( .A(n_358), .Y(n_636) );
INVx3_ASAP7_75t_L g645 ( .A(n_358), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_360), .A2(n_558), .B1(n_625), .B2(n_637), .C(n_646), .Y(n_624) );
INVx2_ASAP7_75t_L g1078 ( .A(n_360), .Y(n_1078) );
INVx2_ASAP7_75t_L g1435 ( .A(n_360), .Y(n_1435) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g539 ( .A(n_361), .Y(n_539) );
OAI33xp33_ASAP7_75t_L g748 ( .A1(n_361), .A2(n_749), .A3(n_750), .B1(n_757), .B2(n_760), .B3(n_766), .Y(n_748) );
NAND3x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .C(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g421 ( .A(n_362), .Y(n_421) );
AND2x4_ASAP7_75t_L g425 ( .A(n_362), .B(n_416), .Y(n_425) );
AND2x4_ASAP7_75t_L g501 ( .A(n_362), .B(n_502), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g843 ( .A(n_362), .B(n_365), .Y(n_843) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g520 ( .A(n_364), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_364), .B(n_443), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_370), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_865) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g543 ( .A(n_371), .Y(n_543) );
CKINVDCx8_ASAP7_75t_R g759 ( .A(n_371), .Y(n_759) );
INVx3_ASAP7_75t_L g1381 ( .A(n_371), .Y(n_1381) );
INVx1_ASAP7_75t_L g1430 ( .A(n_371), .Y(n_1430) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g554 ( .A(n_372), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_387), .B1(n_393), .B2(n_397), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_375), .A2(n_866), .B1(n_870), .B2(n_882), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_375), .A2(n_484), .B1(n_609), .B2(n_1017), .C(n_1018), .Y(n_1016) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g694 ( .A(n_376), .Y(n_694) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g732 ( .A(n_377), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_377), .Y(n_737) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_377), .Y(n_1033) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_378), .A2(n_736), .B1(n_1339), .B2(n_1340), .C(n_1341), .Y(n_1338) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx4_ASAP7_75t_L g592 ( .A(n_379), .Y(n_592) );
BUFx4f_ASAP7_75t_L g695 ( .A(n_379), .Y(n_695) );
BUFx4f_ASAP7_75t_L g734 ( .A(n_379), .Y(n_734) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_379), .Y(n_885) );
BUFx4f_ASAP7_75t_L g935 ( .A(n_379), .Y(n_935) );
OR2x6_ASAP7_75t_L g938 ( .A(n_379), .B(n_939), .Y(n_938) );
OAI221xp5_ASAP7_75t_L g1131 ( .A1(n_379), .A2(n_399), .B1(n_1033), .B2(n_1132), .C(n_1133), .Y(n_1131) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g741 ( .A(n_380), .Y(n_741) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g1014 ( .A(n_383), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g442 ( .A(n_385), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g450 ( .A(n_385), .Y(n_450) );
INVx1_ASAP7_75t_L g1118 ( .A(n_385), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g606 ( .A(n_386), .Y(n_606) );
INVx2_ASAP7_75t_L g618 ( .A(n_386), .Y(n_618) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_386), .Y(n_1015) );
OAI33xp33_ASAP7_75t_L g721 ( .A1(n_387), .A2(n_397), .A3(n_722), .B1(n_728), .B2(n_735), .B3(n_743), .Y(n_721) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_387), .A2(n_697), .A3(n_876), .B1(n_881), .B2(n_883), .B3(n_886), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g1337 ( .A1(n_387), .A2(n_699), .B1(n_1338), .B2(n_1342), .Y(n_1337) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g687 ( .A(n_389), .Y(n_687) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g487 ( .A(n_390), .Y(n_487) );
OR2x6_ASAP7_75t_L g842 ( .A(n_390), .B(n_843), .Y(n_842) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g623 ( .A(n_391), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_391), .B(n_452), .Y(n_941) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g605 ( .A(n_396), .Y(n_605) );
INVx2_ASAP7_75t_L g809 ( .A(n_396), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g932 ( .A1(n_397), .A2(n_933), .B(n_938), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_SL g448 ( .A(n_399), .Y(n_448) );
INVx4_ASAP7_75t_L g612 ( .A(n_399), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_399), .B(n_400), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g1031 ( .A1(n_399), .A2(n_1032), .B(n_1033), .Y(n_1031) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_426), .B(n_432), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_418), .C(n_424), .Y(n_403) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g708 ( .A(n_406), .Y(n_708) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
AND2x4_ASAP7_75t_L g411 ( .A(n_407), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g773 ( .A(n_407), .B(n_409), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g1080 ( .A1(n_407), .A2(n_1081), .B(n_1084), .C(n_1087), .Y(n_1080) );
AND2x4_ASAP7_75t_L g1366 ( .A(n_407), .B(n_409), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_407), .B(n_412), .Y(n_1368) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_410), .A2(n_656), .B1(n_708), .B2(n_709), .Y(n_707) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_411), .A2(n_773), .B1(n_774), .B2(n_775), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_411), .A2(n_773), .B1(n_892), .B2(n_893), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_411), .A2(n_773), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g534 ( .A(n_416), .Y(n_534) );
BUFx3_ASAP7_75t_L g548 ( .A(n_416), .Y(n_548) );
BUFx2_ASAP7_75t_L g559 ( .A(n_416), .Y(n_559) );
INVx2_ASAP7_75t_L g846 ( .A(n_416), .Y(n_846) );
BUFx2_ASAP7_75t_L g968 ( .A(n_416), .Y(n_968) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_416), .Y(n_1077) );
INVx1_ASAP7_75t_L g526 ( .A(n_417), .Y(n_526) );
INVx1_ASAP7_75t_L g711 ( .A(n_419), .Y(n_711) );
INVx2_ASAP7_75t_L g895 ( .A(n_419), .Y(n_895) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g777 ( .A(n_420), .Y(n_777) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_420), .Y(n_1091) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_422), .A2(n_1349), .B1(n_1350), .B2(n_1372), .Y(n_1371) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g712 ( .A(n_423), .Y(n_712) );
INVx1_ASAP7_75t_L g779 ( .A(n_423), .Y(n_779) );
CKINVDCx8_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
CKINVDCx8_ASAP7_75t_R g771 ( .A(n_425), .Y(n_771) );
OAI31xp33_ASAP7_75t_L g1079 ( .A1(n_425), .A2(n_1080), .A3(n_1090), .B(n_1092), .Y(n_1079) );
AOI211xp5_ASAP7_75t_L g1363 ( .A1(n_425), .A2(n_1073), .B(n_1355), .C(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g704 ( .A(n_429), .Y(n_704) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_429), .Y(n_1370) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g705 ( .A(n_431), .Y(n_705) );
INVx1_ASAP7_75t_L g889 ( .A(n_431), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_431), .A2(n_1359), .B1(n_1360), .B2(n_1370), .Y(n_1369) );
OAI31xp33_ASAP7_75t_L g701 ( .A1(n_432), .A2(n_702), .A3(n_706), .B(n_710), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g887 ( .A1(n_432), .A2(n_888), .A3(n_890), .B(n_894), .Y(n_887) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_433), .B(n_435), .Y(n_432) );
AND2x2_ASAP7_75t_L g780 ( .A(n_433), .B(n_435), .Y(n_780) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_433), .B(n_435), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_433), .B(n_435), .Y(n_1374) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
O2A1O1Ixp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_460), .B(n_485), .C(n_488), .Y(n_439) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g802 ( .A(n_442), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_442), .A2(n_458), .B1(n_1414), .B2(n_1415), .Y(n_1413) );
AND2x4_ASAP7_75t_L g458 ( .A(n_443), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g578 ( .A(n_443), .B(n_459), .Y(n_578) );
AND2x2_ASAP7_75t_L g616 ( .A(n_443), .B(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_443), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_449), .B(n_451), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g807 ( .A(n_447), .Y(n_807) );
AOI21xp5_ASAP7_75t_SL g803 ( .A1(n_451), .A2(n_804), .B(n_808), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_451), .A2(n_1402), .B1(n_1405), .B2(n_1406), .C(n_1407), .Y(n_1401) );
INVx1_ASAP7_75t_L g469 ( .A(n_452), .Y(n_469) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_452), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_457), .B2(n_458), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_455), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
AOI221xp5_ASAP7_75t_SL g1408 ( .A1(n_455), .A2(n_1409), .B1(n_1410), .B2(n_1411), .C(n_1412), .Y(n_1408) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g569 ( .A(n_456), .B(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_458), .Y(n_813) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_459), .Y(n_611) );
INVx2_ASAP7_75t_L g1024 ( .A(n_459), .Y(n_1024) );
INVx1_ASAP7_75t_L g1404 ( .A(n_459), .Y(n_1404) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g619 ( .A(n_462), .Y(n_619) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g1406 ( .A(n_464), .Y(n_1406) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g1065 ( .A(n_468), .Y(n_1065) );
INVx1_ASAP7_75t_L g1129 ( .A(n_469), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B1(n_475), .B2(n_479), .C(n_480), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_471), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_471), .A2(n_816), .B1(n_817), .B2(n_818), .C(n_819), .Y(n_815) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g927 ( .A(n_473), .Y(n_927) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_474), .A2(n_530), .B(n_533), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_475), .A2(n_668), .B1(n_683), .B2(n_689), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_475), .A2(n_677), .B1(n_681), .B2(n_689), .Y(n_700) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_477), .A2(n_1035), .B1(n_1036), .B2(n_1037), .Y(n_1034) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g727 ( .A(n_478), .Y(n_727) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_478), .Y(n_747) );
INVx1_ASAP7_75t_L g880 ( .A(n_478), .Y(n_880) );
INVx2_ASAP7_75t_L g929 ( .A(n_478), .Y(n_929) );
INVx2_ASAP7_75t_L g1125 ( .A(n_478), .Y(n_1125) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g603 ( .A(n_484), .Y(n_603) );
INVx3_ASAP7_75t_L g822 ( .A(n_484), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_484), .A2(n_609), .B1(n_694), .B2(n_1120), .C(n_1121), .Y(n_1119) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI31xp67_ASAP7_75t_L g949 ( .A1(n_486), .A2(n_950), .A3(n_960), .B(n_972), .Y(n_949) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_514), .C(n_549), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_504), .Y(n_489) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
AND2x4_ASAP7_75t_L g828 ( .A(n_492), .B(n_495), .Y(n_828) );
INVx2_ASAP7_75t_L g990 ( .A(n_492), .Y(n_990) );
INVx1_ASAP7_75t_L g509 ( .A(n_493), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_493), .Y(n_512) );
OR2x2_ASAP7_75t_L g553 ( .A(n_493), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g971 ( .A(n_494), .Y(n_971) );
INVx5_ASAP7_75t_L g1040 ( .A(n_497), .Y(n_1040) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_503), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
BUFx3_ASAP7_75t_L g532 ( .A(n_499), .Y(n_532) );
INVx8_ASAP7_75t_L g547 ( .A(n_499), .Y(n_547) );
BUFx3_ASAP7_75t_L g835 ( .A(n_499), .Y(n_835) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_499), .Y(n_962) );
AND2x4_ASAP7_75t_L g519 ( .A(n_501), .B(n_520), .Y(n_519) );
AND2x6_ASAP7_75t_L g952 ( .A(n_501), .B(n_517), .Y(n_952) );
AND2x2_ASAP7_75t_L g954 ( .A(n_501), .B(n_525), .Y(n_954) );
INVx1_ASAP7_75t_L g959 ( .A(n_501), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_568), .Y(n_567) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx2_ASAP7_75t_SL g670 ( .A(n_506), .Y(n_670) );
OR2x2_ASAP7_75t_L g852 ( .A(n_506), .B(n_508), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_506), .A2(n_644), .B1(n_863), .B2(n_864), .Y(n_862) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g634 ( .A(n_507), .Y(n_634) );
INVxp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g574 ( .A(n_509), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_511), .B(n_1005), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_511), .B(n_1101), .Y(n_1100) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x4_ASAP7_75t_L g992 ( .A(n_512), .B(n_993), .Y(n_992) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_512), .B(n_993), .Y(n_1443) );
INVx2_ASAP7_75t_SL g639 ( .A(n_513), .Y(n_639) );
INVx3_ASAP7_75t_L g679 ( .A(n_513), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_527), .Y(n_514) );
INVx2_ASAP7_75t_L g581 ( .A(n_516), .Y(n_581) );
NAND2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_519), .Y(n_516) );
AND2x2_ASAP7_75t_L g849 ( .A(n_517), .B(n_519), .Y(n_849) );
AND2x4_ASAP7_75t_SL g1008 ( .A(n_517), .B(n_519), .Y(n_1008) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g522 ( .A(n_519), .B(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g558 ( .A(n_519), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_SL g1010 ( .A(n_519), .B(n_523), .Y(n_1010) );
OR2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_522), .A2(n_581), .B1(n_582), .B2(n_583), .C(n_584), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_522), .A2(n_848), .B1(n_849), .B2(n_850), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g1439 ( .A1(n_522), .A2(n_558), .B1(n_1008), .B2(n_1407), .C(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_529), .B1(n_537), .B2(n_540), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g1375 ( .A1(n_528), .A2(n_537), .B1(n_1376), .B2(n_1379), .Y(n_1375) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g1434 ( .A(n_532), .Y(n_1434) );
INVx1_ASAP7_75t_L g541 ( .A(n_535), .Y(n_541) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g575 ( .A(n_536), .Y(n_575) );
BUFx2_ASAP7_75t_L g867 ( .A(n_536), .Y(n_867) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_543), .B2(n_544), .C(n_545), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_543), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_543), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_543), .A2(n_639), .B1(n_870), .B2(n_871), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_546), .A2(n_628), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
INVx8_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_547), .Y(n_957) );
INVx3_ASAP7_75t_L g985 ( .A(n_547), .Y(n_985) );
INVx2_ASAP7_75t_L g993 ( .A(n_547), .Y(n_993) );
A2O1A1Ixp33_ASAP7_75t_L g955 ( .A1(n_548), .A2(n_956), .B(n_957), .C(n_958), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_548), .A2(n_1062), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_557), .Y(n_549) );
AOI21xp33_ASAP7_75t_SL g825 ( .A1(n_551), .A2(n_826), .B(n_827), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g1436 ( .A1(n_551), .A2(n_1437), .B(n_1438), .Y(n_1436) );
INVx8_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g995 ( .A(n_553), .Y(n_995) );
INVx1_ASAP7_75t_L g914 ( .A(n_555), .Y(n_914) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g854 ( .A(n_558), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_558), .A2(n_1008), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1110 ( .A1(n_558), .A2(n_1008), .B1(n_1010), .B2(n_1111), .C(n_1112), .Y(n_1110) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AO22x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_648), .B1(n_649), .B2(n_714), .Y(n_561) );
INVx1_ASAP7_75t_SL g714 ( .A(n_562), .Y(n_714) );
XNOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_579), .Y(n_564) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_569), .A2(n_577), .B1(n_947), .B2(n_948), .Y(n_946) );
AND2x4_ASAP7_75t_L g577 ( .A(n_570), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g758 ( .A(n_575), .Y(n_758) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND3xp33_ASAP7_75t_SL g579 ( .A(n_580), .B(n_585), .C(n_624), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_582), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_614), .B(n_620), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_599), .C(n_607), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_590), .C(n_598), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_SL g1061 ( .A1(n_589), .A2(n_598), .B(n_1062), .C(n_1063), .Y(n_1061) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g600 ( .A(n_592), .Y(n_600) );
INVx2_ASAP7_75t_L g609 ( .A(n_592), .Y(n_609) );
INVx2_ASAP7_75t_L g882 ( .A(n_592), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_594), .A2(n_596), .B1(n_1103), .B2(n_1111), .Y(n_1128) );
INVx1_ASAP7_75t_L g1066 ( .A(n_596), .Y(n_1066) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_602), .C(n_604), .Y(n_599) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_610), .C(n_613), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_608), .A2(n_632), .B1(n_633), .B2(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g916 ( .A(n_617), .B(n_917), .Y(n_916) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g1060 ( .A(n_618), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g824 ( .A(n_621), .Y(n_824) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI31xp33_ASAP7_75t_L g1012 ( .A1(n_622), .A2(n_1013), .A3(n_1019), .B(n_1029), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_622), .Y(n_1047) );
OAI31xp33_ASAP7_75t_L g1115 ( .A1(n_622), .A2(n_1116), .A3(n_1122), .B(n_1130), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1416 ( .A(n_622), .Y(n_1416) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g676 ( .A(n_626), .Y(n_676) );
INVx8_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx3_ASAP7_75t_L g1420 ( .A(n_627), .Y(n_1420) );
INVx5_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g964 ( .A(n_628), .Y(n_964) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_628), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_629), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_965) );
BUFx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx5_ASAP7_75t_L g838 ( .A(n_630), .Y(n_838) );
BUFx3_ASAP7_75t_L g840 ( .A(n_630), .Y(n_840) );
BUFx12f_ASAP7_75t_L g1082 ( .A(n_630), .Y(n_1082) );
BUFx4f_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g767 ( .A(n_636), .Y(n_767) );
INVx2_ASAP7_75t_L g974 ( .A(n_636), .Y(n_974) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g981 ( .A1(n_644), .A2(n_934), .B(n_982), .C(n_984), .Y(n_981) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI33xp33_ASAP7_75t_L g831 ( .A1(n_647), .A2(n_832), .A3(n_836), .B1(n_839), .B2(n_841), .B3(n_844), .Y(n_831) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_647), .A2(n_841), .A3(n_998), .B1(n_999), .B2(n_1000), .B3(n_1003), .Y(n_997) );
NAND3xp33_ASAP7_75t_L g1096 ( .A(n_647), .B(n_1097), .C(n_1098), .Y(n_1096) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_665), .C(n_701), .Y(n_651) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_662), .Y(n_795) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g796 ( .A(n_664), .Y(n_796) );
NOR2xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_686), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_669), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_671), .A2(n_685), .B1(n_694), .B2(n_695), .Y(n_696) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_675), .A2(n_680), .B1(n_694), .B2(n_695), .Y(n_693) );
OAI33xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .A3(n_693), .B1(n_696), .B2(n_697), .B3(n_700), .Y(n_686) );
INVx1_ASAP7_75t_L g931 ( .A(n_687), .Y(n_931) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_692), .Y(n_878) );
INVx4_ASAP7_75t_L g1036 ( .A(n_692), .Y(n_1036) );
OAI22xp33_ASAP7_75t_SL g883 ( .A1(n_694), .A2(n_864), .B1(n_874), .B2(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_798), .B2(n_855), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_768), .C(n_781), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_748), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_726), .B2(n_727), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_723), .A2(n_738), .B1(n_751), .B2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_726), .A2(n_742), .B1(n_751), .B2(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_733), .B2(n_734), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_729), .A2(n_744), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g1343 ( .A(n_731), .Y(n_1343) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_733), .A2(n_745), .B1(n_761), .B2(n_763), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B1(n_739), .B2(n_742), .Y(n_735) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_736), .A2(n_934), .B1(n_935), .B2(n_936), .C(n_937), .Y(n_933) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx5_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g919 ( .A(n_741), .B(n_918), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_741), .B(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_741), .B(n_1128), .Y(n_1127) );
INVx5_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_SL g1425 ( .A(n_753), .Y(n_1425) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_758), .A2(n_759), .B1(n_1057), .B2(n_1075), .C(n_1076), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_759), .A2(n_977), .B1(n_979), .B2(n_980), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g1068 ( .A1(n_759), .A2(n_1069), .B1(n_1070), .B2(n_1071), .C(n_1072), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_759), .A2(n_1419), .B1(n_1420), .B2(n_1421), .Y(n_1418) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI31xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .A3(n_776), .B(n_780), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_774), .A2(n_790), .B1(n_791), .B2(n_793), .Y(n_789) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI31xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .A3(n_794), .B(n_797), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g1351 ( .A(n_785), .B(n_1352), .C(n_1356), .Y(n_1351) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g1352 ( .A1(n_791), .A2(n_1353), .B1(n_1354), .B2(n_1355), .Y(n_1352) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI31xp33_ASAP7_75t_SL g896 ( .A1(n_797), .A2(n_897), .A3(n_899), .B(n_902), .Y(n_896) );
INVx1_ASAP7_75t_L g855 ( .A(n_798), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_825), .C(n_829), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_814), .B(n_823), .Y(n_800) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g922 ( .A(n_806), .Y(n_922) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g1398 ( .A(n_828), .Y(n_1398) );
NOR3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_851), .C(n_853), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_831), .B(n_847), .Y(n_830) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g1106 ( .A(n_841), .B(n_1107), .C(n_1108), .Y(n_1106) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx3_ASAP7_75t_L g975 ( .A(n_843), .Y(n_975) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g1073 ( .A(n_846), .Y(n_1073) );
INVx1_ASAP7_75t_L g1099 ( .A(n_846), .Y(n_1099) );
INVx2_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_904), .B1(n_905), .B2(n_1136), .Y(n_857) );
INVx1_ASAP7_75t_L g1136 ( .A(n_858), .Y(n_1136) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_887), .C(n_896), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_875), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_863), .A2(n_873), .B1(n_877), .B2(n_879), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_868), .A2(n_871), .B1(n_877), .B2(n_879), .Y(n_886) );
INVx2_ASAP7_75t_SL g877 ( .A(n_878), .Y(n_877) );
BUFx3_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OAI221xp5_ASAP7_75t_L g1342 ( .A1(n_885), .A2(n_1343), .B1(n_1344), .B2(n_1345), .C(n_1346), .Y(n_1342) );
INVx3_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
BUFx3_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OA22x2_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B1(n_1042), .B2(n_1135), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
XOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_986), .Y(n_908) );
XNOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NAND4xp75_ASAP7_75t_L g911 ( .A(n_912), .B(n_920), .C(n_946), .D(n_949), .Y(n_911) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
AOI211x1_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_931), .B(n_932), .C(n_942), .Y(n_920) );
BUFx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_924), .A2(n_1005), .B1(n_1011), .B2(n_1023), .C(n_1025), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g1123 ( .A1(n_924), .A2(n_1023), .B1(n_1101), .B2(n_1112), .C(n_1124), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_924), .B(n_1357), .Y(n_1356) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_928), .B2(n_930), .Y(n_925) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OAI211xp5_ASAP7_75t_SL g1052 ( .A1(n_935), .A2(n_1053), .B(n_1054), .C(n_1055), .Y(n_1052) );
OAI211xp5_ASAP7_75t_SL g1056 ( .A1(n_935), .A2(n_1057), .B(n_1058), .C(n_1059), .Y(n_1056) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
NAND2x2_ASAP7_75t_L g943 ( .A(n_940), .B(n_944), .Y(n_943) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_SL g944 ( .A(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_947), .A2(n_948), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx4_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
AOI21xp33_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_965), .B(n_969), .Y(n_960) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI21xp5_ASAP7_75t_SL g972 ( .A1(n_973), .A2(n_976), .B(n_981), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g1428 ( .A1(n_977), .A2(n_1429), .B1(n_1430), .B2(n_1431), .C(n_1432), .Y(n_1428) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_978), .Y(n_1069) );
XNOR2x1_ASAP7_75t_L g986 ( .A(n_987), .B(n_1041), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_988), .B(n_1006), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_997), .C(n_1004), .Y(n_988) );
AOI222xp33_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B1(n_992), .B2(n_994), .C1(n_995), .C2(n_996), .Y(n_989) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_990), .A2(n_992), .B1(n_995), .B2(n_1103), .C1(n_1104), .C2(n_1105), .Y(n_1102) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
NAND3xp33_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1012), .C(n_1038), .Y(n_1006) );
OAI21xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1022), .B(n_1026), .Y(n_1019) );
OAI21xp5_ASAP7_75t_SL g1122 ( .A1(n_1020), .A2(n_1123), .B(n_1126), .Y(n_1122) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1049 ( .A1(n_1021), .A2(n_1050), .B(n_1051), .Y(n_1049) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1040), .B(n_1114), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1040), .B(n_1415), .Y(n_1441) );
XNOR2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1093), .Y(n_1042) );
XOR2xp5_ASAP7_75t_L g1135 ( .A(n_1043), .B(n_1093), .Y(n_1135) );
XNOR2x1_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1079), .Y(n_1045) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1048), .B(n_1067), .Y(n_1046) );
NAND4xp25_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1052), .C(n_1056), .D(n_1061), .Y(n_1048) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1091), .Y(n_1372) );
XNOR2x1_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1134), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1109), .Y(n_1094) );
NAND4xp25_ASAP7_75t_SL g1095 ( .A(n_1096), .B(n_1100), .C(n_1102), .D(n_1106), .Y(n_1095) );
NAND3xp33_ASAP7_75t_SL g1109 ( .A(n_1110), .B(n_1113), .C(n_1115), .Y(n_1109) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1143), .Y(n_1137) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1138), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1141), .Y(n_1138) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1139), .B(n_1142), .Y(n_1392) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1139), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
NOR2xp33_ASAP7_75t_L g1449 ( .A(n_1142), .B(n_1446), .Y(n_1449) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1332), .B1(n_1333), .B2(n_1384), .C(n_1390), .Y(n_1145) );
NOR2xp67_ASAP7_75t_SL g1146 ( .A(n_1147), .B(n_1270), .Y(n_1146) );
NAND4xp25_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1226), .C(n_1250), .D(n_1264), .Y(n_1147) );
OAI21xp5_ASAP7_75t_L g1148 ( .A1(n_1149), .A2(n_1210), .B(n_1216), .Y(n_1148) );
OAI321xp33_ASAP7_75t_L g1149 ( .A1(n_1150), .A2(n_1175), .A3(n_1186), .B1(n_1190), .B2(n_1193), .C(n_1196), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1151), .B(n_1228), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1167), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1152), .B(n_1194), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1152), .B(n_1168), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1152), .B(n_1242), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1152), .B(n_1243), .Y(n_1316) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1153), .B(n_1215), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1153), .B(n_1169), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1153), .B(n_1243), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1153), .B(n_1279), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1153), .B(n_1243), .Y(n_1302) );
NAND2xp5_ASAP7_75t_SL g1311 ( .A(n_1153), .B(n_1201), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_1153), .B(n_1201), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1162), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1154), .B(n_1162), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
AND2x6_ASAP7_75t_L g1160 ( .A(n_1156), .B(n_1161), .Y(n_1160) );
AND2x6_ASAP7_75t_L g1163 ( .A(n_1156), .B(n_1164), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1156), .B(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1156), .B(n_1166), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1156), .B(n_1166), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1156), .B(n_1157), .Y(n_1221) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_1157), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1160), .Y(n_1223) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1172), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1169), .B(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1169), .Y(n_1243) );
AOI321xp33_ASAP7_75t_L g1264 ( .A1(n_1169), .A2(n_1227), .A3(n_1260), .B1(n_1265), .B2(n_1267), .C(n_1269), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1169), .B(n_1172), .Y(n_1279) );
NAND2x1p5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1172), .Y(n_1195) );
NOR2xp33_ASAP7_75t_L g1199 ( .A(n_1172), .B(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1172), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1172), .B(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1176), .B(n_1230), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1181), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1177), .B(n_1186), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1177), .B(n_1192), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1177), .B(n_1186), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1177), .B(n_1209), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1177), .B(n_1182), .Y(n_1261) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1177), .Y(n_1277) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1177), .Y(n_1300) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1178), .B(n_1209), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1181), .B(n_1192), .Y(n_1191) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1181), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1181), .B(n_1230), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1181), .B(n_1231), .Y(n_1255) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1182), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1185), .Y(n_1182) );
INVx3_ASAP7_75t_L g1192 ( .A(n_1186), .Y(n_1192) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1186), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
OAI322xp33_ASAP7_75t_L g1295 ( .A1(n_1191), .A2(n_1193), .A3(n_1233), .B1(n_1296), .B2(n_1298), .C1(n_1299), .C2(n_1300), .Y(n_1295) );
CKINVDCx14_ASAP7_75t_R g1284 ( .A(n_1192), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1192), .B(n_1266), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1192), .B(n_1247), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1192), .B(n_1208), .Y(n_1330) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1193), .Y(n_1256) );
AOI21xp33_ASAP7_75t_SL g1257 ( .A1(n_1193), .A2(n_1258), .B(n_1259), .Y(n_1257) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1194), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1194), .B(n_1233), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1194), .B(n_1297), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1194), .B(n_1311), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1199), .B1(n_1205), .B2(n_1206), .Y(n_1196) );
OAI21xp5_ASAP7_75t_L g1293 ( .A1(n_1197), .A2(n_1241), .B(n_1294), .Y(n_1293) );
CKINVDCx14_ASAP7_75t_R g1197 ( .A(n_1198), .Y(n_1197) );
NOR3xp33_ASAP7_75t_L g1269 ( .A(n_1198), .B(n_1201), .C(n_1240), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1198), .B(n_1204), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1204), .Y(n_1200) );
INVx4_ASAP7_75t_L g1207 ( .A(n_1201), .Y(n_1207) );
INVx4_ASAP7_75t_L g1231 ( .A(n_1201), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1201), .B(n_1252), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1201), .B(n_1302), .Y(n_1317) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1201), .B(n_1261), .Y(n_1319) );
AND2x4_ASAP7_75t_SL g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1205), .B(n_1231), .Y(n_1281) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1206), .Y(n_1213) );
AOI21xp33_ASAP7_75t_L g1280 ( .A1(n_1206), .A2(n_1215), .B(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1206), .B(n_1263), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
CKINVDCx5p33_ASAP7_75t_R g1228 ( .A(n_1207), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1207), .B(n_1214), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1207), .B(n_1232), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1207), .B(n_1316), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1208), .B(n_1212), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1271 ( .A1(n_1208), .A2(n_1243), .B1(n_1249), .B2(n_1272), .C(n_1273), .Y(n_1271) );
NOR3xp33_ASAP7_75t_L g1309 ( .A(n_1208), .B(n_1310), .C(n_1312), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_1208), .A2(n_1277), .B1(n_1315), .B2(n_1317), .Y(n_1314) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
AOI21xp33_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1213), .B(n_1214), .Y(n_1210) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1211), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1212), .B(n_1238), .Y(n_1237) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_1212), .A2(n_1251), .B1(n_1253), .B2(n_1254), .C(n_1257), .Y(n_1250) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1212), .Y(n_1321) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1214), .Y(n_1275) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
OAI321xp33_ASAP7_75t_L g1270 ( .A1(n_1217), .A2(n_1218), .A3(n_1271), .B1(n_1282), .B2(n_1285), .C(n_1308), .Y(n_1270) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1220), .B(n_1231), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1222), .B1(n_1223), .B2(n_1224), .C(n_1225), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_1221), .Y(n_1332) );
O2A1O1Ixp33_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1229), .B(n_1234), .C(n_1235), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1228), .B(n_1246), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1228), .B(n_1265), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1232), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1230), .B(n_1263), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_1231), .Y(n_1230) );
NAND2xp5_ASAP7_75t_SL g1274 ( .A(n_1231), .B(n_1275), .Y(n_1274) );
NAND2x1_ASAP7_75t_L g1287 ( .A(n_1231), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1232), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1233), .B(n_1242), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1233), .B(n_1278), .Y(n_1307) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1234), .Y(n_1312) );
OAI221xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1239), .B1(n_1240), .B2(n_1244), .C(n_1248), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
OAI21xp5_ASAP7_75t_SL g1248 ( .A1(n_1237), .A2(n_1245), .B(n_1249), .Y(n_1248) );
INVxp67_ASAP7_75t_L g1303 ( .A(n_1238), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1239), .B(n_1328), .Y(n_1327) );
OAI32xp33_ASAP7_75t_L g1329 ( .A1(n_1240), .A2(n_1247), .A3(n_1268), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1242), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1242), .B(n_1255), .C(n_1263), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1242), .B(n_1323), .Y(n_1331) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_1247), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_1247), .A2(n_1274), .B1(n_1276), .B2(n_1278), .C(n_1280), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1256), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1262), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1261), .B(n_1263), .Y(n_1328) );
OAI21xp33_ASAP7_75t_L g1313 ( .A1(n_1263), .A2(n_1314), .B(n_1318), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1265 ( .A(n_1266), .Y(n_1265) );
OAI322xp33_ASAP7_75t_L g1320 ( .A1(n_1266), .A2(n_1268), .A3(n_1307), .B1(n_1321), .B2(n_1322), .C1(n_1325), .C2(n_1326), .Y(n_1320) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
AOI21xp33_ASAP7_75t_L g1282 ( .A1(n_1272), .A2(n_1283), .B(n_1284), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_1276), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1279), .B(n_1323), .Y(n_1322) );
CKINVDCx14_ASAP7_75t_R g1292 ( .A(n_1283), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1283), .B(n_1319), .Y(n_1318) );
O2A1O1Ixp33_ASAP7_75t_L g1301 ( .A1(n_1284), .A2(n_1302), .B(n_1303), .C(n_1304), .Y(n_1301) );
NOR5xp2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1289), .C(n_1295), .D(n_1301), .E(n_1305), .Y(n_1285) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1288), .Y(n_1326) );
A2O1A1Ixp33_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1291), .B(n_1292), .C(n_1293), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1307), .Y(n_1305) );
NOR5xp2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1313), .C(n_1320), .D(n_1327), .E(n_1329), .Y(n_1308) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NOR4xp25_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1347), .C(n_1362), .D(n_1375), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g1379 ( .A1(n_1340), .A2(n_1380), .B1(n_1381), .B2(n_1382), .C(n_1383), .Y(n_1379) );
AOI21xp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1358), .B(n_1361), .Y(n_1347) );
AOI31xp33_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1369), .A3(n_1371), .B(n_1373), .Y(n_1362) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVxp67_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
CKINVDCx20_ASAP7_75t_R g1384 ( .A(n_1385), .Y(n_1384) );
CKINVDCx20_ASAP7_75t_R g1385 ( .A(n_1386), .Y(n_1385) );
INVx3_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
BUFx3_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVxp33_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_SL g1396 ( .A(n_1397), .B(n_1436), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1399), .B1(n_1400), .B2(n_1416), .C(n_1417), .Y(n_1397) );
NAND3xp33_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1408), .C(n_1413), .Y(n_1400) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_1404), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1411), .B(n_1443), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_1423), .A2(n_1424), .B1(n_1426), .B2(n_1427), .Y(n_1422) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
NAND3xp33_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1441), .C(n_1442), .Y(n_1438) );
OAI21xp5_ASAP7_75t_L g1445 ( .A1(n_1446), .A2(n_1447), .B(n_1448), .Y(n_1445) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
endmodule