module fake_jpeg_25386_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_48),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_58),
.B1(n_70),
.B2(n_47),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_21),
.B1(n_17),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_62),
.B1(n_73),
.B2(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_30),
.B1(n_32),
.B2(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_29),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_42),
.B1(n_34),
.B2(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_18),
.B1(n_22),
.B2(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_89),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_18),
.B1(n_22),
.B2(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_95),
.C(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_22),
.B1(n_39),
.B2(n_2),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_77),
.B1(n_10),
.B2(n_11),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_15),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_39),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_13),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_105),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_1),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_72),
.B1(n_68),
.B2(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_77),
.B1(n_65),
.B2(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_1),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_104),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_1),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_71),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_47),
.C(n_5),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_4),
.C(n_6),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_99),
.C(n_102),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_65),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_106),
.B(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_101),
.B1(n_92),
.B2(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_71),
.Y(n_122)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_82),
.B1(n_77),
.B2(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_80),
.B(n_10),
.C(n_11),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_47),
.C(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_86),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g132 ( 
.A(n_121),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_81),
.C(n_89),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_138),
.C(n_143),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_95),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

OAI31xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_88),
.A3(n_104),
.B(n_83),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_140),
.A3(n_120),
.B1(n_115),
.B2(n_133),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_79),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_89),
.C(n_78),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_144),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_153),
.B1(n_125),
.B2(n_109),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_98),
.C(n_107),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_108),
.B(n_137),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_123),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_86),
.B1(n_66),
.B2(n_12),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_159),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_172),
.B(n_127),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_120),
.B(n_115),
.C(n_108),
.D(n_113),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_108),
.C(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_171),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_149),
.C(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_127),
.C(n_144),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_110),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_162),
.C(n_156),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_144),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_185),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_127),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_183),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_118),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_159),
.B1(n_158),
.B2(n_154),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_193),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_156),
.C(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_165),
.B(n_157),
.C(n_162),
.D(n_160),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_164),
.C(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_177),
.B1(n_178),
.B2(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_203),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_189),
.A2(n_168),
.B1(n_185),
.B2(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_194),
.C(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_188),
.C(n_206),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_191),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_196),
.B(n_194),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_R g217 ( 
.A1(n_211),
.A2(n_167),
.B(n_179),
.C(n_155),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_193),
.B(n_197),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_199),
.B(n_204),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_215),
.B(n_216),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_199),
.C(n_192),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_208),
.B(n_171),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.B(n_168),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_218),
.A2(n_211),
.B(n_180),
.Y(n_221)
);

AOI321xp33_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_222),
.A3(n_127),
.B1(n_180),
.B2(n_12),
.C(n_7),
.Y(n_223)
);

AOI211xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_109),
.B(n_11),
.C(n_7),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_86),
.Y(n_225)
);


endmodule