module real_aes_6706_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_725, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_725;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g444 ( .A1(n_0), .A2(n_182), .B(n_445), .C(n_448), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_1), .B(n_439), .Y(n_449) );
INVx1_ASAP7_75t_L g687 ( .A(n_2), .Y(n_687) );
INVx1_ASAP7_75t_L g217 ( .A(n_3), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_4), .B(n_134), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_5), .A2(n_434), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_6), .A2(n_157), .B(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_7), .A2(n_38), .B1(n_127), .B2(n_151), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_8), .B(n_157), .Y(n_229) );
AND2x6_ASAP7_75t_L g142 ( .A(n_9), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_10), .A2(n_142), .B(n_425), .C(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_11), .B(n_39), .Y(n_688) );
INVx1_ASAP7_75t_L g123 ( .A(n_12), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_13), .B(n_132), .Y(n_165) );
INVx1_ASAP7_75t_L g209 ( .A(n_14), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g705 ( .A1(n_15), .A2(n_75), .B1(n_706), .B2(n_707), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_15), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_16), .B(n_134), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_17), .B(n_158), .Y(n_196) );
AO32x2_ASAP7_75t_L g179 ( .A1(n_18), .A2(n_156), .A3(n_157), .B1(n_180), .B2(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_19), .B(n_127), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_20), .B(n_158), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_21), .A2(n_55), .B1(n_127), .B2(n_151), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g154 ( .A1(n_22), .A2(n_82), .B1(n_127), .B2(n_132), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_23), .B(n_127), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_24), .A2(n_156), .B(n_425), .C(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_25), .A2(n_156), .B(n_425), .C(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_26), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_27), .B(n_119), .Y(n_238) );
OAI22xp5_ASAP7_75t_SL g679 ( .A1(n_28), .A2(n_93), .B1(n_680), .B2(n_681), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_28), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_29), .A2(n_678), .B1(n_679), .B2(n_682), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_29), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_30), .A2(n_434), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_31), .B(n_119), .Y(n_144) );
INVx2_ASAP7_75t_L g129 ( .A(n_32), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_33), .A2(n_431), .B(n_457), .C(n_458), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_34), .B(n_127), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_35), .B(n_119), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_36), .A2(n_43), .B1(n_415), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_36), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_37), .B(n_167), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_40), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_41), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_42), .B(n_134), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g109 ( .A1(n_43), .A2(n_110), .B1(n_415), .B2(n_416), .Y(n_109) );
INVx1_ASAP7_75t_L g415 ( .A(n_43), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_44), .B(n_434), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_45), .A2(n_431), .B(n_457), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_46), .B(n_127), .Y(n_224) );
INVx1_ASAP7_75t_L g446 ( .A(n_47), .Y(n_446) );
AOI22xp5_ASAP7_75t_SL g105 ( .A1(n_48), .A2(n_106), .B1(n_685), .B2(n_689), .Y(n_105) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_49), .A2(n_90), .B1(n_151), .B2(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g509 ( .A(n_50), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_51), .B(n_127), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_52), .B(n_127), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_53), .B(n_434), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_54), .B(n_215), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_56), .A2(n_60), .B1(n_127), .B2(n_132), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_57), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_58), .B(n_127), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_59), .B(n_127), .Y(n_237) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_62), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_63), .B(n_439), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_64), .A2(n_212), .B(n_215), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_65), .B(n_127), .Y(n_218) );
INVx1_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_67), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_68), .B(n_134), .Y(n_462) );
AO32x2_ASAP7_75t_L g148 ( .A1(n_69), .A2(n_149), .A3(n_155), .B1(n_156), .B2(n_157), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_70), .B(n_135), .Y(n_499) );
INVx1_ASAP7_75t_L g236 ( .A(n_71), .Y(n_236) );
INVx1_ASAP7_75t_L g130 ( .A(n_72), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_73), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_74), .B(n_461), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_75), .A2(n_104), .B1(n_692), .B2(n_701), .C1(n_716), .C2(n_722), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_75), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_76), .A2(n_425), .B(n_427), .C(n_431), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_77), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_78), .B(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_79), .Y(n_523) );
INVx1_ASAP7_75t_L g696 ( .A(n_80), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_81), .B(n_460), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_83), .B(n_151), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_84), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_85), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_87), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_88), .B(n_153), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_89), .B(n_132), .Y(n_225) );
INVx2_ASAP7_75t_L g108 ( .A(n_91), .Y(n_108) );
OR2x2_ASAP7_75t_L g700 ( .A(n_91), .B(n_685), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_92), .A2(n_102), .B1(n_132), .B2(n_133), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_93), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_94), .B(n_434), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_95), .Y(n_459) );
INVxp67_ASAP7_75t_L g526 ( .A(n_96), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_97), .B(n_132), .Y(n_234) );
INVx1_ASAP7_75t_L g428 ( .A(n_98), .Y(n_428) );
INVx1_ASAP7_75t_L g495 ( .A(n_99), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_100), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g511 ( .A(n_101), .B(n_119), .Y(n_511) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp33_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_677), .B1(n_683), .B2(n_684), .Y(n_106) );
INVx1_ASAP7_75t_L g683 ( .A(n_107), .Y(n_683) );
AO22x2_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_109), .B1(n_417), .B2(n_676), .Y(n_107) );
INVx1_ASAP7_75t_L g676 ( .A(n_108), .Y(n_676) );
NOR2x2_ASAP7_75t_L g691 ( .A(n_108), .B(n_685), .Y(n_691) );
INVx1_ASAP7_75t_L g416 ( .A(n_110), .Y(n_416) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_110), .A2(n_416), .B1(n_709), .B2(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_336), .Y(n_110) );
NAND3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_285), .C(n_327), .Y(n_111) );
AOI211xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_190), .B(n_239), .C(n_261), .Y(n_112) );
OAI211xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_145), .B(n_173), .C(n_185), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_115), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g348 ( .A(n_115), .B(n_265), .Y(n_348) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g250 ( .A(n_116), .B(n_176), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_116), .B(n_161), .Y(n_367) );
INVx1_ASAP7_75t_L g385 ( .A(n_116), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_116), .B(n_282), .Y(n_394) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g277 ( .A(n_117), .B(n_161), .Y(n_277) );
AND2x2_ASAP7_75t_L g335 ( .A(n_117), .B(n_282), .Y(n_335) );
INVx1_ASAP7_75t_L g379 ( .A(n_117), .Y(n_379) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g256 ( .A(n_118), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g264 ( .A(n_118), .Y(n_264) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_118), .Y(n_304) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_144), .Y(n_118) );
INVx2_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_119), .A2(n_162), .B(n_172), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_119), .A2(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g478 ( .A(n_119), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_119), .A2(n_506), .B(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_L g158 ( .A(n_120), .B(n_121), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_137), .B(n_142), .Y(n_124) );
O2A1O1Ixp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_130), .B(n_131), .C(n_134), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_127), .Y(n_430) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_128), .Y(n_152) );
AND2x6_ASAP7_75t_L g425 ( .A(n_128), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_129), .Y(n_133) );
INVx1_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
INVx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_134), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_134), .A2(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_134), .B(n_526), .Y(n_525) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g149 ( .A1(n_135), .A2(n_150), .B1(n_153), .B2(n_154), .Y(n_149) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx1_ASAP7_75t_L g426 ( .A(n_136), .Y(n_426) );
AND2x2_ASAP7_75t_L g435 ( .A(n_136), .B(n_216), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g212 ( .A(n_140), .Y(n_212) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g461 ( .A(n_141), .Y(n_461) );
BUFx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_142), .A2(n_163), .B(n_168), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_142), .A2(n_208), .B(n_213), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_142), .A2(n_223), .B(n_226), .Y(n_222) );
INVx4_ASAP7_75t_SL g432 ( .A(n_142), .Y(n_432) );
AND2x4_ASAP7_75t_L g434 ( .A(n_142), .B(n_435), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_142), .B(n_435), .Y(n_496) );
INVxp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_159), .Y(n_146) );
AND2x2_ASAP7_75t_L g243 ( .A(n_147), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g276 ( .A(n_147), .Y(n_276) );
OR2x2_ASAP7_75t_L g402 ( .A(n_147), .B(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_147), .B(n_161), .Y(n_406) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx1_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g265 ( .A(n_148), .B(n_178), .Y(n_265) );
AND2x2_ASAP7_75t_L g305 ( .A(n_148), .B(n_179), .Y(n_305) );
INVx2_ASAP7_75t_L g448 ( .A(n_152), .Y(n_448) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_152), .Y(n_463) );
INVx2_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_153), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_153), .A2(n_182), .B1(n_199), .B2(n_200), .Y(n_198) );
INVx4_ASAP7_75t_L g447 ( .A(n_153), .Y(n_447) );
INVx1_ASAP7_75t_L g475 ( .A(n_155), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_156), .B(n_198), .C(n_201), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_156), .A2(n_232), .B(n_235), .Y(n_231) );
INVx4_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_157), .A2(n_222), .B(n_229), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_157), .A2(n_485), .B(n_486), .Y(n_484) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_157), .Y(n_520) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVxp67_ASAP7_75t_L g347 ( .A(n_159), .Y(n_347) );
AND2x4_ASAP7_75t_L g372 ( .A(n_159), .B(n_265), .Y(n_372) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_160), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g177 ( .A(n_161), .B(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g251 ( .A(n_161), .B(n_179), .Y(n_251) );
INVx1_ASAP7_75t_L g257 ( .A(n_161), .Y(n_257) );
INVx2_ASAP7_75t_L g283 ( .A(n_161), .Y(n_283) );
AND2x2_ASAP7_75t_L g299 ( .A(n_161), .B(n_300), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_166), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .Y(n_168) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_171), .A2(n_214), .B(n_236), .C(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_174), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx2_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
AND2x2_ASAP7_75t_L g362 ( .A(n_176), .B(n_178), .Y(n_362) );
AND2x2_ASAP7_75t_L g279 ( .A(n_177), .B(n_264), .Y(n_279) );
AND2x2_ASAP7_75t_L g378 ( .A(n_177), .B(n_379), .Y(n_378) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_178), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g403 ( .A(n_178), .B(n_264), .Y(n_403) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g189 ( .A(n_179), .Y(n_189) );
AND2x2_ASAP7_75t_L g282 ( .A(n_179), .B(n_283), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_182), .A2(n_214), .B(n_217), .C(n_218), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_182), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g206 ( .A(n_184), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_184), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
AND2x2_ASAP7_75t_L g328 ( .A(n_187), .B(n_263), .Y(n_328) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_188), .B(n_264), .Y(n_313) );
INVx2_ASAP7_75t_L g312 ( .A(n_189), .Y(n_312) );
OAI222xp33_ASAP7_75t_L g316 ( .A1(n_189), .A2(n_256), .B1(n_317), .B2(n_319), .C1(n_320), .C2(n_323), .Y(n_316) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g241 ( .A(n_194), .Y(n_241) );
OR2x2_ASAP7_75t_L g352 ( .A(n_194), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
NOR2x1_ASAP7_75t_L g325 ( .A(n_195), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_195), .B(n_245), .Y(n_331) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
AO21x1_ASAP7_75t_L g291 ( .A1(n_198), .A2(n_201), .B(n_292), .Y(n_291) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_201), .A2(n_423), .B(n_436), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_201), .B(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g439 ( .A(n_201), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_201), .B(n_465), .Y(n_464) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_201), .A2(n_494), .B(n_501), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_202), .A2(n_295), .B1(n_334), .B2(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_220), .Y(n_202) );
INVx3_ASAP7_75t_L g267 ( .A(n_203), .Y(n_267) );
OR2x2_ASAP7_75t_L g400 ( .A(n_203), .B(n_276), .Y(n_400) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g273 ( .A(n_204), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g289 ( .A(n_204), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_204), .B(n_245), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_204), .B(n_221), .Y(n_353) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g244 ( .A(n_205), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g248 ( .A(n_205), .B(n_221), .Y(n_248) );
AND2x2_ASAP7_75t_L g324 ( .A(n_205), .B(n_271), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_205), .B(n_230), .Y(n_364) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_219), .Y(n_205) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_206), .A2(n_231), .B(n_238), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .C(n_212), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_210), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_210), .A2(n_499), .B(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_212), .A2(n_428), .B(n_429), .C(n_430), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_214), .A2(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_220), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g280 ( .A(n_220), .B(n_241), .Y(n_280) );
AND2x2_ASAP7_75t_L g284 ( .A(n_220), .B(n_274), .Y(n_284) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
INVx3_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
AND2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g405 ( .A(n_221), .B(n_388), .Y(n_405) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
INVx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
AND2x2_ASAP7_75t_L g315 ( .A(n_230), .B(n_291), .Y(n_315) );
INVx1_ASAP7_75t_L g358 ( .A(n_230), .Y(n_358) );
OR2x2_ASAP7_75t_L g389 ( .A(n_230), .B(n_291), .Y(n_389) );
AND2x2_ASAP7_75t_L g409 ( .A(n_230), .B(n_245), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_242), .B(n_246), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g247 ( .A(n_241), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_241), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g366 ( .A(n_243), .Y(n_366) );
INVx2_ASAP7_75t_SL g260 ( .A(n_244), .Y(n_260) );
AND2x2_ASAP7_75t_L g380 ( .A(n_244), .B(n_274), .Y(n_380) );
INVx2_ASAP7_75t_L g326 ( .A(n_245), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_245), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B1(n_252), .B2(n_258), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_248), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g414 ( .A(n_248), .Y(n_414) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g339 ( .A(n_250), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_250), .B(n_282), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_251), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g355 ( .A(n_251), .B(n_304), .Y(n_355) );
INVx2_ASAP7_75t_L g411 ( .A(n_251), .Y(n_411) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g281 ( .A(n_254), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_254), .B(n_299), .Y(n_332) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_256), .B(n_276), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g393 ( .A(n_259), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_SL g343 ( .A1(n_260), .A2(n_344), .B(n_346), .C(n_349), .Y(n_343) );
OR2x2_ASAP7_75t_L g370 ( .A(n_260), .B(n_274), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_266), .B1(n_268), .B2(n_275), .C(n_278), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_263), .B(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g361 ( .A(n_263), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
INVx1_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_267), .B(n_322), .Y(n_321) );
INVxp67_ASAP7_75t_L g375 ( .A(n_267), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_267), .B(n_315), .Y(n_391) );
INVx2_ASAP7_75t_L g377 ( .A(n_268), .Y(n_377) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g318 ( .A(n_270), .B(n_289), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_270), .A2(n_286), .B(n_328), .C(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g296 ( .A(n_271), .B(n_291), .Y(n_296) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_275), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g344 ( .A(n_276), .B(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B1(n_281), .B2(n_284), .Y(n_278) );
INVx1_ASAP7_75t_L g398 ( .A(n_280), .Y(n_398) );
INVx1_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
INVx1_ASAP7_75t_L g396 ( .A(n_284), .Y(n_396) );
AOI211xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_289), .B(n_293), .C(n_316), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g359 ( .A(n_289), .Y(n_359) );
AND2x2_ASAP7_75t_L g408 ( .A(n_289), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .B(n_306), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g322 ( .A(n_296), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_296), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g314 ( .A(n_297), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g390 ( .A(n_297), .Y(n_390) );
OAI32xp33_ASAP7_75t_L g401 ( .A1(n_297), .A2(n_349), .A3(n_356), .B1(n_397), .B2(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_299), .B(n_302), .Y(n_298) );
INVx1_ASAP7_75t_SL g369 ( .A(n_299), .Y(n_369) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g309 ( .A(n_305), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B(n_314), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_308), .A2(n_356), .B1(n_382), .B2(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_312), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g342 ( .A(n_326), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_335), .A2(n_377), .B1(n_378), .B2(n_380), .C(n_381), .Y(n_376) );
NAND5xp2_ASAP7_75t_L g336 ( .A(n_337), .B(n_360), .C(n_376), .D(n_386), .E(n_404), .Y(n_336) );
AOI211xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_343), .C(n_350), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g407 ( .A(n_344), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_354), .B2(n_356), .Y(n_350) );
INVx1_ASAP7_75t_SL g383 ( .A(n_353), .Y(n_383) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI322xp33_ASAP7_75t_L g365 ( .A1(n_356), .A2(n_366), .A3(n_367), .B1(n_368), .B2(n_369), .C1(n_370), .C2(n_371), .Y(n_365) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_358), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_358), .B(n_383), .Y(n_382) );
AOI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B(n_365), .C(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_369), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_395) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_394), .B1(n_395), .B2(n_399), .C(n_401), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B(n_391), .C(n_392), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g413 ( .A(n_389), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_407), .B2(n_408), .C(n_410), .Y(n_404) );
AOI21xp33_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B(n_413), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_619), .Y(n_417) );
AND4x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_559), .C(n_574), .D(n_599), .Y(n_418) );
NOR2xp33_ASAP7_75t_SL g419 ( .A(n_420), .B(n_532), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_450), .B(n_512), .Y(n_420) );
AND2x2_ASAP7_75t_L g562 ( .A(n_421), .B(n_467), .Y(n_562) );
AND2x2_ASAP7_75t_L g575 ( .A(n_421), .B(n_466), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_421), .B(n_451), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_421), .Y(n_629) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_438), .Y(n_421) );
INVx2_ASAP7_75t_L g546 ( .A(n_422), .Y(n_546) );
BUFx2_ASAP7_75t_L g573 ( .A(n_422), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_433), .Y(n_423) );
INVx5_ASAP7_75t_L g443 ( .A(n_425), .Y(n_443) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_SL g441 ( .A1(n_432), .A2(n_442), .B(n_443), .C(n_444), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_432), .A2(n_443), .B(n_523), .C(n_524), .Y(n_522) );
BUFx2_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
AND2x2_ASAP7_75t_L g513 ( .A(n_438), .B(n_467), .Y(n_513) );
INVx2_ASAP7_75t_L g529 ( .A(n_438), .Y(n_529) );
AND2x2_ASAP7_75t_L g538 ( .A(n_438), .B(n_466), .Y(n_538) );
AND2x2_ASAP7_75t_L g617 ( .A(n_438), .B(n_546), .Y(n_617) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_449), .Y(n_438) );
INVx2_ASAP7_75t_L g457 ( .A(n_443), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_479), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_451), .B(n_544), .Y(n_582) );
INVx1_ASAP7_75t_L g670 ( .A(n_451), .Y(n_670) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_466), .Y(n_451) );
AND2x2_ASAP7_75t_L g528 ( .A(n_452), .B(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g542 ( .A(n_452), .B(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_452), .Y(n_571) );
OR2x2_ASAP7_75t_L g603 ( .A(n_452), .B(n_545), .Y(n_603) );
AND2x2_ASAP7_75t_L g611 ( .A(n_452), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g644 ( .A(n_452), .B(n_613), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_452), .B(n_513), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_452), .B(n_573), .Y(n_669) );
AND2x2_ASAP7_75t_L g675 ( .A(n_452), .B(n_562), .Y(n_675) );
INVx5_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g535 ( .A(n_453), .Y(n_535) );
AND2x2_ASAP7_75t_L g565 ( .A(n_453), .B(n_545), .Y(n_565) );
AND2x2_ASAP7_75t_L g598 ( .A(n_453), .B(n_558), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_453), .B(n_467), .Y(n_618) );
AND2x2_ASAP7_75t_L g652 ( .A(n_453), .B(n_518), .Y(n_652) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_464), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_462), .C(n_463), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_460), .A2(n_463), .B(n_509), .C(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g558 ( .A(n_466), .B(n_529), .Y(n_558) );
AND2x2_ASAP7_75t_L g569 ( .A(n_466), .B(n_565), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_466), .B(n_545), .Y(n_608) );
INVx2_ASAP7_75t_L g623 ( .A(n_466), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_466), .B(n_557), .Y(n_646) );
AND2x2_ASAP7_75t_L g665 ( .A(n_466), .B(n_617), .Y(n_665) );
INVx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
AND2x2_ASAP7_75t_L g572 ( .A(n_467), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g613 ( .A(n_467), .B(n_529), .Y(n_613) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_476), .Y(n_467) );
AOI21xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_471), .B(n_475), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
AND2x2_ASAP7_75t_L g536 ( .A(n_481), .B(n_519), .Y(n_536) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_482), .B(n_493), .Y(n_516) );
OR2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_519), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_482), .B(n_519), .Y(n_554) );
AND2x2_ASAP7_75t_L g581 ( .A(n_482), .B(n_518), .Y(n_581) );
AND2x2_ASAP7_75t_L g633 ( .A(n_482), .B(n_492), .Y(n_633) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_483), .B(n_503), .Y(n_541) );
AND2x2_ASAP7_75t_L g577 ( .A(n_483), .B(n_493), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_490), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g567 ( .A(n_491), .B(n_549), .Y(n_567) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
OAI322xp33_ASAP7_75t_L g532 ( .A1(n_492), .A2(n_533), .A3(n_537), .B1(n_539), .B2(n_542), .C1(n_547), .C2(n_555), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_492), .B(n_518), .Y(n_540) );
OR2x2_ASAP7_75t_L g550 ( .A(n_492), .B(n_504), .Y(n_550) );
AND2x2_ASAP7_75t_L g552 ( .A(n_492), .B(n_504), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_492), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_492), .B(n_519), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_492), .B(n_648), .Y(n_647) );
INVx5_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_493), .B(n_536), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_503), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g530 ( .A(n_503), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_503), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g592 ( .A(n_503), .B(n_519), .Y(n_592) );
AOI211xp5_ASAP7_75t_SL g620 ( .A1(n_503), .A2(n_621), .B(n_624), .C(n_636), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_503), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g658 ( .A(n_503), .B(n_633), .Y(n_658) );
INVx5_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g586 ( .A(n_504), .B(n_519), .Y(n_586) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_504), .Y(n_595) );
AND2x2_ASAP7_75t_L g635 ( .A(n_504), .B(n_633), .Y(n_635) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_504), .B(n_536), .Y(n_666) );
AND2x2_ASAP7_75t_L g673 ( .A(n_504), .B(n_632), .Y(n_673) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_528), .B2(n_530), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_513), .B(n_535), .Y(n_583) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g531 ( .A(n_516), .Y(n_531) );
OR2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_SL g639 ( .A1(n_516), .A2(n_640), .B1(n_642), .B2(n_643), .C(n_645), .Y(n_639) );
INVx2_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
AND2x2_ASAP7_75t_L g551 ( .A(n_518), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g641 ( .A(n_518), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_518), .B(n_633), .Y(n_654) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVxp67_ASAP7_75t_L g596 ( .A(n_519), .Y(n_596) );
AND2x2_ASAP7_75t_L g632 ( .A(n_519), .B(n_633), .Y(n_632) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_519) );
AND2x2_ASAP7_75t_L g634 ( .A(n_528), .B(n_573), .Y(n_634) );
AND2x2_ASAP7_75t_L g544 ( .A(n_529), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_529), .B(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_531), .B(n_578), .Y(n_615) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g621 ( .A(n_534), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
OR2x2_ASAP7_75t_L g607 ( .A(n_535), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g672 ( .A(n_535), .B(n_617), .Y(n_672) );
INVx2_ASAP7_75t_L g605 ( .A(n_536), .Y(n_605) );
NAND4xp25_ASAP7_75t_SL g668 ( .A(n_537), .B(n_669), .C(n_670), .D(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_538), .B(n_602), .Y(n_637) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_SL g674 ( .A(n_541), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_SL g636 ( .A1(n_542), .A2(n_605), .B(n_609), .C(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g631 ( .A(n_544), .B(n_623), .Y(n_631) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_545), .Y(n_557) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_546), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_550), .B(n_551), .C(n_553), .Y(n_547) );
AND2x2_ASAP7_75t_L g568 ( .A(n_548), .B(n_552), .Y(n_568) );
OAI322xp33_ASAP7_75t_SL g606 ( .A1(n_548), .A2(n_607), .A3(n_609), .B1(n_610), .B2(n_614), .C1(n_615), .C2(n_616), .Y(n_606) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g628 ( .A(n_550), .B(n_554), .Y(n_628) );
INVx1_ASAP7_75t_L g609 ( .A(n_552), .Y(n_609) );
INVx1_ASAP7_75t_SL g627 ( .A(n_554), .Y(n_627) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_566), .B1(n_568), .B2(n_569), .C1(n_570), .C2(n_725), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
OAI322xp33_ASAP7_75t_L g649 ( .A1(n_561), .A2(n_623), .A3(n_628), .B1(n_650), .B2(n_651), .C1(n_653), .C2(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_562), .A2(n_576), .B1(n_600), .B2(n_604), .C(n_606), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g579 ( .A1(n_567), .A2(n_580), .B1(n_582), .B2(n_583), .C1(n_584), .C2(n_587), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_569), .A2(n_576), .B1(n_646), .B2(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_579), .C(n_590), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_576), .A2(n_613), .B(n_656), .C(n_659), .Y(n_655) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g585 ( .A(n_577), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g648 ( .A(n_581), .Y(n_648) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_588), .B(n_613), .Y(n_642) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_597), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_591), .A2(n_660), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_659) );
INVxp33_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_595), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_602), .B(n_613), .Y(n_653) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g664 ( .A(n_617), .B(n_623), .Y(n_664) );
AND4x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_638), .C(n_655), .D(n_667), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI221xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_630) );
INVx1_ASAP7_75t_L g660 ( .A(n_631), .Y(n_660) );
INVx1_ASAP7_75t_SL g650 ( .A(n_635), .Y(n_650) );
NOR2xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_649), .Y(n_638) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_651), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_658), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g684 ( .A(n_677), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx3_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
NAND2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_697), .Y(n_694) );
INVx1_ASAP7_75t_SL g721 ( .A(n_695), .Y(n_721) );
INVx1_ASAP7_75t_L g720 ( .A(n_697), .Y(n_720) );
OA21x2_ASAP7_75t_L g723 ( .A1(n_697), .A2(n_712), .B(n_721), .Y(n_723) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g712 ( .A(n_700), .Y(n_712) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_700), .Y(n_714) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_712), .B(n_713), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
XNOR2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_714), .B(n_715), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
endmodule