module real_jpeg_22078_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_0),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_102),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_102),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_1),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_158),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_158),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_158),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_3),
.A2(n_34),
.B1(n_64),
.B2(n_65),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_22),
.B1(n_64),
.B2(n_65),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_4),
.A2(n_22),
.B1(n_46),
.B2(n_47),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_107),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_107),
.Y(n_247)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_7),
.B(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_130),
.B(n_156),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_9),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_90),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_11),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_282)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_47),
.B(n_60),
.C(n_87),
.D(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_12),
.B(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_12),
.A2(n_108),
.B(n_110),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_12),
.A2(n_31),
.B(n_42),
.C(n_146),
.D(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_12),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_12),
.B(n_35),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_30),
.B(n_32),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_127),
.Y(n_205)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_76),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_74),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_36),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_21),
.A2(n_25),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_23),
.A2(n_27),
.B(n_127),
.C(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_25),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_25),
.B(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_26),
.A2(n_29),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_26),
.A2(n_29),
.B1(n_216),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_26),
.A2(n_207),
.B(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_26),
.A2(n_29),
.B1(n_54),
.B2(n_291),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_29),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_29),
.A2(n_217),
.B(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_35),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_69),
.C(n_71),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_37),
.A2(n_38),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_316),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_50),
.B1(n_167),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_202),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_45),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_42),
.A2(n_45),
.B1(n_244),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_42),
.A2(n_45),
.B1(n_263),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_44),
.Y(n_154)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_46),
.B(n_48),
.Y(n_153)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_47),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_50),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_50),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_50),
.A2(n_168),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_52),
.A2(n_53),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_58),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_58),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_67),
.B1(n_101),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_59),
.A2(n_144),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_59),
.A2(n_67),
.B1(n_199),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_59),
.A2(n_67),
.B1(n_229),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_59),
.A2(n_67),
.B1(n_238),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_60),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_60),
.A2(n_63),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_65),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_64),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_67),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_103),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_68),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_69),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_334),
.B(n_340),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_307),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_342),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_255),
.A3(n_295),
.B1(n_301),
.B2(n_306),
.C(n_343),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_210),
.C(n_251),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_182),
.B(n_209),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_161),
.B(n_181),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_138),
.B(n_160),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_113),
.B(n_137),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_85),
.B(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_108),
.A2(n_121),
.B1(n_157),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_108),
.A2(n_109),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_108),
.A2(n_192),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_108),
.A2(n_121),
.B1(n_227),
.B2(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_108),
.A2(n_121),
.B(n_236),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_117),
.B(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_109),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_124),
.B(n_136),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_127),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B(n_135),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_128),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_151),
.B2(n_159),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_150),
.C(n_159),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_178),
.C(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_176),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_170),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_195),
.C(n_196),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_191),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_211),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_231),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_231),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_230),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_230),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_228),
.Y(n_240)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_249),
.B2(n_250),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_239),
.C(n_250),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_237),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_273),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_256),
.B(n_273),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.C(n_272),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_257),
.A2(n_258),
.B1(n_266),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_268),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_286),
.B(n_290),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_269),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_293),
.B2(n_294),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_284),
.B2(n_285),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_285),
.C(n_294),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_281),
.B(n_283),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_281),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_283),
.A2(n_309),
.B1(n_318),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_292),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_288),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_320),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_320),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_318),
.C(n_319),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_311),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_316),
.C(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_322),
.C(n_326),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_314),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);


endmodule