module fake_netlist_6_872_n_804 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_804);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_804;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_60),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_49),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_28),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_23),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_81),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_16),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_36),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_80),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_41),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_25),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_9),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_21),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_18),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_40),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_27),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_26),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_37),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_57),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_87),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_61),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_31),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_70),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_39),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_65),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_0),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_163),
.A2(n_83),
.B(n_156),
.Y(n_220)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_202),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_165),
.B(n_173),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_161),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_0),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_1),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_175),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_2),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_3),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_169),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_170),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_224),
.B(n_191),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_224),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_167),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_210),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_224),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_171),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_224),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_233),
.B(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_233),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_180),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_182),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_192),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_223),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_235),
.Y(n_292)
);

AO21x2_ASAP7_75t_L g293 ( 
.A1(n_218),
.A2(n_197),
.B(n_195),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

CKINVDCx6p67_ASAP7_75t_R g296 ( 
.A(n_233),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_233),
.B(n_208),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_200),
.Y(n_302)
);

AND3x2_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_212),
.C(n_211),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_216),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_238),
.A2(n_212),
.B1(n_211),
.B2(n_208),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_257),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_245),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_265),
.B(n_241),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_257),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_258),
.C(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_279),
.B(n_245),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_257),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_244),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_237),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_298),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_255),
.B1(n_247),
.B2(n_241),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_237),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_305),
.A2(n_250),
.B1(n_254),
.B2(n_252),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_237),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_266),
.B1(n_293),
.B2(n_285),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_227),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_267),
.B(n_237),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_267),
.B(n_201),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_222),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_275),
.B(n_243),
.Y(n_336)
);

BUFx2_ASAP7_75t_R g337 ( 
.A(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_293),
.B(n_243),
.Y(n_339)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_228),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_229),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_248),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_301),
.B(n_246),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_277),
.B(n_204),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_277),
.B(n_249),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_206),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_281),
.B(n_252),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_222),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_260),
.B(n_253),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_263),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_263),
.B(n_253),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_295),
.B(n_209),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_292),
.A2(n_254),
.B1(n_235),
.B2(n_242),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_296),
.B(n_221),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_272),
.B(n_256),
.Y(n_363)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_221),
.C(n_232),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_295),
.B(n_256),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_300),
.B(n_256),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_280),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_256),
.B1(n_242),
.B2(n_239),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_300),
.B(n_232),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_280),
.B(n_232),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_278),
.B(n_288),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_312),
.A2(n_291),
.B(n_306),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_239),
.Y(n_374)
);

OAI321xp33_ASAP7_75t_L g375 ( 
.A1(n_329),
.A2(n_239),
.A3(n_242),
.B1(n_306),
.B2(n_307),
.C(n_274),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_327),
.B(n_307),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_220),
.B(n_264),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_264),
.Y(n_378)
);

AOI33xp33_ASAP7_75t_L g379 ( 
.A1(n_329),
.A2(n_274),
.A3(n_283),
.B1(n_287),
.B2(n_264),
.B3(n_269),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_312),
.A2(n_309),
.B(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_269),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_319),
.A2(n_269),
.B(n_270),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_327),
.B(n_291),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_331),
.A2(n_270),
.B(n_274),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_283),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_287),
.B1(n_283),
.B2(n_270),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_3),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_330),
.B(n_287),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_326),
.A2(n_288),
.B(n_278),
.C(n_291),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_336),
.A2(n_278),
.B(n_288),
.C(n_6),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_336),
.A2(n_291),
.B(n_271),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_288),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_271),
.B(n_5),
.C(n_6),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_352),
.A2(n_271),
.B(n_86),
.Y(n_399)
);

AO21x1_ASAP7_75t_L g400 ( 
.A1(n_320),
.A2(n_4),
.B(n_5),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_335),
.B(n_342),
.Y(n_401)
);

NOR2x1_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_271),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_316),
.B(n_271),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_353),
.B(n_7),
.Y(n_404)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_361),
.B(n_7),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_311),
.B(n_348),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_340),
.A2(n_92),
.B(n_153),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_91),
.B(n_151),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_324),
.B(n_22),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_24),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_349),
.B(n_8),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_323),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_334),
.B(n_10),
.Y(n_415)
);

BUFx12f_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_29),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_30),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_337),
.A2(n_97),
.B1(n_149),
.B2(n_148),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_340),
.A2(n_94),
.B(n_147),
.Y(n_420)
);

AOI21xp33_ASAP7_75t_L g421 ( 
.A1(n_346),
.A2(n_11),
.B(n_12),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_317),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_340),
.A2(n_93),
.B(n_145),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_359),
.B(n_33),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_333),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_343),
.A2(n_98),
.B(n_143),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_345),
.A2(n_85),
.B(n_142),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_328),
.B(n_35),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_355),
.A2(n_84),
.B(n_141),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_368),
.B(n_358),
.Y(n_430)
);

OAI21xp33_ASAP7_75t_L g431 ( 
.A1(n_341),
.A2(n_12),
.B(n_13),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_357),
.A2(n_99),
.B(n_139),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_13),
.Y(n_433)
);

O2A1O1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_369),
.A2(n_366),
.B(n_365),
.C(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_38),
.Y(n_435)
);

CKINVDCx11_ASAP7_75t_R g436 ( 
.A(n_371),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_351),
.B(n_14),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_363),
.A2(n_100),
.B(n_138),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_365),
.A2(n_82),
.B(n_137),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_42),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_14),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_377),
.A2(n_394),
.B(n_373),
.Y(n_442)
);

AOI31xp33_ASAP7_75t_L g443 ( 
.A1(n_419),
.A2(n_369),
.A3(n_366),
.B(n_17),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_15),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_317),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_377),
.A2(n_434),
.B(n_403),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_317),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_382),
.A2(n_317),
.B(n_102),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_380),
.B(n_101),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_379),
.B(n_77),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_390),
.B(n_103),
.Y(n_451)
);

OAI21x1_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_76),
.B(n_136),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_416),
.Y(n_453)
);

AOI221x1_ASAP7_75t_L g454 ( 
.A1(n_389),
.A2(n_75),
.B1(n_135),
.B2(n_134),
.C(n_133),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_382),
.A2(n_157),
.B(n_72),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_395),
.Y(n_456)
);

NAND2x1_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_71),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_378),
.A2(n_73),
.B(n_131),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_396),
.A2(n_69),
.B(n_128),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_407),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_405),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_391),
.A2(n_435),
.B(n_428),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_381),
.A2(n_376),
.B(n_422),
.Y(n_465)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_422),
.A2(n_384),
.B(n_401),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_374),
.B(n_19),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_19),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_105),
.B(n_126),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_385),
.B(n_104),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_392),
.A2(n_68),
.B(n_125),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_425),
.B(n_20),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_386),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_106),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_412),
.A2(n_21),
.B1(n_43),
.B2(n_44),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_397),
.B(n_45),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_431),
.A2(n_46),
.B(n_47),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_409),
.A2(n_132),
.B(n_50),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_375),
.A2(n_48),
.B(n_51),
.Y(n_486)
);

OAI21x1_ASAP7_75t_SL g487 ( 
.A1(n_426),
.A2(n_52),
.B(n_53),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_440),
.A2(n_124),
.B(n_56),
.Y(n_490)
);

AOI221x1_ASAP7_75t_L g491 ( 
.A1(n_398),
.A2(n_54),
.B1(n_58),
.B2(n_63),
.C(n_66),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_375),
.A2(n_393),
.B(n_399),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_421),
.B(n_67),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_417),
.A2(n_107),
.B(n_109),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_418),
.A2(n_110),
.B(n_111),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_113),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_424),
.A2(n_114),
.B(n_115),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_406),
.B(n_116),
.Y(n_498)
);

AO31x2_ASAP7_75t_L g499 ( 
.A1(n_441),
.A2(n_117),
.A3(n_118),
.B(n_120),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_448),
.A2(n_442),
.B(n_446),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_472),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_423),
.B1(n_420),
.B2(n_408),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_456),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_458),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_471),
.A2(n_427),
.B(n_438),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_413),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_463),
.A2(n_429),
.B(n_432),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_439),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_475),
.B(n_123),
.Y(n_509)
);

OAI21x1_ASAP7_75t_SL g510 ( 
.A1(n_486),
.A2(n_452),
.B(n_487),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_485),
.A2(n_121),
.B(n_122),
.Y(n_511)
);

BUFx4_ASAP7_75t_SL g512 ( 
.A(n_464),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_455),
.A2(n_449),
.B(n_473),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_444),
.B(n_476),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_471),
.A2(n_492),
.B(n_449),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_461),
.A2(n_475),
.B1(n_480),
.B2(n_469),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_462),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_466),
.B(n_443),
.C(n_498),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_461),
.B(n_478),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_460),
.A2(n_490),
.B(n_465),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

INVx4_ASAP7_75t_SL g522 ( 
.A(n_461),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_492),
.A2(n_450),
.B(n_491),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_474),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_453),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_477),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_459),
.A2(n_467),
.B(n_450),
.Y(n_528)
);

BUFx2_ASAP7_75t_SL g529 ( 
.A(n_479),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_468),
.A2(n_494),
.B(n_486),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_494),
.A2(n_451),
.B(n_470),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_495),
.A2(n_483),
.B(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_489),
.A2(n_497),
.B(n_496),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_493),
.B(n_481),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_484),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_454),
.A2(n_481),
.B(n_499),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_499),
.B(n_390),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_472),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_458),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_448),
.A2(n_442),
.B(n_377),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_458),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_448),
.A2(n_442),
.B(n_377),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_471),
.A2(n_385),
.B(n_377),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_488),
.B(n_383),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_518),
.A2(n_539),
.B1(n_527),
.B2(n_514),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_527),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_547),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_519),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_523),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_514),
.A2(n_537),
.B1(n_539),
.B2(n_551),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_528),
.A2(n_500),
.B(n_513),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_546),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_546),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_548),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_501),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_500),
.Y(n_569)
);

AOI21x1_ASAP7_75t_L g570 ( 
.A1(n_528),
.A2(n_513),
.B(n_549),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_539),
.A2(n_542),
.B1(n_510),
.B2(n_531),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_524),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_545),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_548),
.Y(n_576)
);

BUFx2_ASAP7_75t_R g577 ( 
.A(n_525),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_548),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_522),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_548),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_530),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_506),
.B(n_539),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_535),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_530),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_543),
.Y(n_588)
);

OAI222xp33_ASAP7_75t_L g589 ( 
.A1(n_516),
.A2(n_542),
.B1(n_502),
.B2(n_509),
.C1(n_525),
.C2(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_530),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_531),
.A2(n_533),
.B1(n_508),
.B2(n_529),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_520),
.A2(n_549),
.B(n_507),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_531),
.B(n_508),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_550),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_520),
.A2(n_507),
.B(n_534),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_553),
.A2(n_515),
.B1(n_533),
.B2(n_540),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_583),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_554),
.B(n_517),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_554),
.B(n_517),
.Y(n_601)
);

AO31x2_ASAP7_75t_L g602 ( 
.A1(n_595),
.A2(n_540),
.A3(n_541),
.B(n_515),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_562),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_573),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_556),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_568),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_543),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_556),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_568),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_583),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_572),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_561),
.A2(n_508),
.B1(n_521),
.B2(n_509),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_566),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_559),
.Y(n_616)
);

NAND2x1_ASAP7_75t_L g617 ( 
.A(n_567),
.B(n_544),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_559),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_558),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_521),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_564),
.B(n_515),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_561),
.B(n_544),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_583),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_585),
.B(n_550),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_564),
.B(n_536),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_565),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_565),
.B(n_536),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_585),
.B(n_505),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_557),
.B(n_590),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_576),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_589),
.B(n_505),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_594),
.B(n_511),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_511),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_594),
.B(n_534),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_595),
.A2(n_512),
.A3(n_569),
.B(n_574),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_576),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_576),
.A2(n_567),
.B1(n_578),
.B2(n_591),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_586),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_590),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_586),
.B(n_571),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_575),
.A2(n_579),
.B1(n_582),
.B2(n_581),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_619),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_552),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_621),
.B(n_552),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_630),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_604),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_578),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_606),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_620),
.B(n_592),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_641),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_607),
.B(n_581),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_641),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_SL g657 ( 
.A1(n_632),
.A2(n_576),
.B1(n_578),
.B2(n_567),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_636),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_599),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_629),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_613),
.A2(n_577),
.B1(n_582),
.B2(n_575),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_624),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_633),
.B(n_560),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_635),
.B(n_587),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_600),
.B(n_579),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_633),
.B(n_560),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_625),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_625),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_632),
.A2(n_580),
.B1(n_576),
.B2(n_567),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_619),
.B(n_574),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_622),
.A2(n_580),
.B1(n_578),
.B2(n_574),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_631),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_605),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_608),
.B(n_587),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_597),
.B(n_587),
.C(n_569),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_628),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_612),
.B(n_569),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_634),
.B(n_570),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_637),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_631),
.B(n_570),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_615),
.B(n_563),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_644),
.B(n_593),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_663),
.B(n_602),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_682),
.B(n_634),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_679),
.B(n_651),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_659),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_652),
.B(n_601),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_663),
.B(n_602),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_658),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_658),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_683),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_664),
.B(n_602),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_664),
.B(n_602),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_R g697 ( 
.A(n_665),
.B(n_639),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_650),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_646),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_667),
.B(n_597),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_673),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_666),
.B(n_637),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_683),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_670),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_667),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_666),
.B(n_637),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_649),
.B(n_618),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_678),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_667),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_678),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_654),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_674),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_655),
.B(n_616),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_661),
.A2(n_634),
.B1(n_623),
.B2(n_609),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_679),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_653),
.B(n_651),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_647),
.B(n_637),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_717),
.A2(n_675),
.B1(n_662),
.B2(n_660),
.C(n_677),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_708),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_715),
.A2(n_681),
.B1(n_657),
.B2(n_669),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_686),
.Y(n_723)
);

NAND2x1_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_679),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_698),
.B(n_662),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_691),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_687),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_716),
.B(n_679),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_687),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_705),
.B(n_684),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_SL g731 ( 
.A(n_699),
.B(n_672),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_692),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_716),
.B(n_648),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_706),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_702),
.B(n_648),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_693),
.B(n_684),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_714),
.B(n_660),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_729),
.B(n_718),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_721),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_726),
.Y(n_741)
);

OAI31xp33_ASAP7_75t_L g742 ( 
.A1(n_720),
.A2(n_689),
.A3(n_675),
.B(n_686),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_720),
.Y(n_743)
);

AOI221xp5_ASAP7_75t_L g744 ( 
.A1(n_719),
.A2(n_693),
.B1(n_704),
.B2(n_711),
.C(n_709),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_732),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_725),
.A2(n_643),
.B(n_672),
.C(n_703),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_734),
.Y(n_747)
);

AOI21xp33_ASAP7_75t_L g748 ( 
.A1(n_731),
.A2(n_697),
.B(n_700),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_735),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_733),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_735),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_723),
.A2(n_718),
.B1(n_702),
.B2(n_707),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_742),
.A2(n_724),
.B1(n_722),
.B2(n_738),
.C(n_723),
.Y(n_753)
);

AO22x1_ASAP7_75t_L g754 ( 
.A1(n_743),
.A2(n_727),
.B1(n_723),
.B2(n_728),
.Y(n_754)
);

OAI322xp33_ASAP7_75t_L g755 ( 
.A1(n_743),
.A2(n_737),
.A3(n_730),
.B1(n_713),
.B2(n_695),
.C1(n_694),
.C2(n_700),
.Y(n_755)
);

OAI31xp33_ASAP7_75t_L g756 ( 
.A1(n_748),
.A2(n_727),
.A3(n_728),
.B(n_686),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_746),
.A2(n_744),
.B(n_752),
.C(n_727),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_745),
.B(n_736),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_750),
.B(n_733),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_758),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_759),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_740),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_753),
.B(n_672),
.Y(n_763)
);

NOR4xp25_ASAP7_75t_L g764 ( 
.A(n_755),
.B(n_741),
.C(n_747),
.D(n_749),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_754),
.B(n_739),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_751),
.Y(n_766)
);

OAI211xp5_ASAP7_75t_SL g767 ( 
.A1(n_760),
.A2(n_756),
.B(n_752),
.C(n_671),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_764),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_763),
.A2(n_696),
.B(n_688),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_769),
.B(n_765),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_766),
.B(n_765),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_770),
.A2(n_701),
.B(n_696),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_772),
.B(n_768),
.Y(n_774)
);

OAI322xp33_ASAP7_75t_L g775 ( 
.A1(n_771),
.A2(n_767),
.A3(n_694),
.B1(n_695),
.B2(n_680),
.C1(n_713),
.C2(n_706),
.Y(n_775)
);

NAND4xp75_ASAP7_75t_L g776 ( 
.A(n_773),
.B(n_610),
.C(n_598),
.D(n_645),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_774),
.B(n_736),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_776),
.B(n_707),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_775),
.Y(n_779)
);

NOR2x1_ASAP7_75t_L g780 ( 
.A(n_774),
.B(n_627),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_774),
.A2(n_701),
.B1(n_710),
.B2(n_712),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_780),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_777),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_778),
.B(n_710),
.Y(n_784)
);

AOI31xp33_ASAP7_75t_L g785 ( 
.A1(n_779),
.A2(n_610),
.A3(n_598),
.B(n_640),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_781),
.B(n_712),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_779),
.A2(n_617),
.B1(n_682),
.B2(n_642),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_782),
.Y(n_788)
);

OAI22x1_ASAP7_75t_L g789 ( 
.A1(n_783),
.A2(n_682),
.B1(n_642),
.B2(n_639),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_785),
.A2(n_784),
.B(n_787),
.Y(n_790)
);

AOI31xp33_ASAP7_75t_L g791 ( 
.A1(n_786),
.A2(n_680),
.A3(n_614),
.B(n_603),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_790),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_SL g793 ( 
.A1(n_788),
.A2(n_639),
.B(n_638),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_790),
.A2(n_682),
.B1(n_638),
.B2(n_677),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_789),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_792),
.A2(n_791),
.B(n_603),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_795),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_794),
.A2(n_690),
.B1(n_685),
.B2(n_676),
.Y(n_798)
);

OAI31xp33_ASAP7_75t_L g799 ( 
.A1(n_797),
.A2(n_793),
.A3(n_656),
.B(n_654),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_798),
.B(n_685),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_799),
.A2(n_796),
.B(n_596),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_801),
.A2(n_800),
.B(n_626),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_802),
.B(n_614),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_803),
.A2(n_611),
.B1(n_626),
.B2(n_668),
.Y(n_804)
);


endmodule