module fake_jpeg_29680_n_97 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_39),
.C(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_51),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_19),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_56),
.B1(n_6),
.B2(n_7),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_3),
.B(n_4),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_6),
.Y(n_64)
);

BUFx2_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_48),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_10),
.C(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_9),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_23),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_26),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_17),
.C(n_21),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_69),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_90),
.A3(n_79),
.B1(n_76),
.B2(n_61),
.C1(n_82),
.C2(n_59),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_82),
.B(n_81),
.C(n_79),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_87),
.Y(n_97)
);


endmodule