module fake_jpeg_16171_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_0),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_16),
.B(n_19),
.C(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_3),
.B1(n_11),
.B2(n_6),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_5),
.B(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_48),
.B(n_23),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_46),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_23),
.B1(n_14),
.B2(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_16),
.B1(n_19),
.B2(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_26),
.A2(n_24),
.B(n_22),
.C(n_14),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_20),
.B(n_7),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_64),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_50),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_5),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_68),
.C(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_78),
.B1(n_54),
.B2(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_75),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_85),
.C(n_89),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_86),
.B(n_67),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_66),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_64),
.B(n_77),
.C(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_90),
.B1(n_78),
.B2(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_95),
.C(n_96),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_58),
.B1(n_43),
.B2(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_87),
.B1(n_86),
.B2(n_83),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_56),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_86),
.B1(n_81),
.B2(n_67),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_94),
.B1(n_31),
.B2(n_34),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_96),
.C(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_105),
.C(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_95),
.C(n_94),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_101),
.B(n_9),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_20),
.B(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_8),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_20),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_108),
.Y(n_113)
);


endmodule