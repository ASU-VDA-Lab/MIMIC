module fake_netlist_6_15_n_1812 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1812);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1812;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_12),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_54),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_21),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_70),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_58),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_57),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_12),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_42),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_15),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_20),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_23),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_28),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_118),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_2),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_34),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_19),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_82),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_56),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_86),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_68),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_34),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_84),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_91),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_15),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_100),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_24),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_130),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_40),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_121),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_115),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_73),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_25),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_71),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_110),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_53),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_67),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_3),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_85),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_122),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_62),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_40),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_113),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_42),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_87),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_75),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_95),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_38),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_36),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_127),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_21),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_29),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_43),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_18),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_7),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_64),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_101),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_30),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_99),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_14),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_63),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_47),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_117),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_123),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_145),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_4),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_88),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_148),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_6),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_44),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_173),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_160),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_173),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_251),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_250),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_164),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_173),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_165),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_173),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_155),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_173),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_173),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_185),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_213),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_173),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_262),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_166),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_262),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_156),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_233),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_232),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_187),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_167),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_248),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_232),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_208),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_168),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_234),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_189),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_208),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_220),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_276),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_236),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_260),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_258),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_175),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_157),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_224),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_182),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_224),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_183),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_193),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_197),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_198),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_161),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_286),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_180),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_180),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_186),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_186),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_286),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_311),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_276),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_317),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_199),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_339),
.B(n_287),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_204),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_373),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_322),
.B(n_169),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_321),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_312),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_314),
.A2(n_162),
.B(n_154),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_320),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_322),
.B(n_189),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_338),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_319),
.A2(n_163),
.B1(n_270),
.B2(n_297),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_205),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_318),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_346),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_318),
.B(n_287),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_323),
.A2(n_162),
.B(n_154),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_R g419 ( 
.A(n_350),
.B(n_206),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_357),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_316),
.A2(n_230),
.B1(n_188),
.B2(n_306),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_325),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_362),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_337),
.B(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_326),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_313),
.B(n_176),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_330),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_341),
.B(n_177),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_364),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_215),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_398),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_386),
.B(n_313),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_366),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_408),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_395),
.Y(n_455)
);

AND3x2_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_352),
.C(n_192),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_400),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_328),
.C(n_327),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_406),
.B(n_192),
.C(n_177),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_398),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_427),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_431),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_194),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

AOI22x1_ASAP7_75t_L g481 ( 
.A1(n_382),
.A2(n_379),
.B1(n_378),
.B2(n_377),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_405),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_381),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_401),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_391),
.B(n_368),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_408),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_435),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_428),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_394),
.B(n_324),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_386),
.B(n_363),
.Y(n_494)
);

BUFx6f_ASAP7_75t_SL g495 ( 
.A(n_386),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_383),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_410),
.B(n_315),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_394),
.B(n_369),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_397),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_424),
.A2(n_316),
.B1(n_358),
.B2(n_363),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_370),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_414),
.B(n_342),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_417),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

AND3x1_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_216),
.C(n_203),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_390),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_385),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_443),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_389),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_386),
.B(n_358),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_386),
.B(n_375),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_389),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_434),
.A2(n_371),
.B1(n_243),
.B2(n_280),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_393),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_393),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_382),
.B(n_375),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_382),
.B(n_380),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_345),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_380),
.A2(n_229),
.B1(n_275),
.B2(n_273),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_423),
.B(n_436),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_419),
.B(n_375),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

NAND3xp33_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_200),
.C(n_194),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_387),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_444),
.B(n_202),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_444),
.B(n_294),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_405),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_416),
.B(n_203),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_399),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_403),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_412),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_434),
.A2(n_256),
.B1(n_211),
.B2(n_308),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_392),
.B(n_200),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_403),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_404),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_439),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_412),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_404),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_410),
.B(n_329),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_412),
.B(n_303),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_406),
.A2(n_229),
.B1(n_216),
.B2(n_247),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_418),
.A2(n_210),
.B(n_201),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_401),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_419),
.B(n_176),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_412),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_412),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_409),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_409),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_422),
.A2(n_222),
.B1(n_212),
.B2(n_210),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_411),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_412),
.B(n_218),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_440),
.Y(n_584)
);

INVxp33_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_412),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_438),
.B(n_345),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_440),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_415),
.B(n_430),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_415),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_387),
.B(n_352),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_454),
.Y(n_593)
);

BUFx6f_ASAP7_75t_SL g594 ( 
.A(n_461),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_499),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_413),
.C(n_422),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_396),
.C(n_384),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_540),
.A2(n_421),
.B1(n_426),
.B2(n_360),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_490),
.B(n_421),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_542),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_493),
.B(n_415),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_554),
.B(n_415),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_544),
.B(n_426),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_544),
.B(n_424),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_343),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_544),
.B(n_424),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_499),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_516),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_555),
.B(n_415),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_452),
.B(n_415),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_495),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_511),
.B(n_424),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_480),
.B(n_347),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_509),
.B(n_415),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_557),
.B(n_158),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_539),
.B(n_418),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_532),
.B(n_476),
.Y(n_617)
);

OAI221xp5_ASAP7_75t_L g618 ( 
.A1(n_543),
.A2(n_295),
.B1(n_261),
.B2(n_266),
.C(n_271),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_542),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_587),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_476),
.B(n_418),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_503),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_247),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_476),
.B(n_418),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_476),
.A2(n_418),
.B1(n_417),
.B2(n_392),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_503),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_528),
.B(n_170),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_507),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_497),
.B(n_392),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_507),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_558),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_497),
.B(n_392),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_558),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_488),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_462),
.A2(n_273),
.B(n_261),
.C(n_266),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_480),
.B(n_384),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_498),
.B(n_392),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_592),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_590),
.B(n_221),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_507),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_462),
.B(n_223),
.Y(n_643)
);

BUFx5_ASAP7_75t_L g644 ( 
.A(n_500),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_566),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_548),
.B(n_571),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_515),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_566),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_506),
.B(n_396),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_504),
.B(n_417),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_569),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_548),
.B(n_225),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_548),
.B(n_226),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_569),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_518),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_510),
.B(n_417),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_510),
.B(n_417),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_578),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_513),
.B(n_519),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_489),
.A2(n_228),
.B1(n_252),
.B2(n_305),
.Y(n_663)
);

INVxp33_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_513),
.B(n_417),
.Y(n_665)
);

AND2x4_ASAP7_75t_SL g666 ( 
.A(n_461),
.B(n_176),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_502),
.A2(n_235),
.B1(n_237),
.B2(n_239),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_578),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_429),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_534),
.B(n_171),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_492),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_572),
.A2(n_263),
.B1(n_201),
.B2(n_212),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_523),
.B(n_240),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_523),
.B(n_429),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_449),
.A2(n_265),
.B1(n_227),
.B2(n_231),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_567),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_494),
.A2(n_265),
.B1(n_227),
.B2(n_231),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_524),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_484),
.B(n_222),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_525),
.B(n_242),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_241),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_580),
.A2(n_550),
.B(n_463),
.C(n_579),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_526),
.B(n_529),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_581),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_522),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_524),
.B(n_430),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_574),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_547),
.B(n_172),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_526),
.B(n_241),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_529),
.B(n_253),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_535),
.B(n_253),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_564),
.B(n_437),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_535),
.B(n_255),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_470),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_541),
.B(n_255),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_531),
.A2(n_281),
.B1(n_244),
.B2(n_249),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_541),
.B(n_257),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_557),
.A2(n_283),
.B1(n_279),
.B2(n_299),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_549),
.B(n_257),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_581),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_551),
.B(n_492),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_580),
.A2(n_271),
.B1(n_304),
.B2(n_295),
.C(n_275),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_549),
.B(n_552),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_508),
.B(n_288),
.C(n_184),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_583),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_552),
.B(n_553),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_564),
.B(n_437),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_463),
.A2(n_442),
.B(n_441),
.C(n_306),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_530),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_553),
.B(n_583),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_550),
.A2(n_263),
.B1(n_292),
.B2(n_293),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_461),
.B(n_441),
.Y(n_714)
);

NAND2x1_ASAP7_75t_L g715 ( 
.A(n_453),
.B(n_442),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_545),
.B(n_292),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_530),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_576),
.B(n_300),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_576),
.B(n_293),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_481),
.A2(n_304),
.B1(n_181),
.B2(n_214),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_533),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_575),
.B(n_179),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_537),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_195),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_564),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_456),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_501),
.B(n_196),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_570),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_481),
.B(n_207),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_378),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_538),
.B(n_559),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_585),
.A2(n_379),
.B(n_367),
.C(n_365),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_538),
.A2(n_559),
.B(n_560),
.C(n_565),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_560),
.B(n_209),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_565),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_584),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_584),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_588),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_576),
.B(n_176),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_564),
.A2(n_181),
.B1(n_214),
.B2(n_282),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_591),
.B(n_181),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_495),
.A2(n_181),
.B1(n_214),
.B2(n_278),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_591),
.B(n_214),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_588),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_589),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_589),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_517),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_446),
.B(n_217),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_461),
.B(n_367),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_445),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_446),
.B(n_219),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_564),
.A2(n_285),
.B1(n_245),
.B2(n_246),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_446),
.B(n_238),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_447),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_582),
.A2(n_290),
.B1(n_264),
.B2(n_267),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_447),
.B(n_259),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_445),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_586),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_445),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_451),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_678),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_601),
.B(n_451),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_595),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_617),
.B(n_467),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_595),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_632),
.B(n_459),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_607),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_607),
.Y(n_770)
);

AO22x1_ASAP7_75t_L g771 ( 
.A1(n_596),
.A2(n_458),
.B1(n_460),
.B2(n_505),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_657),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_599),
.B(n_467),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_622),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_598),
.B(n_562),
.C(n_268),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_621),
.B(n_586),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_SL g777 ( 
.A(n_670),
.B(n_284),
.C(n_272),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_694),
.B(n_517),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_622),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_459),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_678),
.Y(n_782)
);

AND3x2_ASAP7_75t_SL g783 ( 
.A(n_670),
.B(n_9),
.C(n_13),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_676),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_647),
.Y(n_785)
);

NAND2x1_ASAP7_75t_L g786 ( 
.A(n_759),
.B(n_751),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_611),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_704),
.A2(n_472),
.B1(n_477),
.B2(n_471),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_645),
.B(n_466),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_627),
.Y(n_790)
);

OAI21xp33_ASAP7_75t_L g791 ( 
.A1(n_664),
.A2(n_289),
.B(n_277),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_634),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_671),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_603),
.A2(n_586),
.B1(n_446),
.B2(n_568),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_610),
.B(n_467),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_703),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_694),
.B(n_448),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_631),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_467),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_614),
.B(n_448),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_644),
.B(n_448),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_625),
.B(n_448),
.Y(n_803)
);

CKINVDCx8_ASAP7_75t_R g804 ( 
.A(n_636),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_648),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_644),
.B(n_464),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_648),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_649),
.B(n_466),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_652),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_653),
.B(n_469),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_686),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_686),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_694),
.B(n_464),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_656),
.B(n_469),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_661),
.B(n_471),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_668),
.B(n_472),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_652),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_687),
.B(n_349),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_679),
.B(n_477),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_594),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_685),
.B(n_485),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_605),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_631),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_693),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_593),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_600),
.A2(n_269),
.B1(n_307),
.B2(n_296),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_693),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_631),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_711),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_702),
.B(n_485),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_707),
.B(n_486),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_711),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_720),
.Y(n_833)
);

NOR2x1p5_ASAP7_75t_L g834 ( 
.A(n_638),
.B(n_298),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_748),
.B(n_464),
.Y(n_835)
);

NOR2x2_ASAP7_75t_L g836 ( 
.A(n_623),
.B(n_301),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_619),
.B(n_486),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_720),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_736),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_650),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_603),
.A2(n_512),
.B1(n_473),
.B2(n_568),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_620),
.A2(n_487),
.B1(n_465),
.B2(n_468),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_624),
.B(n_487),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_631),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_736),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_642),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_644),
.B(n_464),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_473),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_628),
.B(n_473),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_628),
.B(n_473),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_642),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_594),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_751),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_758),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_758),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_672),
.A2(n_713),
.B1(n_618),
.B2(n_616),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_717),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_722),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_642),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_714),
.B(n_482),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_644),
.B(n_482),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_757),
.B(n_602),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_688),
.B(n_349),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_728),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_673),
.A2(n_520),
.B1(n_521),
.B2(n_568),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_724),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_755),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_608),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_626),
.A2(n_479),
.B1(n_496),
.B2(n_457),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_611),
.B(n_354),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_643),
.A2(n_479),
.B1(n_496),
.B2(n_457),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_609),
.A2(n_453),
.B(n_577),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_757),
.B(n_482),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_643),
.A2(n_465),
.B1(n_468),
.B2(n_474),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_SL g877 ( 
.A(n_728),
.B(n_302),
.C(n_354),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_669),
.B(n_674),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_761),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_613),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_709),
.B(n_482),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_760),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_732),
.Y(n_884)
);

AND3x1_ASAP7_75t_SL g885 ( 
.A(n_689),
.B(n_355),
.C(n_361),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_629),
.B(n_712),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_644),
.B(n_512),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_727),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_709),
.B(n_512),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_611),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_660),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_729),
.A2(n_355),
.B1(n_361),
.B2(n_365),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_760),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_644),
.B(n_512),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_684),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_735),
.B(n_723),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_689),
.B(n_474),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_723),
.B(n_520),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_683),
.A2(n_573),
.B(n_455),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_705),
.Y(n_900)
);

AND3x2_ASAP7_75t_SL g901 ( 
.A(n_741),
.B(n_14),
.C(n_17),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_708),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_666),
.B(n_475),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_637),
.B(n_520),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_726),
.B(n_623),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_737),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_662),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_698),
.B(n_573),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_660),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_637),
.B(n_521),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_739),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_730),
.A2(n_491),
.B1(n_475),
.B2(n_455),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_725),
.B(n_521),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_700),
.B(n_491),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_660),
.Y(n_915)
);

O2A1O1Ixp5_ASAP7_75t_L g916 ( 
.A1(n_716),
.A2(n_455),
.B(n_561),
.C(n_556),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_739),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

AND2x4_ASAP7_75t_SL g919 ( 
.A(n_623),
.B(n_597),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_747),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_630),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_731),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_612),
.B(n_561),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_738),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_696),
.B(n_556),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_680),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_666),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_662),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_680),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_721),
.A2(n_556),
.B1(n_577),
.B2(n_536),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_746),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_749),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_604),
.A2(n_606),
.B1(n_675),
.B2(n_706),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_633),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_752),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_715),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_R g938 ( 
.A(n_615),
.B(n_79),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_651),
.B(n_577),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_673),
.B(n_681),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_658),
.B(n_577),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_639),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_681),
.B(n_536),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_734),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_659),
.B(n_536),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_771),
.B(n_800),
.C(n_796),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_879),
.B(n_733),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_777),
.A2(n_677),
.B1(n_754),
.B2(n_752),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_763),
.A2(n_733),
.B(n_612),
.C(n_744),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_763),
.B(n_756),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_772),
.B(n_784),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_762),
.Y(n_952)
);

OAI22x1_ASAP7_75t_L g953 ( 
.A1(n_778),
.A2(n_743),
.B1(n_604),
.B2(n_606),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_796),
.B(n_753),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_896),
.A2(n_710),
.B(n_754),
.C(n_654),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_869),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_766),
.A2(n_718),
.B(n_655),
.C(n_654),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_906),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_856),
.A2(n_934),
.B1(n_895),
.B2(n_902),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_826),
.A2(n_744),
.B(n_742),
.C(n_740),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_891),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_899),
.A2(n_646),
.B(n_665),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_906),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_918),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_856),
.A2(n_697),
.B1(n_692),
.B2(n_682),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_762),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_773),
.B(n_742),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_918),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_778),
.A2(n_663),
.B1(n_667),
.B2(n_655),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_SL g970 ( 
.A1(n_940),
.A2(n_646),
.B(n_718),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_800),
.B(n_740),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_826),
.A2(n_719),
.B(n_701),
.C(n_699),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_840),
.B(n_641),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_817),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_825),
.B(n_641),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_787),
.B(n_695),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_818),
.B(n_719),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_804),
.Y(n_978)
);

CKINVDCx10_ASAP7_75t_R g979 ( 
.A(n_864),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_877),
.A2(n_691),
.B(n_690),
.C(n_22),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_900),
.B(n_453),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_865),
.B(n_536),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_870),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_859),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_865),
.B(n_915),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_878),
.A2(n_863),
.B(n_886),
.Y(n_986)
);

INVx3_ASAP7_75t_SL g987 ( 
.A(n_820),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_764),
.A2(n_527),
.B(n_478),
.Y(n_988)
);

INVx6_ASAP7_75t_L g989 ( 
.A(n_890),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_880),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_785),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_913),
.A2(n_527),
.B(n_478),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_936),
.A2(n_478),
.B(n_470),
.C(n_514),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_825),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_822),
.B(n_782),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_935),
.B(n_478),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_849),
.A2(n_470),
.B(n_514),
.C(n_484),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_942),
.B(n_470),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_835),
.A2(n_17),
.B(n_19),
.C(n_22),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_775),
.A2(n_470),
.B1(n_514),
.B2(n_484),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_884),
.B(n_514),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_782),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_920),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_921),
.B(n_514),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_795),
.A2(n_484),
.B(n_66),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_849),
.A2(n_484),
.B(n_26),
.C(n_27),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_894),
.A2(n_72),
.B(n_146),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_874),
.A2(n_65),
.B(n_140),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_24),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_921),
.B(n_897),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_898),
.A2(n_153),
.B(n_137),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_890),
.B(n_129),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_835),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_809),
.B(n_31),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_765),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_SL g1016 ( 
.A1(n_907),
.A2(n_32),
.B(n_33),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_875),
.A2(n_83),
.B(n_124),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_809),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_928),
.B(n_77),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_866),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_891),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_920),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_793),
.B(n_125),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_SL g1024 ( 
.A(n_927),
.B(n_35),
.C(n_36),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_850),
.B(n_108),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_801),
.A2(n_107),
.B(n_106),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_850),
.B(n_103),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_916),
.A2(n_98),
.B(n_94),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_799),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_853),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_891),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_922),
.B(n_848),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_801),
.A2(n_93),
.B(n_92),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_L g1034 ( 
.A1(n_766),
.A2(n_38),
.B(n_44),
.C(n_45),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_925),
.A2(n_45),
.B(n_46),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_791),
.A2(n_46),
.B(n_48),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_854),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_775),
.B(n_49),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_891),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_859),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_922),
.B(n_49),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_859),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_905),
.B(n_50),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_888),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_859),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_933),
.B(n_54),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_855),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_860),
.B(n_933),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_798),
.B(n_813),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_864),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_915),
.B(n_798),
.Y(n_1052)
);

AO21x2_ASAP7_75t_L g1053 ( 
.A1(n_795),
.A2(n_908),
.B(n_923),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_837),
.A2(n_843),
.B(n_858),
.C(n_857),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_923),
.A2(n_934),
.B(n_914),
.C(n_944),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_802),
.A2(n_806),
.B(n_847),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_864),
.B(n_905),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_802),
.A2(n_806),
.B(n_847),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_767),
.B(n_769),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_790),
.B(n_792),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_868),
.B(n_903),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_888),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_861),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_SL g1064 ( 
.A(n_938),
.B(n_852),
.C(n_901),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_929),
.B(n_932),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_861),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_797),
.B(n_805),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_813),
.A2(n_882),
.B1(n_889),
.B2(n_885),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_872),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_872),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_872),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_862),
.A2(n_887),
.B(n_930),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_892),
.Y(n_1073)
);

AND3x2_ASAP7_75t_L g1074 ( 
.A(n_901),
.B(n_783),
.C(n_882),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_768),
.A2(n_789),
.B(n_815),
.C(n_816),
.Y(n_1075)
);

AOI221x1_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_910),
.B1(n_943),
.B2(n_831),
.C(n_819),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_811),
.B(n_829),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_787),
.B(n_890),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_909),
.B(n_890),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_871),
.A2(n_931),
.B1(n_842),
.B2(n_788),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_812),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_824),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_919),
.B(n_924),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_909),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_SL g1085 ( 
.A1(n_1038),
.A2(n_945),
.B(n_941),
.C(n_939),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_952),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1055),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_956),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_990),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1010),
.B(n_950),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_959),
.B(n_808),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1052),
.B(n_985),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1030),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1065),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1073),
.B(n_938),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1080),
.A2(n_959),
.B1(n_947),
.B2(n_1010),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_974),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1037),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1015),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_965),
.A2(n_851),
.B(n_828),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_970),
.A2(n_912),
.B(n_873),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1057),
.B(n_770),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_SL g1103 ( 
.A1(n_1080),
.A2(n_861),
.B(n_844),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_977),
.B(n_830),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1036),
.A2(n_810),
.B1(n_814),
.B2(n_821),
.C(n_780),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_971),
.A2(n_1025),
.B1(n_1027),
.B2(n_954),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_1028),
.A2(n_1053),
.B(n_1027),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_960),
.A2(n_867),
.B(n_931),
.C(n_839),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_965),
.A2(n_1025),
.B(n_955),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_967),
.B(n_845),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_953),
.A2(n_833),
.A3(n_827),
.B(n_779),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1072),
.A2(n_876),
.B(n_873),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1032),
.B(n_774),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_994),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1081),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1082),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_946),
.A2(n_871),
.B1(n_842),
.B2(n_788),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1076),
.A2(n_838),
.A3(n_781),
.B(n_807),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1053),
.A2(n_851),
.B(n_799),
.Y(n_1119)
);

AO22x2_ASAP7_75t_L g1120 ( 
.A1(n_1064),
.A2(n_783),
.B1(n_885),
.B2(n_836),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_995),
.B(n_828),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_988),
.A2(n_828),
.B(n_786),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1005),
.A2(n_832),
.B(n_911),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_1028),
.A2(n_794),
.B(n_841),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_SL g1125 ( 
.A1(n_1023),
.A2(n_823),
.B(n_846),
.C(n_803),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_975),
.B(n_823),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1049),
.B(n_917),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1059),
.B(n_893),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1002),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_962),
.A2(n_828),
.B(n_844),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_973),
.B(n_846),
.Y(n_1131)
);

BUFx8_ASAP7_75t_L g1132 ( 
.A(n_1062),
.Y(n_1132)
);

AO21x1_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_883),
.B(n_803),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1014),
.B(n_861),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_981),
.A2(n_937),
.B(n_803),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1043),
.B(n_926),
.C(n_803),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1059),
.B(n_776),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1084),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_997),
.A2(n_803),
.A3(n_776),
.B(n_937),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_993),
.A2(n_776),
.A3(n_937),
.B(n_1006),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1083),
.A2(n_776),
.B1(n_969),
.B2(n_951),
.Y(n_1141)
);

NAND3x1_ASAP7_75t_L g1142 ( 
.A(n_1044),
.B(n_1009),
.C(n_1047),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_978),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1019),
.A2(n_998),
.A3(n_996),
.B(n_1047),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_991),
.B(n_1061),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1060),
.Y(n_1146)
);

AND2x2_ASAP7_75t_SL g1147 ( 
.A(n_948),
.B(n_976),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1074),
.A2(n_1041),
.B1(n_1051),
.B2(n_1068),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_957),
.A2(n_1054),
.B(n_972),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_966),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_1019),
.A2(n_1008),
.B(n_1077),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1018),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1020),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1060),
.B(n_1077),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1067),
.Y(n_1155)
);

AND2x6_ASAP7_75t_L g1156 ( 
.A(n_961),
.B(n_1021),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_998),
.B(n_1048),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1041),
.B(n_958),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_983),
.B(n_1050),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_1035),
.A2(n_1011),
.B1(n_1017),
.B2(n_1033),
.C(n_1026),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1029),
.B(n_989),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1069),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_999),
.A2(n_1013),
.B(n_980),
.C(n_1034),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1070),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1024),
.B(n_1071),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_963),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_985),
.B(n_1052),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_964),
.B(n_1022),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1079),
.B(n_961),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_989),
.B(n_1079),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1007),
.A2(n_1001),
.B(n_1000),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_987),
.B(n_968),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_982),
.A2(n_1004),
.B(n_1012),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1003),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1016),
.A2(n_1004),
.B1(n_1046),
.B2(n_1042),
.C(n_1066),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1063),
.A2(n_984),
.B(n_1040),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_984),
.B(n_1040),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_979),
.B(n_1045),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1063),
.A2(n_1066),
.B(n_1046),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1063),
.A2(n_989),
.B(n_1066),
.Y(n_1181)
);

AOI221x1_ASAP7_75t_L g1182 ( 
.A1(n_1042),
.A2(n_1046),
.B1(n_1021),
.B2(n_1031),
.C(n_1039),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_961),
.B(n_1021),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1031),
.B(n_1039),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1031),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1039),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1078),
.B(n_599),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_SL g1188 ( 
.A(n_1063),
.B(n_1080),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_956),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_959),
.B(n_879),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1010),
.B(n_879),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1055),
.A2(n_959),
.B(n_970),
.Y(n_1192)
);

AO21x2_ASAP7_75t_L g1193 ( 
.A1(n_1055),
.A2(n_1028),
.B(n_795),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_961),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1055),
.A2(n_959),
.A3(n_953),
.B(n_1076),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_992),
.A2(n_1058),
.B(n_1056),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_950),
.B(n_599),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_971),
.A2(n_960),
.B(n_950),
.C(n_670),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_992),
.A2(n_1058),
.B(n_1056),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_989),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_952),
.Y(n_1201)
);

AOI221x1_ASAP7_75t_L g1202 ( 
.A1(n_959),
.A2(n_953),
.B1(n_1055),
.B2(n_1036),
.C(n_775),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1055),
.A2(n_959),
.B(n_970),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_986),
.A2(n_879),
.B(n_863),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_R g1205 ( 
.A(n_974),
.B(n_483),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_989),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_959),
.B(n_879),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_986),
.A2(n_879),
.B(n_863),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1063),
.B(n_1029),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_959),
.A3(n_953),
.B(n_1076),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_956),
.Y(n_1211)
);

NOR2x1_ASAP7_75t_SL g1212 ( 
.A(n_1063),
.B(n_1080),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_946),
.B1(n_1038),
.B2(n_971),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_SL g1214 ( 
.A(n_1063),
.B(n_1080),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_989),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_950),
.A2(n_570),
.B1(n_329),
.B2(n_343),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_971),
.A2(n_960),
.B(n_950),
.C(n_670),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_992),
.A2(n_1058),
.B(n_1056),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1029),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_950),
.B(n_321),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1010),
.B(n_879),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_992),
.A2(n_1058),
.B(n_1056),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_971),
.A2(n_960),
.B(n_950),
.C(n_670),
.Y(n_1223)
);

BUFx8_ASAP7_75t_L g1224 ( 
.A(n_1062),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_992),
.A2(n_1058),
.B(n_1056),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1109),
.A2(n_1208),
.B(n_1204),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1088),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1189),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1086),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1222),
.A2(n_1225),
.B(n_1123),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1096),
.B(n_1090),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1149),
.A2(n_1087),
.B(n_1100),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1118),
.Y(n_1233)
);

INVx4_ASAP7_75t_SL g1234 ( 
.A(n_1111),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1209),
.Y(n_1235)
);

CKINVDCx9p33_ASAP7_75t_R g1236 ( 
.A(n_1178),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1119),
.A2(n_1112),
.B(n_1122),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1089),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1135),
.A2(n_1101),
.B(n_1130),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1211),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1099),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1101),
.A2(n_1173),
.B(n_1203),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1192),
.A2(n_1203),
.B(n_1125),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1200),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1118),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1118),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1170),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1143),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1198),
.B(n_1223),
.C(n_1217),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1191),
.B(n_1221),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1097),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1138),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1106),
.A2(n_1197),
.B1(n_1190),
.B2(n_1207),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1209),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1111),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1106),
.A2(n_1142),
.B(n_1163),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1146),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_L g1262 ( 
.A(n_1220),
.B(n_1202),
.C(n_1216),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1157),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1093),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1098),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1192),
.A2(n_1133),
.B(n_1085),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1213),
.A2(n_1147),
.B1(n_1095),
.B2(n_1205),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1175),
.A2(n_1160),
.B(n_1108),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1157),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1188),
.A2(n_1212),
.B(n_1214),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1134),
.B(n_1092),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1091),
.A2(n_1096),
.B(n_1207),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1201),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1190),
.A2(n_1091),
.B(n_1103),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1094),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1155),
.B(n_1110),
.Y(n_1276)
);

CKINVDCx6p67_ASAP7_75t_R g1277 ( 
.A(n_1200),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1175),
.A2(n_1137),
.B(n_1158),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1153),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1137),
.A2(n_1124),
.B(n_1171),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1107),
.A2(n_1193),
.B(n_1151),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1200),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1139),
.Y(n_1283)
);

AO32x2_ASAP7_75t_L g1284 ( 
.A1(n_1117),
.A2(n_1210),
.A3(n_1195),
.B1(n_1107),
.B2(n_1144),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1105),
.A2(n_1126),
.B(n_1141),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_SL g1286 ( 
.A1(n_1158),
.A2(n_1154),
.B(n_1127),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1195),
.B(n_1210),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1128),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1111),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1171),
.A2(n_1124),
.B(n_1128),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1166),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1193),
.A2(n_1151),
.B(n_1117),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1168),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1154),
.A2(n_1113),
.B(n_1127),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1201),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1215),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1132),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1132),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1148),
.A2(n_1187),
.B1(n_1114),
.B2(n_1104),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1139),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1215),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1113),
.A2(n_1176),
.B(n_1181),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1104),
.B(n_1145),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1182),
.A2(n_1180),
.B(n_1131),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1177),
.A2(n_1121),
.B(n_1168),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1174),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1215),
.B(n_1219),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1136),
.A2(n_1120),
.B1(n_1165),
.B2(n_1164),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1219),
.A2(n_1184),
.B(n_1179),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1092),
.B(n_1170),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1139),
.Y(n_1312)
);

NOR2x1_ASAP7_75t_L g1313 ( 
.A(n_1206),
.B(n_1172),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1120),
.B(n_1210),
.Y(n_1314)
);

OAI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1159),
.A2(n_1162),
.B1(n_1150),
.B2(n_1152),
.C(n_1102),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1184),
.A2(n_1186),
.B(n_1167),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1144),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1224),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1194),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1185),
.B(n_1169),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1186),
.A2(n_1183),
.B(n_1140),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1169),
.B(n_1195),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1194),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1194),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1161),
.B(n_1206),
.C(n_1140),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1140),
.A2(n_1161),
.B(n_1156),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1156),
.A2(n_1198),
.B1(n_1217),
.B2(n_1223),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1156),
.A2(n_1217),
.B(n_1198),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1156),
.A2(n_1220),
.B1(n_424),
.B2(n_666),
.Y(n_1329)
);

CKINVDCx8_ASAP7_75t_R g1330 ( 
.A(n_1097),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1149),
.A2(n_1109),
.B(n_1123),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1198),
.A2(n_1223),
.B(n_1217),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_596),
.B1(n_1038),
.B2(n_1147),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1196),
.A2(n_1218),
.B(n_1199),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1118),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1170),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1209),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1143),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1118),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1088),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1198),
.A2(n_1223),
.B(n_1217),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1086),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1201),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1146),
.B(n_1198),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1213),
.A2(n_596),
.B1(n_1038),
.B2(n_1147),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1088),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1196),
.A2(n_1218),
.B(n_1199),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1200),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1146),
.B(n_1198),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1149),
.A2(n_1109),
.B(n_1087),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1198),
.A2(n_1223),
.B(n_1217),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1118),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1213),
.A2(n_596),
.B1(n_1038),
.B2(n_1147),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1088),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1109),
.A2(n_1133),
.A3(n_1106),
.B(n_1149),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1196),
.A2(n_1218),
.B(n_1199),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1088),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1118),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1149),
.A2(n_1087),
.B(n_1109),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1198),
.A2(n_1217),
.B1(n_1223),
.B2(n_1090),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1088),
.Y(n_1361)
);

CKINVDCx6p67_ASAP7_75t_R g1362 ( 
.A(n_1250),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1276),
.B(n_1254),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1307),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_SL g1365 ( 
.A(n_1325),
.B(n_1327),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1238),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1246),
.A2(n_1360),
.B(n_1296),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1249),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1226),
.A2(n_1274),
.B(n_1332),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1249),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1276),
.B(n_1303),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1266),
.A2(n_1245),
.B(n_1341),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1314),
.B(n_1344),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1271),
.B(n_1267),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1295),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1314),
.B(n_1344),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1262),
.A2(n_1333),
.B1(n_1345),
.B2(n_1353),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1231),
.B(n_1343),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1349),
.B(n_1322),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1309),
.A2(n_1315),
.B1(n_1251),
.B2(n_1329),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1275),
.B(n_1349),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1246),
.A2(n_1296),
.B(n_1351),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1260),
.A2(n_1285),
.B(n_1328),
.C(n_1243),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1231),
.B(n_1278),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1240),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1249),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1299),
.A2(n_1244),
.B1(n_1273),
.B2(n_1313),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1257),
.A2(n_1286),
.B(n_1294),
.C(n_1241),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1359),
.A2(n_1350),
.B(n_1268),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1242),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1250),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1286),
.A2(n_1294),
.B(n_1342),
.C(n_1241),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1278),
.B(n_1287),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1252),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1271),
.B(n_1311),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1261),
.B(n_1293),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1249),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1359),
.A2(n_1350),
.B(n_1268),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1229),
.A2(n_1342),
.B1(n_1227),
.B2(n_1228),
.C(n_1361),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1311),
.B(n_1229),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1244),
.A2(n_1292),
.B(n_1239),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1249),
.B(n_1336),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1236),
.A2(n_1277),
.B(n_1270),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1338),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_L g1405 ( 
.A(n_1277),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1244),
.A2(n_1320),
.B1(n_1261),
.B2(n_1336),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1253),
.A2(n_1270),
.B(n_1340),
.C(n_1357),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1282),
.B(n_1301),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1266),
.A2(n_1245),
.B(n_1243),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1278),
.B(n_1287),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1246),
.A2(n_1301),
.B(n_1348),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1306),
.B(n_1346),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1282),
.A2(n_1348),
.B(n_1308),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1306),
.B(n_1354),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1336),
.A2(n_1319),
.B1(n_1256),
.B2(n_1288),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1330),
.A2(n_1234),
.B(n_1298),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1292),
.A2(n_1239),
.B(n_1281),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1288),
.B(n_1265),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1284),
.B(n_1355),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1326),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1319),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1230),
.A2(n_1290),
.B(n_1237),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1336),
.A2(n_1256),
.B1(n_1330),
.B2(n_1308),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1336),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_SL g1428 ( 
.A1(n_1234),
.A2(n_1298),
.B(n_1304),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1284),
.B(n_1355),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1230),
.A2(n_1290),
.B(n_1237),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1264),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1308),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1272),
.B(n_1355),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1316),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1272),
.B(n_1355),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1310),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1297),
.A2(n_1279),
.B1(n_1318),
.B2(n_1255),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1355),
.B(n_1323),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1324),
.B(n_1305),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1310),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1284),
.B(n_1259),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1305),
.B(n_1316),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_L g1443 ( 
.A(n_1235),
.B(n_1258),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1321),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1318),
.A2(n_1317),
.B(n_1281),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1235),
.B(n_1258),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1304),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1234),
.A2(n_1284),
.B(n_1297),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1235),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1279),
.A2(n_1255),
.B1(n_1258),
.B2(n_1337),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1337),
.A2(n_1312),
.B1(n_1300),
.B2(n_1283),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1337),
.B(n_1259),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1289),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1302),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1233),
.A2(n_1358),
.B(n_1339),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1283),
.B(n_1312),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1300),
.A2(n_1358),
.B(n_1352),
.C(n_1339),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1247),
.B(n_1248),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1280),
.B(n_1232),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1331),
.B(n_1352),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1248),
.B(n_1335),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1334),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1434),
.Y(n_1463)
);

INVxp33_ASAP7_75t_SL g1464 ( 
.A(n_1437),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1453),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1384),
.B(n_1356),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1444),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1369),
.B(n_1422),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1384),
.B(n_1393),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1393),
.B(n_1412),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1419),
.A2(n_1389),
.B(n_1398),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1412),
.B(n_1379),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1433),
.A2(n_1435),
.B(n_1383),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1377),
.A2(n_1380),
.B1(n_1365),
.B2(n_1387),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1378),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1401),
.A2(n_1459),
.B(n_1447),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1458),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1461),
.Y(n_1479)
);

CKINVDCx6p67_ASAP7_75t_R g1480 ( 
.A(n_1362),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1461),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1422),
.B(n_1436),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1440),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1454),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1426),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1442),
.A2(n_1430),
.B(n_1424),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1402),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1421),
.B(n_1429),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1381),
.B(n_1371),
.Y(n_1492)
);

AOI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1424),
.A2(n_1430),
.B(n_1372),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1439),
.B(n_1456),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1363),
.B(n_1366),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1455),
.A2(n_1460),
.B(n_1457),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1421),
.A2(n_1429),
.B(n_1460),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1385),
.B(n_1390),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1411),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1394),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1427),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1372),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1372),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1431),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1445),
.A2(n_1451),
.B(n_1441),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1396),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1388),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1441),
.A2(n_1456),
.B(n_1409),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1375),
.A2(n_1362),
.B1(n_1364),
.B2(n_1391),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1462),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1443),
.A2(n_1382),
.B(n_1367),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1452),
.B(n_1462),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1392),
.A2(n_1420),
.B(n_1443),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1407),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1400),
.B(n_1402),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1399),
.A2(n_1415),
.B(n_1406),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1408),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1470),
.B(n_1402),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_L g1520 ( 
.A(n_1511),
.B(n_1446),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1470),
.B(n_1374),
.Y(n_1521)
);

BUFx2_ASAP7_75t_SL g1522 ( 
.A(n_1511),
.Y(n_1522)
);

INVx3_ASAP7_75t_SL g1523 ( 
.A(n_1480),
.Y(n_1523)
);

NOR4xp25_ASAP7_75t_SL g1524 ( 
.A(n_1507),
.B(n_1423),
.C(n_1449),
.D(n_1428),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1482),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1475),
.A2(n_1464),
.B1(n_1517),
.B2(n_1507),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1470),
.B(n_1368),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1476),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.B(n_1368),
.Y(n_1530)
);

NAND4xp25_ASAP7_75t_L g1531 ( 
.A(n_1475),
.B(n_1404),
.C(n_1450),
.D(n_1425),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1500),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1497),
.B(n_1370),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1517),
.A2(n_1391),
.B1(n_1417),
.B2(n_1405),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1501),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1509),
.A2(n_1426),
.B1(n_1395),
.B2(n_1405),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1502),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1370),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1471),
.B(n_1386),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1504),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1484),
.Y(n_1541)
);

NAND4xp25_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1410),
.C(n_1413),
.D(n_1403),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1386),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1497),
.B(n_1397),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1499),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1471),
.B(n_1397),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1432),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1497),
.B(n_1432),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1426),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1473),
.B(n_1405),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1473),
.B(n_1418),
.Y(n_1552)
);

OR2x6_ASAP7_75t_SL g1553 ( 
.A(n_1550),
.B(n_1512),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1539),
.B(n_1471),
.Y(n_1555)
);

AOI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1526),
.A2(n_1495),
.B1(n_1492),
.B2(n_1506),
.C(n_1515),
.Y(n_1556)
);

OAI31xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1531),
.A2(n_1483),
.A3(n_1486),
.B(n_1473),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1549),
.B(n_1490),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1526),
.A2(n_1480),
.B1(n_1510),
.B2(n_1512),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1549),
.B(n_1490),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_L g1561 ( 
.A1(n_1531),
.A2(n_1510),
.B(n_1495),
.C(n_1468),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1549),
.B(n_1490),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1505),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1534),
.B(n_1468),
.C(n_1515),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1547),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1522),
.A2(n_1505),
.B1(n_1496),
.B2(n_1514),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1519),
.B(n_1505),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1534),
.A2(n_1506),
.B1(n_1498),
.B2(n_1465),
.C(n_1494),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1536),
.B(n_1465),
.C(n_1477),
.Y(n_1571)
);

AOI222xp33_ASAP7_75t_L g1572 ( 
.A1(n_1528),
.A2(n_1486),
.B1(n_1483),
.B2(n_1494),
.C1(n_1513),
.C2(n_1498),
.Y(n_1572)
);

OAI33xp33_ASAP7_75t_L g1573 ( 
.A1(n_1547),
.A2(n_1550),
.A3(n_1543),
.B1(n_1540),
.B2(n_1532),
.B3(n_1535),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1539),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1522),
.A2(n_1494),
.B1(n_1483),
.B2(n_1486),
.C(n_1466),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1463),
.C(n_1466),
.D(n_1485),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_R g1579 ( 
.A(n_1523),
.B(n_1487),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1546),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1545),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1508),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1523),
.A2(n_1512),
.B1(n_1489),
.B2(n_1487),
.Y(n_1583)
);

NOR4xp25_ASAP7_75t_SL g1584 ( 
.A(n_1524),
.B(n_1463),
.C(n_1485),
.D(n_1467),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1523),
.A2(n_1489),
.B1(n_1487),
.B2(n_1494),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1520),
.B(n_1469),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1552),
.A2(n_1489),
.B1(n_1494),
.B2(n_1505),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1523),
.A2(n_1469),
.B1(n_1487),
.B2(n_1474),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1521),
.B(n_1513),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1545),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1552),
.A2(n_1505),
.B1(n_1514),
.B2(n_1516),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1545),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1541),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1527),
.B(n_1508),
.Y(n_1594)
);

AOI222xp33_ASAP7_75t_L g1595 ( 
.A1(n_1552),
.A2(n_1513),
.B1(n_1481),
.B2(n_1479),
.C1(n_1478),
.C2(n_1466),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1521),
.B(n_1518),
.Y(n_1596)
);

AOI33xp33_ASAP7_75t_L g1597 ( 
.A1(n_1524),
.A2(n_1503),
.A3(n_1518),
.B1(n_1481),
.B2(n_1479),
.B3(n_1478),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1581),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1566),
.B(n_1548),
.Y(n_1599)
);

AO21x2_ASAP7_75t_L g1600 ( 
.A1(n_1571),
.A2(n_1493),
.B(n_1472),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1591),
.A2(n_1493),
.B(n_1488),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1581),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1593),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1593),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_SL g1605 ( 
.A(n_1584),
.B(n_1469),
.C(n_1551),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1563),
.B(n_1568),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1570),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1555),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1590),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1555),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1563),
.B(n_1530),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1592),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1592),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1567),
.B(n_1542),
.C(n_1520),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1582),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1575),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_L g1619 ( 
.A(n_1565),
.B(n_1542),
.C(n_1502),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1578),
.Y(n_1621)
);

BUFx8_ASAP7_75t_L g1622 ( 
.A(n_1561),
.Y(n_1622)
);

NOR2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1577),
.B(n_1529),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1587),
.A2(n_1488),
.B(n_1499),
.Y(n_1624)
);

AO21x1_ASAP7_75t_L g1625 ( 
.A1(n_1559),
.A2(n_1537),
.B(n_1548),
.Y(n_1625)
);

INVx4_ASAP7_75t_SL g1626 ( 
.A(n_1586),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1568),
.B(n_1530),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1570),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1596),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1553),
.Y(n_1632)
);

BUFx8_ASAP7_75t_L g1633 ( 
.A(n_1554),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1594),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

AND2x6_ASAP7_75t_SL g1636 ( 
.A(n_1564),
.B(n_1551),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1632),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1632),
.B(n_1553),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1631),
.B(n_1557),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1604),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1609),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1616),
.A2(n_1569),
.B(n_1556),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1623),
.Y(n_1643)
);

NAND4xp75_ASAP7_75t_L g1644 ( 
.A(n_1625),
.B(n_1624),
.C(n_1616),
.D(n_1619),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1606),
.B(n_1558),
.Y(n_1645)
);

OR2x6_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1586),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1527),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1611),
.B(n_1521),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1631),
.B(n_1572),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1623),
.B(n_1529),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1604),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1606),
.B(n_1558),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1604),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1630),
.B(n_1595),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1529),
.Y(n_1655)
);

AO221x1_ASAP7_75t_L g1656 ( 
.A1(n_1621),
.A2(n_1588),
.B1(n_1583),
.B2(n_1585),
.C(n_1525),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1603),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1611),
.B(n_1560),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1576),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1603),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1606),
.B(n_1626),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1626),
.B(n_1560),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1626),
.B(n_1562),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1605),
.B(n_1586),
.Y(n_1664)
);

OAI31xp33_ASAP7_75t_L g1665 ( 
.A1(n_1609),
.A2(n_1588),
.A3(n_1551),
.B(n_1548),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1626),
.B(n_1562),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1622),
.B(n_1579),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1608),
.B(n_1508),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1618),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1508),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1636),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1629),
.B(n_1508),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1554),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1618),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1636),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1633),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1629),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1598),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1626),
.B(n_1554),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1650),
.B(n_1626),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1675),
.A2(n_1605),
.B1(n_1586),
.B2(n_1599),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1641),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1640),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1637),
.B(n_1625),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1651),
.Y(n_1685)
);

AOI32xp33_ASAP7_75t_L g1686 ( 
.A1(n_1671),
.A2(n_1622),
.A3(n_1625),
.B1(n_1599),
.B2(n_1627),
.Y(n_1686)
);

NAND2xp67_ASAP7_75t_SL g1687 ( 
.A(n_1638),
.B(n_1661),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1664),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1638),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1642),
.B(n_1635),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1650),
.B(n_1612),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1650),
.A2(n_1628),
.B(n_1602),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1661),
.B(n_1612),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1644),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1644),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1676),
.B(n_1612),
.Y(n_1696)
);

NAND2x1_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1653),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1667),
.B(n_1607),
.Y(n_1699)
);

AOI322xp5_ASAP7_75t_L g1700 ( 
.A1(n_1675),
.A2(n_1627),
.A3(n_1635),
.B1(n_1530),
.B2(n_1538),
.C1(n_1544),
.C2(n_1533),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1678),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1657),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1634),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1627),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1674),
.B(n_1634),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1677),
.B(n_1634),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1668),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1668),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1648),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1670),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1713)
);

AOI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1665),
.A2(n_1601),
.B(n_1573),
.C(n_1622),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1713),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1654),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

CKINVDCx16_ASAP7_75t_R g1719 ( 
.A(n_1713),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1699),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1699),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1649),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1690),
.B(n_1659),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1688),
.B(n_1662),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.B(n_1684),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1699),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_L g1727 ( 
.A(n_1694),
.B(n_1646),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1685),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1711),
.B(n_1658),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1658),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1696),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1694),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1695),
.B(n_1655),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1695),
.A2(n_1646),
.B1(n_1656),
.B2(n_1622),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1680),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1727),
.B(n_1695),
.C(n_1686),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1719),
.B(n_1707),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1716),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1736),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1718),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1738),
.A2(n_1697),
.B1(n_1714),
.B2(n_1646),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1725),
.A2(n_1697),
.B(n_1714),
.C(n_1705),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1736),
.B(n_1739),
.Y(n_1749)
);

OAI321xp33_ASAP7_75t_L g1750 ( 
.A1(n_1717),
.A2(n_1686),
.A3(n_1680),
.B1(n_1687),
.B2(n_1705),
.C(n_1691),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1704),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1737),
.A2(n_1700),
.B(n_1687),
.C(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1724),
.B(n_1704),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1730),
.B(n_1693),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1717),
.A2(n_1700),
.B(n_1692),
.C(n_1597),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1722),
.A2(n_1673),
.B(n_1679),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1730),
.B(n_1673),
.Y(n_1757)
);

OAI332xp33_ASAP7_75t_L g1758 ( 
.A1(n_1720),
.A2(n_1706),
.A3(n_1702),
.B1(n_1698),
.B2(n_1708),
.B3(n_1703),
.C1(n_1672),
.C2(n_1701),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1751),
.B(n_1734),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1741),
.B(n_1735),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1744),
.B(n_1734),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1744),
.B(n_1721),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1744),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1753),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1749),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1754),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1741),
.B(n_1726),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1740),
.B(n_1731),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1758),
.B(n_1728),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1742),
.B(n_1731),
.Y(n_1770)
);

AOI222xp33_ASAP7_75t_L g1771 ( 
.A1(n_1768),
.A2(n_1750),
.B1(n_1745),
.B2(n_1752),
.C1(n_1755),
.C2(n_1743),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1769),
.A2(n_1747),
.B1(n_1745),
.B2(n_1757),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1769),
.A2(n_1748),
.B1(n_1755),
.B2(n_1746),
.C(n_1756),
.Y(n_1773)
);

AOI211x1_ASAP7_75t_SL g1774 ( 
.A1(n_1762),
.A2(n_1708),
.B(n_1701),
.C(n_1712),
.Y(n_1774)
);

OAI22xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1763),
.A2(n_1732),
.B1(n_1733),
.B2(n_1729),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1760),
.A2(n_1767),
.B(n_1761),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1765),
.A2(n_1732),
.B1(n_1702),
.B2(n_1706),
.C(n_1703),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1770),
.A2(n_1692),
.B(n_1701),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1759),
.B(n_1679),
.Y(n_1779)
);

OAI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1771),
.A2(n_1764),
.B(n_1766),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1773),
.A2(n_1712),
.B(n_1710),
.C(n_1709),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1775),
.Y(n_1782)
);

OAI322xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1777),
.A2(n_1712),
.A3(n_1710),
.B1(n_1709),
.B2(n_1634),
.C1(n_1620),
.C2(n_1617),
.Y(n_1783)
);

OAI32xp33_ASAP7_75t_L g1784 ( 
.A1(n_1774),
.A2(n_1672),
.A3(n_1670),
.B1(n_1710),
.B2(n_1709),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1776),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1782),
.Y(n_1786)
);

INVx8_ASAP7_75t_L g1787 ( 
.A(n_1781),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1784),
.B(n_1779),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1783),
.B(n_1772),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1780),
.B(n_1778),
.C(n_1666),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1788),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1789),
.A2(n_1666),
.B1(n_1663),
.B2(n_1662),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1785),
.A2(n_1663),
.B1(n_1633),
.B2(n_1600),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1790),
.A2(n_1617),
.B1(n_1620),
.B2(n_1607),
.C(n_1628),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1786),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1795),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1791),
.B(n_1787),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1792),
.B(n_1787),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1796),
.B(n_1794),
.C(n_1793),
.Y(n_1799)
);

AOI322xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1798),
.A3(n_1797),
.B1(n_1607),
.B2(n_1628),
.C1(n_1652),
.C2(n_1645),
.Y(n_1800)
);

OR3x2_ASAP7_75t_L g1801 ( 
.A(n_1800),
.B(n_1647),
.C(n_1597),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1801),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1628),
.B1(n_1647),
.B2(n_1617),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1803),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1804),
.A2(n_1617),
.B1(n_1620),
.B2(n_1610),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_SL g1807 ( 
.A(n_1805),
.B(n_1645),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1620),
.B1(n_1652),
.B2(n_1633),
.Y(n_1808)
);

AOI22x1_ASAP7_75t_L g1809 ( 
.A1(n_1806),
.A2(n_1610),
.B1(n_1615),
.B2(n_1614),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1808),
.A2(n_1809),
.B(n_1598),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1633),
.B1(n_1614),
.B2(n_1613),
.Y(n_1811)
);

AOI211xp5_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1598),
.B(n_1615),
.C(n_1613),
.Y(n_1812)
);


endmodule