module fake_jpeg_319_n_246 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_246);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_1),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_17),
.B1(n_26),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_30),
.B1(n_29),
.B2(n_14),
.Y(n_103)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_22),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_26),
.B1(n_18),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_67),
.B1(n_79),
.B2(n_14),
.Y(n_117)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_22),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_69),
.Y(n_94)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_23),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_88),
.Y(n_93)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_40),
.B(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_91),
.Y(n_100)
);

XNOR2x1_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_25),
.B1(n_16),
.B2(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_95),
.A2(n_53),
.B1(n_78),
.B2(n_66),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_52),
.A2(n_29),
.B1(n_14),
.B2(n_5),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_109),
.B(n_50),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_29),
.B1(n_14),
.B2(n_5),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_4),
.C(n_5),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_55),
.B1(n_60),
.B2(n_53),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_3),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_126),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_69),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_134),
.Y(n_161)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_139),
.B1(n_142),
.B2(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_90),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_84),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_98),
.C(n_118),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_101),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_51),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_146),
.B(n_107),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_90),
.B1(n_66),
.B2(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_74),
.B1(n_83),
.B2(n_49),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_83),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_64),
.B1(n_51),
.B2(n_68),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_93),
.A2(n_68),
.B(n_89),
.C(n_64),
.D(n_14),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_115),
.B1(n_97),
.B2(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

CKINVDCx10_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_172),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_140),
.B1(n_126),
.B2(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_95),
.B1(n_94),
.B2(n_118),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_163),
.B(n_170),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_104),
.B(n_106),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_106),
.B1(n_89),
.B2(n_94),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_120),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_120),
.B(n_8),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_4),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_134),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_188),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_188),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_152),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_193),
.C(n_201),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_155),
.C(n_149),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_158),
.B1(n_149),
.B2(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_159),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_204),
.C(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_158),
.B1(n_163),
.B2(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_170),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_136),
.B(n_124),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_176),
.B1(n_183),
.B2(n_185),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_178),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_156),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.C(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_192),
.C(n_200),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_196),
.C(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_223),
.C(n_175),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_201),
.C(n_205),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_206),
.B(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_166),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_210),
.A3(n_216),
.B1(n_199),
.B2(n_212),
.C1(n_195),
.C2(n_186),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NAND4xp25_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_190),
.C(n_169),
.D(n_212),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_166),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_145),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_232),
.C(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_229),
.B1(n_231),
.B2(n_136),
.Y(n_240)
);

NOR4xp25_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.C(n_235),
.D(n_190),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_238),
.A3(n_240),
.B1(n_241),
.B2(n_169),
.C1(n_239),
.C2(n_150),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_243),
.C(n_125),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_128),
.Y(n_246)
);


endmodule