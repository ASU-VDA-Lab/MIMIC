module fake_netlist_1_9967_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_SL g3 ( .A(n_1), .Y(n_3) );
BUFx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
OR3x4_ASAP7_75t_SL g5 ( .A(n_3), .B(n_0), .C(n_1), .Y(n_5) );
AOI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_2), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_4), .B1(n_5), .B2(n_0), .C(n_6), .Y(n_8) );
NOR2x1_ASAP7_75t_L g9 ( .A(n_8), .B(n_4), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_4), .B(n_2), .Y(n_11) );
endmodule