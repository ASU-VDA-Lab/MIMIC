module fake_netlist_5_552_n_21 (n_8, n_4, n_5, n_7, n_0, n_2, n_3, n_6, n_1, n_21);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_2;
input n_3;
input n_6;
input n_1;

output n_21;

wire n_16;
wire n_12;
wire n_9;
wire n_18;
wire n_10;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_14;
wire n_13;
wire n_20;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_7),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVxp67_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

OA21x2_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_0),
.B(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

O2A1O1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_10),
.B(n_12),
.C(n_11),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_15),
.A2(n_9),
.B(n_13),
.Y(n_17)
);

AOI221xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.B1(n_13),
.B2(n_4),
.C(n_5),
.Y(n_18)
);

AOI221xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_13),
.B1(n_3),
.B2(n_2),
.C(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

AOI222xp33_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_19),
.B1(n_13),
.B2(n_3),
.C1(n_8),
.C2(n_6),
.Y(n_21)
);


endmodule