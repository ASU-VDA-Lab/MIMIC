module fake_ibex_1874_n_2086 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2086);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2086;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_2083;
wire n_886;
wire n_1010;
wire n_883;
wire n_2044;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2013;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_519;
wire n_1843;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_313),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_164),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_73),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_209),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_335),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_88),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_205),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_299),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_0),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_4),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_173),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_373),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_224),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_277),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_194),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_360),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_62),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_349),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_420),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_38),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_263),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_239),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_289),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_82),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_264),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_244),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_366),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_42),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_377),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_203),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_290),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_136),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_293),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_213),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_186),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_417),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_384),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_398),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_159),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_16),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_94),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_334),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_188),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_28),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_66),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_91),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_369),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_356),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_387),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_124),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_106),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_97),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_350),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_190),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_159),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_167),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_274),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_148),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_352),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_111),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_316),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_305),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_307),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_60),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_132),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_256),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_241),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_107),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_37),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_192),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_28),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_140),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_61),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_406),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_354),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_372),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_23),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_273),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_340),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_298),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_59),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_278),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_312),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_261),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_104),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_79),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_66),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_302),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_332),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_351),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_123),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_64),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_410),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_180),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_144),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_20),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_403),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_99),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_275),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_133),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_284),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_371),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_91),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_50),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_136),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_228),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_42),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_201),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_121),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_131),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_149),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_191),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_1),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_135),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_246),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_220),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_132),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_359),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_160),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_232),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_124),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_282),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_393),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_144),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_143),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_243),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_229),
.Y(n_555)
);

CKINVDCx14_ASAP7_75t_R g556 ( 
.A(n_114),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_269),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_242),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_58),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_399),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_170),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_379),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_140),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_311),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_245),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_46),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_266),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_128),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_310),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_186),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_56),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_262),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_94),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_126),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_213),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_392),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_327),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_401),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_361),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_116),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_333),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_242),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_24),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_171),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_315),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_227),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_344),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_267),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_257),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_285),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_173),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_105),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_342),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_78),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_79),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_157),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_370),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_106),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_31),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g600 ( 
.A(n_59),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_247),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_155),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_89),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_396),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_268),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_139),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_122),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_252),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_168),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_62),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_76),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_194),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_29),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_134),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_324),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_80),
.Y(n_616)
);

CKINVDCx14_ASAP7_75t_R g617 ( 
.A(n_378),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_64),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_97),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_227),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_167),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_13),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_328),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_225),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_44),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_281),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_109),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_96),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_418),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_130),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_113),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_321),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_336),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_4),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_26),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_130),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_6),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_113),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_131),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_255),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_204),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_250),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_34),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_191),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_102),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_31),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_5),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_346),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_51),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_129),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_142),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_60),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_168),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_141),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_17),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_177),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_296),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_155),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_260),
.Y(n_659)
);

CKINVDCx16_ASAP7_75t_R g660 ( 
.A(n_304),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_288),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_314),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_223),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_80),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_135),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_137),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_414),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_190),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_347),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_53),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_246),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_139),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_107),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_172),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_196),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_280),
.Y(n_676)
);

BUFx10_ASAP7_75t_L g677 ( 
.A(n_287),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_270),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_48),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_74),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_165),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_276),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_32),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_197),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_251),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_329),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_326),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_196),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_114),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_300),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_162),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_178),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_47),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_368),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_341),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_226),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_380),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_18),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_34),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_26),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_386),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_415),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_226),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_295),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_253),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_363),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_358),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_301),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_600),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_424),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_424),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_555),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_603),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_595),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_423),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_660),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_686),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_696),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_500),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_490),
.B(n_690),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_490),
.B(n_1),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_515),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_549),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_591),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_445),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_431),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_621),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_591),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_445),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_679),
.B(n_2),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_644),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_644),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_698),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_681),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_431),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_690),
.B(n_3),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_468),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_446),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_446),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_468),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_564),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_564),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_491),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_574),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_454),
.B(n_3),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_523),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_528),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_496),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_556),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_528),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_537),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_574),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_537),
.Y(n_757)
);

INVxp33_ASAP7_75t_SL g758 ( 
.A(n_449),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_541),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_542),
.B(n_5),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_652),
.B(n_7),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_572),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_598),
.B(n_7),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_625),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_625),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_686),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_650),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_650),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_433),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_680),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_428),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_572),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_695),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_433),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_444),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_458),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_695),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_439),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_451),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_470),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_471),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_439),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_472),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_574),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_469),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_657),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_432),
.B(n_8),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_669),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_669),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_477),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_482),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_483),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_469),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_493),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_678),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_497),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_481),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_588),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_481),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_596),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_434),
.B(n_436),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_456),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_485),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_485),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_499),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_492),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_520),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_456),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_492),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_522),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_526),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_513),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_678),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_687),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_460),
.B(n_461),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_687),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_760),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_710),
.B(n_715),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_773),
.B(n_447),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_719),
.A2(n_457),
.B(n_453),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_710),
.B(n_450),
.Y(n_821)
);

AND3x2_ASAP7_75t_L g822 ( 
.A(n_731),
.B(n_426),
.C(n_547),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_760),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_719),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_711),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_712),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_773),
.B(n_588),
.Y(n_828)
);

CKINVDCx6p67_ASAP7_75t_R g829 ( 
.A(n_756),
.Y(n_829)
);

XOR2xp5_ASAP7_75t_L g830 ( 
.A(n_709),
.B(n_714),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_766),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_713),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_747),
.B(n_694),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_766),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_798),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_722),
.B(n_464),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_777),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_742),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_717),
.B(n_617),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_779),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_738),
.B(n_596),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_743),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_721),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_723),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_725),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_716),
.B(n_460),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_SL g848 ( 
.A(n_752),
.B(n_694),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_726),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_727),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_802),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_728),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_758),
.A2(n_566),
.B1(n_465),
.B2(n_466),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_732),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_750),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_735),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_753),
.B(n_808),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_718),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_751),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_736),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_754),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_755),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_737),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_757),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_768),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_771),
.B(n_474),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_759),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_709),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_776),
.B(n_422),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_780),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_775),
.B(n_552),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_764),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_765),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_781),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_748),
.B(n_479),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_767),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_801),
.B(n_465),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_770),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_724),
.B(n_740),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_783),
.B(n_480),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_790),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_791),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_784),
.B(n_596),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_800),
.B(n_448),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_792),
.B(n_448),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_794),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_796),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_805),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_807),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

INVx6_ASAP7_75t_L g891 ( 
.A(n_763),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_811),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_787),
.B(n_749),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_761),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_734),
.B(n_466),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_729),
.B(n_467),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_733),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_741),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_744),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_745),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_746),
.B(n_762),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_772),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_786),
.B(n_692),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_788),
.B(n_692),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_789),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_720),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_795),
.B(n_484),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_730),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_813),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_816),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_730),
.A2(n_566),
.B1(n_699),
.B2(n_693),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_739),
.B(n_693),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_739),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_812),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_769),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_769),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_809),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_774),
.B(n_699),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_774),
.Y(n_920)
);

BUFx8_ASAP7_75t_L g921 ( 
.A(n_778),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_778),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_809),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_782),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_782),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_785),
.B(n_448),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_806),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_785),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_793),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_793),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_806),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_797),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_797),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_799),
.B(n_553),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_799),
.B(n_700),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_803),
.B(n_605),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_803),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_804),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_804),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_710),
.B(n_605),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_730),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_722),
.B(n_700),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_760),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_760),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_760),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_815),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_710),
.B(n_605),
.Y(n_947)
);

BUFx8_ASAP7_75t_L g948 ( 
.A(n_715),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_760),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_760),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_718),
.B(n_517),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_760),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_760),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_R g954 ( 
.A(n_758),
.B(n_705),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_779),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_760),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_760),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_760),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_722),
.B(n_706),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_773),
.B(n_486),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_719),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_760),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_760),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_722),
.B(n_708),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_760),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_773),
.B(n_489),
.Y(n_966)
);

INVx6_ASAP7_75t_L g967 ( 
.A(n_760),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_760),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_779),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_760),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_760),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_779),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_710),
.A2(n_427),
.B1(n_430),
.B2(n_425),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_760),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_760),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_758),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_760),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_719),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_773),
.B(n_502),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_719),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_760),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_710),
.B(n_662),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_719),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_719),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_760),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_711),
.B(n_568),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_719),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_760),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_760),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_760),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_946),
.B(n_422),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_967),
.Y(n_992)
);

AO22x2_ASAP7_75t_L g993 ( 
.A1(n_817),
.A2(n_571),
.B1(n_575),
.B2(n_573),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_885),
.B(n_582),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_821),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_818),
.B(n_545),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_940),
.B(n_437),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_947),
.B(n_441),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_826),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_829),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_827),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_982),
.B(n_476),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_832),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_942),
.B(n_452),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_841),
.B(n_478),
.Y(n_1005)
);

INVx8_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_913),
.B(n_583),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_SL g1008 ( 
.A(n_829),
.B(n_455),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_825),
.A2(n_524),
.B1(n_592),
.B2(n_513),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_887),
.B(n_455),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_944),
.B(n_676),
.Y(n_1011)
);

NOR2x1p5_ASAP7_75t_L g1012 ( 
.A(n_976),
.B(n_487),
.Y(n_1012)
);

NOR2x1p5_ASAP7_75t_L g1013 ( 
.A(n_976),
.B(n_910),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_851),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_962),
.Y(n_1015)
);

INVx4_ASAP7_75t_SL g1016 ( 
.A(n_828),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_851),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_840),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_888),
.B(n_459),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_962),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_884),
.B(n_602),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_883),
.B(n_616),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_955),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_869),
.B(n_459),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_986),
.B(n_619),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_963),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_888),
.B(n_462),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_986),
.B(n_624),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_890),
.B(n_462),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_981),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_890),
.B(n_475),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_981),
.A2(n_634),
.B1(n_636),
.B2(n_630),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_981),
.A2(n_641),
.B1(n_642),
.B2(n_638),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_869),
.B(n_697),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_989),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_989),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_870),
.B(n_697),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_865),
.B(n_702),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_989),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_892),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_874),
.B(n_702),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_959),
.B(n_704),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_856),
.Y(n_1046)
);

AND2x2_ASAP7_75t_SL g1047 ( 
.A(n_936),
.B(n_703),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_856),
.Y(n_1048)
);

INVx6_ASAP7_75t_L g1049 ( 
.A(n_892),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_941),
.A2(n_524),
.B1(n_592),
.B2(n_519),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_969),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_892),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_948),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_881),
.B(n_704),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_943),
.A2(n_643),
.B1(n_664),
.B2(n_663),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_871),
.A2(n_671),
.B1(n_672),
.B2(n_666),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_972),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_892),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_823),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_842),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_876),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_954),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_882),
.B(n_708),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_857),
.B(n_494),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_871),
.B(n_673),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_886),
.B(n_510),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_889),
.B(n_516),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_823),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_910),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_936),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_944),
.B(n_676),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_871),
.B(n_858),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_964),
.B(n_707),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_837),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_894),
.B(n_684),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_891),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_971),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_971),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_974),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_974),
.Y(n_1080)
);

AND3x2_ASAP7_75t_L g1081 ( 
.A(n_868),
.B(n_639),
.C(n_519),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_847),
.B(n_495),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_894),
.B(n_685),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_910),
.B(n_688),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_945),
.B(n_985),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_853),
.B(n_498),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_891),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_906),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_867),
.Y(n_1089)
);

OAI221xp5_ASAP7_75t_L g1090 ( 
.A1(n_950),
.A2(n_689),
.B1(n_665),
.B2(n_653),
.C(n_594),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_975),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_973),
.B(n_504),
.Y(n_1092)
);

INVx4_ASAP7_75t_SL g1093 ( 
.A(n_828),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_949),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_949),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_855),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_952),
.A2(n_691),
.B1(n_640),
.B2(n_658),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_855),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_866),
.B(n_508),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_875),
.B(n_677),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_836),
.B(n_957),
.C(n_956),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_838),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_953),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_877),
.B(n_662),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_926),
.B(n_896),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_919),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_899),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_953),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_875),
.B(n_707),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_SL g1110 ( 
.A(n_958),
.B(n_677),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_861),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_935),
.Y(n_1112)
);

INVxp33_ASAP7_75t_L g1113 ( 
.A(n_830),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_921),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_861),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_861),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_879),
.B(n_463),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_953),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_911),
.B(n_895),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_836),
.B(n_473),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_954),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_970),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_861),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_965),
.B(n_968),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_864),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_820),
.A2(n_551),
.B(n_546),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_864),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_912),
.B(n_514),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_921),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_893),
.B(n_488),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_970),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_977),
.B(n_429),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_878),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_878),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_820),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_941),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_839),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_921),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_839),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_988),
.B(n_435),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_843),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_911),
.B(n_531),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_990),
.B(n_438),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_907),
.A2(n_533),
.B1(n_534),
.B2(n_532),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_843),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_828),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_859),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_824),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_907),
.A2(n_536),
.B1(n_538),
.B2(n_535),
.Y(n_1149)
);

CKINVDCx16_ASAP7_75t_R g1150 ( 
.A(n_833),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_898),
.B(n_539),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_903),
.B(n_632),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_831),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_904),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_862),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_900),
.B(n_540),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_897),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_908),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_901),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_844),
.B(n_440),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_845),
.B(n_569),
.Y(n_1161)
);

AND2x6_ASAP7_75t_L g1162 ( 
.A(n_831),
.B(n_834),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_872),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_L g1164 ( 
.A(n_902),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_846),
.B(n_577),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_934),
.B(n_543),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_834),
.B(n_961),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_905),
.B(n_909),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_849),
.B(n_850),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_852),
.B(n_585),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_934),
.B(n_544),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_854),
.B(n_587),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_860),
.B(n_442),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_873),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_863),
.B(n_548),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_880),
.B(n_554),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_880),
.B(n_558),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_1009),
.A2(n_924),
.B1(n_925),
.B2(n_923),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1059),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1068),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1077),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1037),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1014),
.B(n_443),
.Y(n_1183)
);

OAI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1014),
.A2(n_1057),
.B1(n_1017),
.B2(n_1090),
.C(n_996),
.Y(n_1184)
);

AO22x2_ASAP7_75t_L g1185 ( 
.A1(n_1009),
.A2(n_924),
.B1(n_925),
.B2(n_923),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1078),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1079),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1080),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1017),
.A2(n_1057),
.B1(n_1090),
.B2(n_1056),
.C(n_1025),
.Y(n_1189)
);

OR2x6_ASAP7_75t_SL g1190 ( 
.A(n_1000),
.B(n_916),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1091),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_999),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1013),
.B(n_1084),
.Y(n_1193)
);

AO22x2_ASAP7_75t_L g1194 ( 
.A1(n_1070),
.A2(n_931),
.B1(n_933),
.B2(n_927),
.Y(n_1194)
);

AO22x2_ASAP7_75t_L g1195 ( 
.A1(n_1088),
.A2(n_927),
.B1(n_915),
.B2(n_918),
.Y(n_1195)
);

OR2x2_ASAP7_75t_SL g1196 ( 
.A(n_1150),
.B(n_920),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1053),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1003),
.Y(n_1199)
);

AO22x2_ASAP7_75t_L g1200 ( 
.A1(n_1159),
.A2(n_922),
.B1(n_929),
.B2(n_917),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1082),
.B(n_822),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1159),
.A2(n_937),
.B1(n_938),
.B2(n_932),
.Y(n_1202)
);

OAI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_1106),
.A2(n_848),
.B1(n_960),
.B2(n_966),
.C(n_819),
.Y(n_1203)
);

OAI221xp5_ASAP7_75t_L g1204 ( 
.A1(n_1112),
.A2(n_960),
.B1(n_979),
.B2(n_966),
.C(n_819),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1006),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1008),
.A2(n_1110),
.B1(n_1051),
.B2(n_1121),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1105),
.A2(n_951),
.B1(n_979),
.B2(n_561),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1103),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1108),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1006),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1107),
.B(n_1069),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1089),
.Y(n_1212)
);

AO22x2_ASAP7_75t_L g1213 ( 
.A1(n_1097),
.A2(n_914),
.B1(n_916),
.B2(n_928),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1118),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1114),
.Y(n_1215)
);

AO22x2_ASAP7_75t_L g1216 ( 
.A1(n_1097),
.A2(n_930),
.B1(n_668),
.B2(n_670),
.Y(n_1216)
);

AO22x2_ASAP7_75t_L g1217 ( 
.A1(n_1176),
.A2(n_668),
.B1(n_670),
.B2(n_658),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1047),
.B(n_920),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1176),
.A2(n_691),
.B1(n_939),
.B2(n_920),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1122),
.Y(n_1220)
);

NOR2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1129),
.B(n_1138),
.Y(n_1221)
);

OAI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1112),
.A2(n_565),
.B1(n_570),
.B2(n_563),
.C(n_559),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1131),
.Y(n_1223)
);

AO22x2_ASAP7_75t_L g1224 ( 
.A1(n_1177),
.A2(n_939),
.B1(n_604),
.B2(n_615),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1040),
.B(n_978),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1158),
.Y(n_1226)
);

OAI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1128),
.A2(n_1007),
.B1(n_995),
.B2(n_1019),
.C(n_1060),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1050),
.A2(n_939),
.B1(n_626),
.B2(n_629),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1072),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1137),
.Y(n_1230)
);

OAI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1144),
.A2(n_586),
.B1(n_589),
.B2(n_584),
.C(n_580),
.Y(n_1231)
);

NOR2x1p5_ASAP7_75t_L g1232 ( 
.A(n_1005),
.B(n_599),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1155),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1169),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1169),
.Y(n_1235)
);

AO22x2_ASAP7_75t_L g1236 ( 
.A1(n_1121),
.A2(n_633),
.B1(n_648),
.B2(n_597),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1119),
.B(n_978),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_1157),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_992),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_994),
.B(n_980),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_993),
.Y(n_1241)
);

AO22x2_ASAP7_75t_L g1242 ( 
.A1(n_1081),
.A2(n_1142),
.B1(n_1175),
.B2(n_1101),
.Y(n_1242)
);

OAI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1149),
.A2(n_607),
.B1(n_610),
.B2(n_609),
.C(n_601),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_1081),
.A2(n_661),
.B1(n_667),
.B2(n_659),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1136),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_993),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1061),
.B(n_983),
.Y(n_1247)
);

OAI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1154),
.A2(n_613),
.B1(n_618),
.B2(n_612),
.C(n_611),
.Y(n_1248)
);

OAI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1166),
.A2(n_622),
.B1(n_628),
.B2(n_627),
.C(n_620),
.Y(n_1249)
);

OAI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1171),
.A2(n_635),
.B1(n_645),
.B2(n_637),
.C(n_631),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_993),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1055),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1055),
.Y(n_1253)
);

OAI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_1041),
.A2(n_651),
.B1(n_654),
.B2(n_649),
.C(n_646),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1055),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1148),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_997),
.B(n_655),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_998),
.B(n_656),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1142),
.A2(n_701),
.B1(n_987),
.B2(n_984),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_994),
.B(n_987),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1085),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1012),
.Y(n_1262)
);

AO22x2_ASAP7_75t_L g1263 ( 
.A1(n_1175),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1085),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1064),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1124),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1027),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1027),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1044),
.B(n_674),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1054),
.B(n_683),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1113),
.A2(n_1062),
.B1(n_1086),
.B2(n_1092),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1002),
.B(n_675),
.Y(n_1272)
);

AO22x2_ASAP7_75t_L g1273 ( 
.A1(n_1065),
.A2(n_1030),
.B1(n_1083),
.B2(n_1075),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1168),
.B(n_614),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1062),
.B(n_647),
.Y(n_1275)
);

AO22x2_ASAP7_75t_L g1276 ( 
.A1(n_1065),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1063),
.B(n_1099),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1146),
.B(n_647),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1094),
.Y(n_1279)
);

NAND2x1_ASAP7_75t_L g1280 ( 
.A(n_1162),
.B(n_517),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1095),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1141),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1147),
.Y(n_1284)
);

AO22x2_ASAP7_75t_L g1285 ( 
.A1(n_1075),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_1285)
);

AO22x2_ASAP7_75t_L g1286 ( 
.A1(n_1083),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1024),
.A2(n_503),
.B1(n_505),
.B2(n_501),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1024),
.A2(n_507),
.B1(n_509),
.B2(n_506),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1163),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1174),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1063),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1046),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1164),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1048),
.Y(n_1294)
);

OAI221xp5_ASAP7_75t_L g1295 ( 
.A1(n_1120),
.A2(n_518),
.B1(n_521),
.B2(n_512),
.C(n_511),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1023),
.B(n_517),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1066),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1151),
.B(n_517),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1151),
.B(n_19),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1156),
.A2(n_527),
.B1(n_529),
.B2(n_525),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1067),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1010),
.B(n_530),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_SL g1303 ( 
.A(n_1156),
.Y(n_1303)
);

OAI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1034),
.A2(n_1035),
.B1(n_1117),
.B2(n_1104),
.C(n_1164),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1073),
.B(n_21),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1076),
.A2(n_1087),
.B1(n_1029),
.B2(n_1031),
.Y(n_1306)
);

AO22x2_ASAP7_75t_L g1307 ( 
.A1(n_1021),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_991),
.B(n_550),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1021),
.Y(n_1309)
);

AO22x2_ASAP7_75t_L g1310 ( 
.A1(n_1029),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_1310)
);

AO22x2_ASAP7_75t_L g1311 ( 
.A1(n_1033),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_1311)
);

AO22x2_ASAP7_75t_L g1312 ( 
.A1(n_1033),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1167),
.Y(n_1313)
);

AO22x2_ASAP7_75t_L g1314 ( 
.A1(n_1026),
.A2(n_35),
.B1(n_30),
.B2(n_33),
.Y(n_1314)
);

AO22x2_ASAP7_75t_L g1315 ( 
.A1(n_1036),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1315)
);

OAI221xp5_ASAP7_75t_L g1316 ( 
.A1(n_1130),
.A2(n_562),
.B1(n_567),
.B2(n_560),
.C(n_557),
.Y(n_1316)
);

OAI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1152),
.A2(n_578),
.B1(n_581),
.B2(n_579),
.C(n_576),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1153),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_SL g1319 ( 
.A(n_1011),
.Y(n_1319)
);

AO22x2_ASAP7_75t_L g1320 ( 
.A1(n_1028),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1139),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1011),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1004),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1100),
.B(n_39),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1132),
.Y(n_1325)
);

AO22x2_ASAP7_75t_L g1326 ( 
.A1(n_1028),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_1326)
);

AND2x6_ASAP7_75t_L g1327 ( 
.A(n_1135),
.B(n_623),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1039),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1328)
);

AO22x2_ASAP7_75t_L g1329 ( 
.A1(n_1109),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1161),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1161),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1165),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1160),
.Y(n_1333)
);

AO22x2_ASAP7_75t_L g1334 ( 
.A1(n_1016),
.A2(n_1093),
.B1(n_1170),
.B2(n_1165),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1045),
.B(n_593),
.C(n_590),
.Y(n_1335)
);

AO22x2_ASAP7_75t_L g1336 ( 
.A1(n_1016),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1336)
);

AO22x2_ASAP7_75t_L g1337 ( 
.A1(n_1016),
.A2(n_52),
.B1(n_49),
.B2(n_51),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1172),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1140),
.B(n_52),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1172),
.Y(n_1340)
);

AO22x2_ASAP7_75t_L g1341 ( 
.A1(n_1093),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1341)
);

BUFx8_ASAP7_75t_L g1342 ( 
.A(n_1071),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1102),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1093),
.A2(n_57),
.B1(n_54),
.B2(n_55),
.Y(n_1344)
);

AO22x2_ASAP7_75t_L g1345 ( 
.A1(n_1015),
.A2(n_61),
.B1(n_57),
.B2(n_58),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1173),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1143),
.Y(n_1347)
);

AO22x2_ASAP7_75t_L g1348 ( 
.A1(n_1020),
.A2(n_67),
.B1(n_63),
.B2(n_65),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1167),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1022),
.B(n_63),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1126),
.B(n_65),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1123),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1032),
.B(n_67),
.Y(n_1353)
);

AO22x2_ASAP7_75t_L g1354 ( 
.A1(n_1038),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1042),
.Y(n_1355)
);

AO22x2_ASAP7_75t_L g1356 ( 
.A1(n_1126),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1234),
.B(n_1235),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1261),
.B(n_1043),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1226),
.B(n_1205),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_SL g1360 ( 
.A(n_1319),
.B(n_1098),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1352),
.B(n_1115),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1206),
.B(n_1115),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1211),
.B(n_1125),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1350),
.B(n_1018),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1193),
.B(n_1264),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_R g1366 ( 
.A(n_1197),
.B(n_1096),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1266),
.B(n_1096),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1297),
.B(n_1116),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1301),
.B(n_1116),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1330),
.B(n_1111),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1331),
.B(n_1332),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1338),
.B(n_1127),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1340),
.B(n_1133),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1309),
.B(n_1299),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1299),
.B(n_1134),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1210),
.B(n_1058),
.Y(n_1376)
);

NAND2xp33_ASAP7_75t_SL g1377 ( 
.A(n_1353),
.B(n_1074),
.Y(n_1377)
);

NAND2xp33_ASAP7_75t_SL g1378 ( 
.A(n_1353),
.B(n_682),
.Y(n_1378)
);

NAND2xp33_ASAP7_75t_SL g1379 ( 
.A(n_1277),
.B(n_71),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1303),
.B(n_71),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1192),
.B(n_1049),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1256),
.B(n_1052),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1287),
.B(n_72),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1288),
.B(n_73),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1241),
.B(n_75),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1300),
.B(n_75),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1198),
.B(n_76),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1265),
.B(n_77),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1237),
.B(n_1322),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1237),
.B(n_78),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1199),
.B(n_81),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1342),
.B(n_1323),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1218),
.B(n_83),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1293),
.B(n_83),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1246),
.B(n_84),
.Y(n_1395)
);

NAND2xp33_ASAP7_75t_SL g1396 ( 
.A(n_1251),
.B(n_85),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1346),
.B(n_86),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1272),
.B(n_87),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1240),
.B(n_88),
.Y(n_1399)
);

NAND2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1252),
.B(n_89),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1273),
.B(n_90),
.Y(n_1401)
);

NAND2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1253),
.B(n_92),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1273),
.B(n_1260),
.Y(n_1403)
);

NAND2xp33_ASAP7_75t_SL g1404 ( 
.A(n_1255),
.B(n_93),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1257),
.B(n_93),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1258),
.B(n_95),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1179),
.B(n_98),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1313),
.B(n_1232),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1212),
.B(n_100),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1184),
.B(n_101),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1259),
.B(n_103),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1238),
.B(n_105),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1229),
.B(n_108),
.Y(n_1413)
);

NAND2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1321),
.B(n_108),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1201),
.B(n_1339),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1339),
.B(n_110),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1267),
.B(n_111),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1182),
.B(n_112),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1324),
.B(n_115),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1268),
.B(n_115),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1324),
.B(n_116),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1305),
.B(n_117),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1189),
.B(n_118),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1269),
.B(n_118),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1305),
.B(n_119),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1270),
.B(n_119),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_SL g1427 ( 
.A(n_1221),
.B(n_120),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1274),
.B(n_123),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1274),
.B(n_125),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1271),
.B(n_126),
.Y(n_1430)
);

NAND2xp33_ASAP7_75t_SL g1431 ( 
.A(n_1262),
.B(n_127),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1183),
.B(n_1333),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1225),
.B(n_137),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1230),
.B(n_138),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1233),
.B(n_141),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1247),
.B(n_145),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1222),
.B(n_146),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1178),
.B(n_147),
.Y(n_1438)
);

NAND2xp33_ASAP7_75t_SL g1439 ( 
.A(n_1318),
.B(n_1302),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1292),
.B(n_150),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_SL g1441 ( 
.A(n_1279),
.B(n_151),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_SL g1442 ( 
.A(n_1281),
.B(n_152),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1347),
.B(n_152),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1325),
.B(n_153),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1215),
.B(n_153),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1207),
.B(n_154),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1349),
.B(n_156),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1343),
.B(n_157),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1282),
.B(n_158),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1294),
.B(n_160),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_SL g1451 ( 
.A(n_1283),
.B(n_161),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1308),
.B(n_162),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1284),
.B(n_163),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1289),
.B(n_164),
.Y(n_1454)
);

NAND2xp33_ASAP7_75t_SL g1455 ( 
.A(n_1290),
.B(n_165),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1180),
.B(n_166),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1335),
.B(n_169),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1208),
.B(n_169),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1249),
.B(n_170),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1209),
.B(n_171),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_SL g1461 ( 
.A(n_1296),
.B(n_174),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1181),
.B(n_174),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1351),
.B(n_175),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1214),
.B(n_176),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1220),
.B(n_179),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1245),
.B(n_1298),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_SL g1467 ( 
.A(n_1298),
.B(n_181),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1186),
.B(n_182),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1185),
.B(n_183),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1223),
.B(n_1187),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1188),
.B(n_1191),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1280),
.B(n_184),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1355),
.B(n_184),
.Y(n_1473)
);

NAND2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1242),
.B(n_185),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1239),
.B(n_187),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1278),
.B(n_189),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1242),
.B(n_193),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1185),
.B(n_193),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1224),
.B(n_195),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_SL g1480 ( 
.A(n_1219),
.B(n_198),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_SL g1481 ( 
.A(n_1236),
.B(n_199),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1306),
.B(n_1236),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1306),
.B(n_1195),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1275),
.B(n_1195),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1275),
.B(n_200),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_SL g1486 ( 
.A(n_1190),
.B(n_200),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1200),
.B(n_201),
.Y(n_1487)
);

NAND2xp33_ASAP7_75t_SL g1488 ( 
.A(n_1334),
.B(n_202),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1200),
.B(n_1202),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1202),
.B(n_1194),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1334),
.B(n_202),
.Y(n_1491)
);

NAND2xp33_ASAP7_75t_SL g1492 ( 
.A(n_1213),
.B(n_204),
.Y(n_1492)
);

NAND2xp33_ASAP7_75t_SL g1493 ( 
.A(n_1213),
.B(n_205),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1336),
.B(n_206),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1217),
.B(n_207),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1337),
.B(n_208),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1248),
.B(n_208),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1304),
.B(n_209),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1203),
.B(n_210),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1196),
.B(n_211),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1337),
.B(n_212),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1228),
.B(n_214),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1228),
.B(n_214),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1341),
.B(n_215),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_SL g1505 ( 
.A(n_1341),
.B(n_216),
.Y(n_1505)
);

AND2x2_ASAP7_75t_SL g1506 ( 
.A(n_1344),
.B(n_217),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1263),
.B(n_1204),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_SL g1508 ( 
.A(n_1344),
.B(n_218),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1217),
.B(n_219),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1295),
.B(n_220),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1231),
.B(n_221),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1263),
.B(n_221),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_SL g1513 ( 
.A(n_1276),
.B(n_222),
.Y(n_1513)
);

NAND2x1p5_ASAP7_75t_L g1514 ( 
.A(n_1327),
.B(n_259),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1243),
.B(n_222),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1250),
.B(n_223),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1317),
.B(n_225),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1316),
.B(n_230),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1216),
.B(n_230),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1216),
.B(n_231),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1254),
.B(n_231),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1276),
.B(n_232),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_SL g1523 ( 
.A(n_1320),
.B(n_233),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1320),
.B(n_234),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1244),
.B(n_234),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1244),
.B(n_235),
.Y(n_1526)
);

NAND2xp33_ASAP7_75t_SL g1527 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1307),
.B(n_1310),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1310),
.B(n_236),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1311),
.B(n_237),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1311),
.B(n_237),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1532)
);

NAND2xp33_ASAP7_75t_SL g1533 ( 
.A(n_1285),
.B(n_1286),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1285),
.B(n_238),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_SL g1535 ( 
.A(n_1286),
.B(n_238),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1329),
.B(n_239),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1312),
.B(n_240),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1329),
.B(n_240),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1312),
.B(n_241),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1345),
.B(n_1348),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1314),
.B(n_244),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1345),
.B(n_1348),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1314),
.B(n_245),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1354),
.B(n_247),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1315),
.B(n_248),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1354),
.B(n_248),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1315),
.B(n_249),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1356),
.B(n_251),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_SL g1549 ( 
.A(n_1356),
.B(n_252),
.Y(n_1549)
);

NAND2xp33_ASAP7_75t_SL g1550 ( 
.A(n_1319),
.B(n_254),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1357),
.B(n_257),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_L g1552 ( 
.A1(n_1528),
.A2(n_258),
.B(n_265),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1364),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1377),
.A2(n_271),
.B(n_272),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1403),
.B(n_1470),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1466),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1483),
.A2(n_279),
.B(n_283),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1361),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1527),
.A2(n_1532),
.B(n_1533),
.C(n_1481),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1365),
.B(n_286),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1389),
.B(n_291),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1415),
.B(n_1507),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1364),
.Y(n_1563)
);

NAND2x1p5_ASAP7_75t_L g1564 ( 
.A(n_1364),
.B(n_292),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1483),
.A2(n_294),
.B(n_297),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1359),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_303),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1439),
.B(n_1461),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1506),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1482),
.A2(n_317),
.A3(n_318),
.B(n_319),
.Y(n_1570)
);

AO32x2_ASAP7_75t_L g1571 ( 
.A1(n_1490),
.A2(n_320),
.A3(n_322),
.B1(n_323),
.B2(n_325),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1495),
.A2(n_330),
.B(n_331),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1543),
.A2(n_337),
.B(n_338),
.C(n_339),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1407),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1407),
.A2(n_1462),
.B(n_1456),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1407),
.B(n_343),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_1456),
.Y(n_1577)
);

AND3x2_ASAP7_75t_L g1578 ( 
.A(n_1495),
.B(n_353),
.C(n_355),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1513),
.A2(n_357),
.B1(n_362),
.B2(n_364),
.Y(n_1579)
);

AO21x1_ASAP7_75t_L g1580 ( 
.A1(n_1494),
.A2(n_1501),
.B(n_1496),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1430),
.B(n_365),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1506),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1392),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1401),
.B(n_381),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1480),
.A2(n_382),
.B(n_383),
.C(n_385),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1456),
.A2(n_388),
.B(n_389),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1522),
.A2(n_390),
.B1(n_391),
.B2(n_394),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1463),
.A2(n_1523),
.B(n_1524),
.C(n_1549),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1459),
.B(n_397),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1509),
.B(n_400),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1509),
.B(n_404),
.Y(n_1591)
);

AO31x2_ASAP7_75t_L g1592 ( 
.A1(n_1478),
.A2(n_405),
.A3(n_408),
.B(n_409),
.Y(n_1592)
);

AOI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1424),
.A2(n_1426),
.B(n_1423),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1358),
.B(n_411),
.Y(n_1594)
);

OA22x2_ASAP7_75t_L g1595 ( 
.A1(n_1519),
.A2(n_412),
.B1(n_413),
.B2(n_416),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1358),
.B(n_419),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1456),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1401),
.Y(n_1598)
);

NOR2xp67_ASAP7_75t_L g1599 ( 
.A(n_1542),
.B(n_1411),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1534),
.A2(n_1535),
.B(n_1512),
.C(n_1505),
.Y(n_1600)
);

OAI22x1_ASAP7_75t_L g1601 ( 
.A1(n_1520),
.A2(n_1547),
.B1(n_1546),
.B2(n_1544),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1419),
.B(n_1421),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1387),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1413),
.B(n_1437),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1387),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1422),
.B(n_1425),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1446),
.A2(n_1420),
.B(n_1417),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1370),
.A2(n_1372),
.B(n_1373),
.Y(n_1609)
);

AOI221x1_ASAP7_75t_L g1610 ( 
.A1(n_1504),
.A2(n_1508),
.B1(n_1492),
.B2(n_1493),
.C(n_1477),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1611)
);

AOI21xp33_ASAP7_75t_L g1612 ( 
.A1(n_1410),
.A2(n_1499),
.B(n_1517),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1525),
.A2(n_1526),
.B(n_1536),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1363),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1368),
.A2(n_1369),
.B(n_1367),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1398),
.B(n_1416),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1391),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1366),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1516),
.A2(n_1497),
.B(n_1515),
.C(n_1511),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1391),
.B(n_1471),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1623)
);

OAI22x1_ASAP7_75t_L g1624 ( 
.A1(n_1529),
.A2(n_1531),
.B1(n_1530),
.B2(n_1537),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1453),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1432),
.B(n_1375),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1539),
.A2(n_1487),
.B(n_1521),
.C(n_1406),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1538),
.A2(n_1479),
.B(n_1541),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1453),
.A2(n_1454),
.B1(n_1428),
.B2(n_1429),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1454),
.B(n_1499),
.Y(n_1630)
);

BUFx8_ASAP7_75t_L g1631 ( 
.A(n_1486),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1510),
.A2(n_1518),
.B(n_1433),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1467),
.B(n_1414),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_L g1634 ( 
.A(n_1485),
.B(n_1500),
.Y(n_1634)
);

OAI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1548),
.A2(n_1541),
.B(n_1538),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1440),
.B(n_1450),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1458),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1460),
.B(n_1464),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1464),
.Y(n_1639)
);

OAI22x1_ASAP7_75t_L g1640 ( 
.A1(n_1502),
.A2(n_1503),
.B1(n_1412),
.B2(n_1548),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1408),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1465),
.A2(n_1384),
.B1(n_1383),
.B2(n_1381),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1405),
.B(n_1445),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1465),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1388),
.B(n_1386),
.Y(n_1645)
);

INVx6_ASAP7_75t_L g1646 ( 
.A(n_1382),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1382),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1474),
.B(n_1400),
.C(n_1404),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1449),
.A2(n_1451),
.B1(n_1455),
.B2(n_1379),
.Y(n_1649)
);

NOR2xp67_ASAP7_75t_L g1650 ( 
.A(n_1457),
.B(n_1476),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1360),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1390),
.B(n_1399),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1397),
.B(n_1452),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1418),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1488),
.A2(n_1491),
.A3(n_1402),
.B(n_1396),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1427),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1447),
.B(n_1393),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1385),
.A2(n_1395),
.B(n_1441),
.C(n_1442),
.Y(n_1659)
);

BUFx2_ASAP7_75t_R g1660 ( 
.A(n_1436),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1448),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1475),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1376),
.Y(n_1663)
);

BUFx10_ASAP7_75t_L g1664 ( 
.A(n_1380),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1394),
.B(n_1409),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1473),
.A2(n_1550),
.B(n_1431),
.C(n_1472),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1378),
.A2(n_1532),
.B(n_1527),
.C(n_1533),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1357),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1371),
.A2(n_1291),
.B(n_1309),
.Y(n_1672)
);

CKINVDCx8_ASAP7_75t_R g1673 ( 
.A(n_1407),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1407),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1357),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1357),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1378),
.A2(n_1357),
.B(n_1377),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1371),
.A2(n_1291),
.B(n_1309),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1543),
.B(n_1545),
.C(n_1549),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1357),
.B(n_1006),
.Y(n_1681)
);

NOR4xp25_ASAP7_75t_L g1682 ( 
.A(n_1519),
.B(n_1520),
.C(n_1489),
.D(n_1540),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1403),
.B(n_1014),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1371),
.A2(n_1291),
.B(n_1309),
.Y(n_1684)
);

AO31x2_ASAP7_75t_L g1685 ( 
.A1(n_1483),
.A2(n_1482),
.A3(n_1478),
.B(n_1438),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1519),
.A2(n_1520),
.B(n_1227),
.C(n_1184),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1687)
);

INVx5_ASAP7_75t_L g1688 ( 
.A(n_1411),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1371),
.A2(n_1291),
.B(n_1309),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1690)
);

AO31x2_ASAP7_75t_L g1691 ( 
.A1(n_1483),
.A2(n_1482),
.A3(n_1478),
.B(n_1438),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1357),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1466),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1374),
.B(n_906),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1403),
.B(n_1014),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1697)
);

O2A1O1Ixp5_ASAP7_75t_L g1698 ( 
.A1(n_1490),
.A2(n_1484),
.B(n_1362),
.C(n_1498),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1357),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1482),
.A2(n_1206),
.B(n_1184),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1514),
.A2(n_1456),
.B(n_1407),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1403),
.B(n_1014),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1357),
.B(n_1234),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1378),
.A2(n_1532),
.B(n_1527),
.C(n_1533),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1357),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1371),
.A2(n_1291),
.B(n_1309),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1675),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1618),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1693),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1669),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1575),
.A2(n_1701),
.B(n_1677),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1673),
.A2(n_1611),
.B1(n_1576),
.B2(n_1574),
.Y(n_1713)
);

NOR2xp67_ASAP7_75t_L g1714 ( 
.A(n_1583),
.B(n_1561),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1687),
.B(n_1683),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1668),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1696),
.B(n_1702),
.Y(n_1718)
);

OAI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1572),
.A2(n_1690),
.B1(n_1697),
.B2(n_1692),
.C(n_1703),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1686),
.A2(n_1588),
.B(n_1593),
.C(n_1600),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1598),
.B(n_1695),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1612),
.A2(n_1630),
.B(n_1613),
.C(n_1700),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1576),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1699),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_L g1725 ( 
.A(n_1561),
.B(n_1688),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1628),
.A2(n_1610),
.B(n_1635),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1681),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1620),
.A2(n_1638),
.B(n_1636),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1705),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1635),
.A2(n_1680),
.B(n_1698),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1631),
.Y(n_1731)
);

OR2x6_ASAP7_75t_L g1732 ( 
.A(n_1681),
.B(n_1576),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1681),
.B(n_1555),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1606),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1551),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1619),
.B(n_1559),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1603),
.B(n_1605),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1621),
.B(n_1672),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1688),
.A2(n_1657),
.B1(n_1694),
.B2(n_1556),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1577),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1629),
.A2(n_1609),
.B(n_1615),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1631),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1552),
.B(n_1648),
.C(n_1572),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_SL g1744 ( 
.A1(n_1670),
.A2(n_1704),
.B(n_1659),
.C(n_1568),
.Y(n_1744)
);

NOR2xp67_ASAP7_75t_L g1745 ( 
.A(n_1601),
.B(n_1640),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1577),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1594),
.A2(n_1596),
.B(n_1597),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1617),
.B(n_1625),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1678),
.B(n_1684),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_R g1750 ( 
.A(n_1664),
.B(n_1651),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1613),
.A2(n_1604),
.B(n_1633),
.C(n_1627),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1567),
.A2(n_1580),
.B(n_1648),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1586),
.B(n_1674),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1558),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1584),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1599),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1639),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1689),
.B(n_1706),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1647),
.Y(n_1759)
);

BUFx4f_ASAP7_75t_SL g1760 ( 
.A(n_1664),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1564),
.Y(n_1761)
);

AOI222xp33_ASAP7_75t_L g1762 ( 
.A1(n_1637),
.A2(n_1644),
.B1(n_1624),
.B2(n_1590),
.C1(n_1591),
.C2(n_1643),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1569),
.A2(n_1582),
.B1(n_1595),
.B2(n_1641),
.Y(n_1763)
);

AOI21xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1682),
.A2(n_1655),
.B(n_1626),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1562),
.B(n_1622),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1649),
.A2(n_1587),
.B1(n_1579),
.B2(n_1602),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1566),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1607),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1685),
.B(n_1691),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1587),
.A2(n_1594),
.B1(n_1596),
.B2(n_1667),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1660),
.B(n_1616),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1645),
.A2(n_1654),
.B1(n_1634),
.B2(n_1666),
.Y(n_1772)
);

BUFx12f_ASAP7_75t_L g1773 ( 
.A(n_1553),
.Y(n_1773)
);

OR2x6_ASAP7_75t_L g1774 ( 
.A(n_1563),
.B(n_1560),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1646),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1563),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1573),
.B(n_1585),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1642),
.A2(n_1632),
.B(n_1608),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1554),
.A2(n_1565),
.B(n_1557),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1634),
.A2(n_1662),
.B1(n_1661),
.B2(n_1653),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1560),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1665),
.B(n_1652),
.Y(n_1782)
);

INVx8_ASAP7_75t_L g1783 ( 
.A(n_1663),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1614),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1589),
.B(n_1581),
.C(n_1650),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1650),
.B(n_1578),
.C(n_1658),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1663),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1691),
.B(n_1571),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1656),
.B(n_1592),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1570),
.B(n_1575),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1671),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1671),
.B(n_1675),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1673),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1623),
.A2(n_1533),
.B1(n_1527),
.B2(n_1532),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1671),
.B(n_1675),
.Y(n_1795)
);

CKINVDCx11_ASAP7_75t_R g1796 ( 
.A(n_1673),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1671),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1575),
.B(n_1701),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1673),
.A2(n_1671),
.B1(n_1675),
.B2(n_1681),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1707),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1719),
.A2(n_1732),
.B1(n_1713),
.B2(n_1723),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1789),
.A2(n_1741),
.B(n_1779),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_R g1803 ( 
.A(n_1796),
.B(n_1707),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1792),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1792),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1709),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1791),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1732),
.Y(n_1808)
);

INVx4_ASAP7_75t_SL g1809 ( 
.A(n_1798),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1798),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1795),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1769),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1798),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1716),
.B(n_1717),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_1731),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1757),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1773),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1722),
.A2(n_1720),
.B(n_1785),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1713),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1718),
.B(n_1715),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1790),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1723),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1724),
.B(n_1729),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1783),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1710),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1736),
.B(n_1756),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1797),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1737),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1754),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1711),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1737),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1783),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1725),
.B(n_1712),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1748),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1712),
.B(n_1745),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1765),
.B(n_1755),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1719),
.A2(n_1794),
.B1(n_1762),
.B2(n_1770),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1733),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1783),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1741),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1740),
.Y(n_1842)
);

BUFx2_ASAP7_75t_SL g1843 ( 
.A(n_1714),
.Y(n_1843)
);

BUFx3_ASAP7_75t_L g1844 ( 
.A(n_1740),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1748),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1788),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1726),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1762),
.A2(n_1770),
.B1(n_1743),
.B2(n_1738),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1743),
.A2(n_1749),
.B1(n_1758),
.B2(n_1721),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1726),
.B(n_1759),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1755),
.B(n_1768),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1782),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1727),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1740),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1752),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1799),
.A2(n_1747),
.B1(n_1781),
.B2(n_1763),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1767),
.B(n_1771),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1784),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1815),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1845),
.B(n_1722),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_R g1861 ( 
.A(n_1836),
.B(n_1750),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1815),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1817),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1820),
.B(n_1734),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1808),
.B(n_1786),
.Y(n_1865)
);

NAND2xp33_ASAP7_75t_R g1866 ( 
.A(n_1836),
.B(n_1793),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1829),
.B(n_1751),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1801),
.B(n_1763),
.Y(n_1868)
);

NAND2xp33_ASAP7_75t_R g1869 ( 
.A(n_1836),
.B(n_1793),
.Y(n_1869)
);

AND2x4_ASAP7_75t_SL g1870 ( 
.A(n_1800),
.B(n_1742),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1809),
.B(n_1774),
.Y(n_1871)
);

XOR2xp5_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1708),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1817),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1807),
.Y(n_1874)
);

XNOR2xp5_ASAP7_75t_L g1875 ( 
.A(n_1820),
.B(n_1776),
.Y(n_1875)
);

NAND2xp33_ASAP7_75t_R g1876 ( 
.A(n_1857),
.B(n_1761),
.Y(n_1876)
);

NAND2xp33_ASAP7_75t_R g1877 ( 
.A(n_1822),
.B(n_1761),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1842),
.B(n_1739),
.Y(n_1878)
);

CKINVDCx8_ASAP7_75t_R g1879 ( 
.A(n_1843),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1825),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1823),
.Y(n_1881)
);

BUFx8_ASAP7_75t_SL g1882 ( 
.A(n_1825),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_R g1883 ( 
.A(n_1840),
.B(n_1760),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1809),
.B(n_1787),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1806),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_R g1886 ( 
.A(n_1822),
.B(n_1730),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_R g1887 ( 
.A(n_1840),
.B(n_1775),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1832),
.B(n_1751),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_R g1889 ( 
.A(n_1833),
.B(n_1746),
.Y(n_1889)
);

NAND2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1838),
.B(n_1739),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_R g1891 ( 
.A(n_1834),
.B(n_1746),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1835),
.B(n_1720),
.Y(n_1892)
);

XNOR2xp5_ASAP7_75t_L g1893 ( 
.A(n_1852),
.B(n_1772),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1830),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1816),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1804),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1812),
.B(n_1764),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_R g1898 ( 
.A(n_1833),
.B(n_1735),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_R g1899 ( 
.A(n_1842),
.B(n_1780),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_R g1900 ( 
.A(n_1844),
.B(n_1854),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_R g1901 ( 
.A(n_1844),
.B(n_1777),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_R g1902 ( 
.A(n_1854),
.B(n_1777),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1809),
.B(n_1753),
.Y(n_1903)
);

NAND2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1848),
.B(n_1778),
.Y(n_1904)
);

XNOR2xp5_ASAP7_75t_L g1905 ( 
.A(n_1849),
.B(n_1805),
.Y(n_1905)
);

INVxp67_ASAP7_75t_SL g1906 ( 
.A(n_1831),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1837),
.B(n_1747),
.Y(n_1907)
);

NAND2xp33_ASAP7_75t_R g1908 ( 
.A(n_1810),
.B(n_1813),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1828),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1853),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1895),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1890),
.A2(n_1868),
.B1(n_1904),
.B2(n_1819),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1881),
.B(n_1850),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1906),
.Y(n_1914)
);

OAI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1879),
.A2(n_1818),
.B1(n_1856),
.B2(n_1744),
.C(n_1843),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1860),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1850),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1860),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1892),
.B(n_1841),
.Y(n_1919)
);

AND2x2_ASAP7_75t_SL g1920 ( 
.A(n_1903),
.B(n_1824),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1884),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1863),
.B(n_1873),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1897),
.B(n_1846),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1897),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1892),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1885),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1877),
.Y(n_1927)
);

NOR2xp67_ASAP7_75t_L g1928 ( 
.A(n_1878),
.B(n_1847),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1864),
.B(n_1802),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1903),
.B(n_1821),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1909),
.B(n_1837),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1867),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1888),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1896),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1888),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1911),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1927),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1927),
.B(n_1898),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1914),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1929),
.B(n_1913),
.Y(n_1940)
);

AND2x4_ASAP7_75t_SL g1941 ( 
.A(n_1921),
.B(n_1871),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1929),
.B(n_1855),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1913),
.B(n_1855),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1921),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1912),
.A2(n_1893),
.B1(n_1905),
.B2(n_1827),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1925),
.B(n_1894),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1917),
.B(n_1802),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1915),
.A2(n_1918),
.B1(n_1916),
.B2(n_1933),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1921),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1921),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1921),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1914),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1930),
.B(n_1821),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1930),
.B(n_1821),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1917),
.B(n_1802),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1946),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1937),
.B(n_1928),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1946),
.B(n_1940),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1939),
.Y(n_1960)
);

NAND2x1_ASAP7_75t_L g1961 ( 
.A(n_1937),
.B(n_1928),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1939),
.Y(n_1962)
);

OR3x2_ASAP7_75t_L g1963 ( 
.A(n_1938),
.B(n_1876),
.C(n_1882),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1948),
.B(n_1916),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1936),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1948),
.B(n_1918),
.Y(n_1966)
);

NOR2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1949),
.B(n_1880),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1940),
.B(n_1923),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1940),
.B(n_1923),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1942),
.B(n_1931),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1939),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1942),
.B(n_1926),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1942),
.B(n_1925),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1938),
.A2(n_1915),
.B(n_1870),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1952),
.B(n_1931),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1952),
.B(n_1926),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1947),
.B(n_1955),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1952),
.B(n_1925),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1943),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1937),
.B(n_1932),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1947),
.B(n_1923),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_R g1982 ( 
.A(n_1963),
.B(n_1883),
.Y(n_1982)
);

AO221x2_ASAP7_75t_L g1983 ( 
.A1(n_1974),
.A2(n_1872),
.B1(n_1803),
.B2(n_1861),
.C(n_1920),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1967),
.B(n_1900),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1964),
.B(n_1859),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1961),
.B(n_1889),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1959),
.A2(n_1891),
.B1(n_1866),
.B2(n_1869),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1959),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1960),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1966),
.B(n_1933),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1972),
.A2(n_1908),
.B1(n_1886),
.B2(n_1951),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1972),
.A2(n_1951),
.B1(n_1949),
.B2(n_1910),
.Y(n_1992)
);

OAI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1976),
.A2(n_1949),
.B1(n_1951),
.B2(n_1944),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1976),
.A2(n_1949),
.B1(n_1951),
.B2(n_1944),
.Y(n_1994)
);

AO221x2_ASAP7_75t_L g1995 ( 
.A1(n_1963),
.A2(n_1922),
.B1(n_1875),
.B2(n_1945),
.C(n_1920),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1958),
.B(n_1901),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1970),
.A2(n_1975),
.B1(n_1979),
.B2(n_1977),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_R g1998 ( 
.A(n_1962),
.B(n_1862),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1998),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1988),
.B(n_1977),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_L g2001 ( 
.A(n_1982),
.B(n_1958),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_L g2002 ( 
.A(n_1987),
.B(n_1958),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1989),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1990),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_SL g2005 ( 
.A1(n_1995),
.A2(n_1920),
.B1(n_1941),
.B2(n_1887),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1985),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_L g2007 ( 
.A(n_1983),
.B(n_1945),
.C(n_1971),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1997),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1992),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1983),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1984),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1986),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1993),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1994),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1991),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1996),
.B(n_1981),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1989),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1988),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_SL g2019 ( 
.A1(n_2010),
.A2(n_1865),
.B(n_1941),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2003),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2003),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1999),
.B(n_1956),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_2007),
.A2(n_1924),
.B1(n_1980),
.B2(n_1957),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2018),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_2018),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2008),
.B(n_1924),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2017),
.Y(n_2027)
);

AOI221xp5_ASAP7_75t_L g2028 ( 
.A1(n_2015),
.A2(n_1980),
.B1(n_1874),
.B2(n_1934),
.C(n_1932),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2000),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2001),
.B(n_1981),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_2011),
.A2(n_1980),
.B(n_1934),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_2005),
.A2(n_1978),
.B1(n_1973),
.B2(n_1968),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2006),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2030),
.B(n_2020),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2021),
.B(n_2009),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2027),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2029),
.B(n_2009),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_2032),
.B(n_2012),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2031),
.B(n_2013),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2033),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2022),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2024),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2019),
.B(n_2002),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2026),
.B(n_2014),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_2025),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2031),
.B(n_2016),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2037),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2045),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2037),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2035),
.Y(n_2050)
);

INVxp33_ASAP7_75t_SL g2051 ( 
.A(n_2035),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2042),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2034),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2045),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2045),
.Y(n_2055)
);

INVx1_ASAP7_75t_SL g2056 ( 
.A(n_2036),
.Y(n_2056)
);

O2A1O1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_2056),
.A2(n_2038),
.B(n_2041),
.C(n_2040),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2048),
.Y(n_2058)
);

AOI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_2051),
.A2(n_2038),
.B1(n_2039),
.B2(n_2046),
.C(n_2044),
.Y(n_2059)
);

OAI221xp5_ASAP7_75t_L g2060 ( 
.A1(n_2047),
.A2(n_2043),
.B1(n_2023),
.B2(n_2032),
.C(n_2046),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2054),
.B(n_2039),
.C(n_2028),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_2051),
.B(n_2026),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_L g2063 ( 
.A(n_2055),
.B(n_2052),
.C(n_2048),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2053),
.B(n_2016),
.C(n_2000),
.D(n_2004),
.Y(n_2064)
);

NOR4xp25_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_2050),
.C(n_2049),
.D(n_2004),
.Y(n_2065)
);

OAI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2059),
.A2(n_1853),
.B1(n_1811),
.B2(n_1978),
.C(n_1858),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_2061),
.A2(n_1826),
.B(n_1969),
.C(n_1968),
.Y(n_2067)
);

NOR3xp33_ASAP7_75t_L g2068 ( 
.A(n_2063),
.B(n_1785),
.C(n_1728),
.Y(n_2068)
);

OAI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2060),
.A2(n_1778),
.B1(n_1950),
.B2(n_1944),
.C(n_1728),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2069),
.B(n_2058),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2066),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_L g2072 ( 
.A(n_2068),
.B(n_2062),
.C(n_2064),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_L g2073 ( 
.A(n_2067),
.B(n_1969),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_R g2074 ( 
.A(n_2071),
.B(n_2065),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_SL g2075 ( 
.A(n_2072),
.B(n_1902),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2075),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2074),
.A2(n_2070),
.B(n_2073),
.C(n_1899),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2076),
.A2(n_1865),
.B1(n_1814),
.B2(n_1953),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2077),
.Y(n_2079)
);

INVxp67_ASAP7_75t_SL g2080 ( 
.A(n_2079),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2080),
.A2(n_2078),
.B1(n_1935),
.B2(n_1932),
.Y(n_2081)
);

OAI222xp33_ASAP7_75t_L g2082 ( 
.A1(n_2081),
.A2(n_1950),
.B1(n_1851),
.B2(n_1935),
.C1(n_1919),
.C2(n_1965),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2082),
.A2(n_1950),
.B1(n_1921),
.B2(n_1935),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2083),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_1941),
.B1(n_1921),
.B2(n_1953),
.C(n_1954),
.Y(n_2085)
);

AOI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_1766),
.B(n_1851),
.C(n_1953),
.Y(n_2086)
);


endmodule