module fake_jpeg_27263_n_11 (n_0, n_2, n_1, n_11);

input n_0;
input n_2;
input n_1;

output n_11;

wire n_3;
wire n_10;
wire n_4;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g3 ( 
.A(n_0),
.Y(n_3)
);

INVx3_ASAP7_75t_L g4 ( 
.A(n_1),
.Y(n_4)
);

INVx3_ASAP7_75t_L g5 ( 
.A(n_1),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_7),
.C(n_8),
.Y(n_9)
);

NOR3xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.C(n_1),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_3),
.Y(n_10)
);

AOI322xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_9),
.C1(n_7),
.C2(n_8),
.Y(n_11)
);


endmodule