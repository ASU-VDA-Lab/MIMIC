module fake_jpeg_22368_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx2_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_20),
.B(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_22),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_17),
.C(n_20),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_48),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_4),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_42),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_70),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.C(n_19),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_41),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_29),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_61),
.B1(n_54),
.B2(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_81),
.B(n_12),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_19),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_14),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_31),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_66),
.C(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_74),
.A3(n_69),
.B1(n_79),
.B2(n_55),
.C1(n_14),
.C2(n_13),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_31),
.Y(n_96)
);

OA21x2_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_30),
.B(n_6),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_87),
.C(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_95),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_34),
.B1(n_50),
.B2(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_98),
.B(n_7),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_4),
.B(n_6),
.Y(n_98)
);

AOI21x1_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_94),
.B(n_8),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_9),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_50),
.Y(n_104)
);


endmodule