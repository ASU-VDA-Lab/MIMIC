module fake_jpeg_12610_n_420 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_420);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_420;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_58),
.B(n_67),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_68),
.Y(n_112)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_20),
.B(n_15),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_14),
.Y(n_74)
);

BUFx6f_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_78),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_91),
.Y(n_118)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_99),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_29),
.B(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_29),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_98),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_101),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_31),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_106),
.Y(n_135)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_47),
.B(n_0),
.CON(n_105),
.SN(n_105)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_107),
.Y(n_174)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_45),
.B(n_40),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_47),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_11),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_117),
.B(n_93),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_43),
.B1(n_51),
.B2(n_41),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_60),
.A2(n_45),
.B1(n_43),
.B2(n_24),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_51),
.B1(n_24),
.B2(n_38),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_51),
.B1(n_24),
.B2(n_38),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_17),
.B1(n_44),
.B2(n_39),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_124),
.A2(n_130),
.B1(n_140),
.B2(n_142),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_72),
.B1(n_87),
.B2(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_125),
.A2(n_139),
.B1(n_152),
.B2(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_44),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_126),
.B(n_172),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_17),
.B1(n_39),
.B2(n_32),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_56),
.A2(n_54),
.B1(n_32),
.B2(n_30),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_131),
.A2(n_153),
.B1(n_157),
.B2(n_164),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_54),
.B1(n_30),
.B2(n_27),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_76),
.B(n_2),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_151),
.B(n_136),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_92),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_101),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_83),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_162),
.B1(n_170),
.B2(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_95),
.A2(n_89),
.B1(n_99),
.B2(n_100),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_96),
.A2(n_105),
.B1(n_69),
.B2(n_62),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_88),
.A2(n_106),
.B1(n_59),
.B2(n_70),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_78),
.A2(n_57),
.B1(n_65),
.B2(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_57),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_65),
.A2(n_53),
.B1(n_42),
.B2(n_37),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_93),
.A2(n_53),
.B1(n_42),
.B2(n_37),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_157),
.B1(n_138),
.B2(n_141),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_179),
.B(n_181),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_118),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_182),
.Y(n_252)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_115),
.B(n_128),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_126),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_206),
.C(n_214),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_112),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_194),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_122),
.B(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_195),
.B(n_202),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_117),
.B(n_137),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_207),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_125),
.B(n_135),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_132),
.B(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_139),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_147),
.B(n_149),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_213),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_219),
.B1(n_221),
.B2(n_173),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx6_ASAP7_75t_SL g273 ( 
.A(n_211),
.Y(n_273)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_156),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_155),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_152),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_141),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_225),
.Y(n_269)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_141),
.A2(n_143),
.B1(n_134),
.B2(n_114),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_143),
.A2(n_114),
.B1(n_163),
.B2(n_178),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_227),
.B1(n_222),
.B2(n_214),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_171),
.A2(n_166),
.B(n_150),
.C(n_155),
.Y(n_224)
);

OR2x2_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_235),
.Y(n_256)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_113),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_226),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_163),
.A2(n_169),
.B1(n_178),
.B2(n_166),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_167),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_136),
.B(n_165),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_159),
.B(n_165),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_159),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_223),
.B1(n_182),
.B2(n_199),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_272),
.B1(n_277),
.B2(n_238),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_171),
.C(n_173),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_247),
.C(n_248),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_188),
.B(n_192),
.C(n_206),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_208),
.A2(n_216),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_185),
.C(n_211),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_267),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_180),
.A2(n_205),
.B1(n_228),
.B2(n_210),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_262),
.A2(n_276),
.B1(n_212),
.B2(n_232),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_185),
.C(n_235),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_219),
.A2(n_183),
.B1(n_189),
.B2(n_190),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_191),
.A2(n_183),
.B1(n_214),
.B2(n_203),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_224),
.A2(n_200),
.B1(n_201),
.B2(n_198),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_281),
.A2(n_286),
.B1(n_291),
.B2(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_186),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_254),
.B(n_230),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_283),
.B(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_197),
.B1(n_236),
.B2(n_233),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_240),
.B(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_289),
.A2(n_271),
.B1(n_242),
.B2(n_274),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_184),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_220),
.B1(n_196),
.B2(n_218),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_225),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_296),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_225),
.B1(n_238),
.B2(n_267),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_256),
.B1(n_245),
.B2(n_276),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_295),
.A2(n_252),
.B1(n_258),
.B2(n_253),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_250),
.B(n_251),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_241),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_298),
.B(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_243),
.B(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_246),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_301),
.B(n_304),
.Y(n_334)
);

BUFx4f_ASAP7_75t_SL g302 ( 
.A(n_273),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_302),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_269),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_264),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_309),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_270),
.B(n_255),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_257),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_252),
.C(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_312),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_291),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_271),
.C(n_249),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_324),
.C(n_327),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_280),
.B1(n_288),
.B2(n_285),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_307),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_329),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_274),
.C(n_275),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_290),
.A2(n_266),
.B(n_279),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_326),
.A2(n_266),
.B(n_279),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_296),
.C(n_295),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_311),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_337),
.B(n_332),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_339),
.B(n_352),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_315),
.A2(n_281),
.B1(n_293),
.B2(n_306),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_353),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_292),
.B(n_306),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_282),
.B1(n_310),
.B2(n_289),
.Y(n_345)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_280),
.B1(n_299),
.B2(n_286),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_354),
.Y(n_372)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_355),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_283),
.B(n_302),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_302),
.B(n_294),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_297),
.B1(n_275),
.B2(n_312),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_316),
.Y(n_356)
);

NOR4xp25_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_330),
.C(n_318),
.D(n_325),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_339),
.A2(n_327),
.B1(n_322),
.B2(n_334),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_362),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_351),
.A2(n_334),
.B1(n_328),
.B2(n_326),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_351),
.A2(n_320),
.B1(n_337),
.B2(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_343),
.B(n_325),
.CI(n_319),
.CON(n_366),
.SN(n_366)
);

AOI322xp5_ASAP7_75t_SL g377 ( 
.A1(n_366),
.A2(n_345),
.A3(n_357),
.B1(n_338),
.B2(n_354),
.C1(n_356),
.C2(n_355),
.Y(n_377)
);

AOI221xp5_ASAP7_75t_L g375 ( 
.A1(n_367),
.A2(n_346),
.B1(n_347),
.B2(n_340),
.C(n_353),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_352),
.A2(n_336),
.B1(n_333),
.B2(n_317),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_330),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_357),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_358),
.B1(n_363),
.B2(n_373),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_377),
.B(n_381),
.Y(n_391)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

BUFx12_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_382),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_365),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_385),
.B1(n_368),
.B2(n_371),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_390),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_367),
.C(n_376),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_359),
.B1(n_373),
.B2(n_360),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_393),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_369),
.C(n_364),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_359),
.C(n_361),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_366),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_374),
.B1(n_382),
.B2(n_379),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_399),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_389),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_398),
.B(n_400),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_379),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_395),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_386),
.A2(n_385),
.B1(n_383),
.B2(n_331),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_388),
.Y(n_403)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_393),
.C(n_391),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_408),
.C(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_401),
.B(n_391),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_406),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_403),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_405),
.B(n_404),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_413),
.Y(n_416)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

AOI221xp5_ASAP7_75t_L g417 ( 
.A1(n_414),
.A2(n_415),
.B1(n_410),
.B2(n_318),
.C(n_344),
.Y(n_417)
);

AOI321xp33_ASAP7_75t_L g418 ( 
.A1(n_417),
.A2(n_341),
.A3(n_349),
.B1(n_416),
.B2(n_378),
.C(n_335),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_418),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_342),
.Y(n_420)
);


endmodule