module fake_ariane_2235_n_1229 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1229);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1229;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1178;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_479;
wire n_836;
wire n_564;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_1152;
wire n_921;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_895;
wire n_583;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_796;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g323 ( 
.A(n_116),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_137),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_153),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_204),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_120),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_176),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_109),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_182),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_25),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_71),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_130),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_164),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_244),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_213),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_181),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_35),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_140),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_114),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_20),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_187),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_52),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_292),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_65),
.Y(n_351)
);

BUFx2_ASAP7_75t_SL g352 ( 
.A(n_122),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_118),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_37),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_174),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_106),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_128),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_219),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_266),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_167),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_7),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_157),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_41),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_17),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_47),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_192),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_216),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_8),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_205),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_193),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_81),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_91),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_129),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_87),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_90),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_26),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_230),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_42),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

INVxp33_ASAP7_75t_R g383 ( 
.A(n_300),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_73),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_61),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_124),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_136),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_224),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_156),
.Y(n_390)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_141),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_165),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_83),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_57),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_7),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_262),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_311),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_98),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_54),
.Y(n_400)
);

BUFx2_ASAP7_75t_SL g401 ( 
.A(n_274),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_173),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_125),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_212),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_131),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_134),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_289),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_158),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_69),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_257),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_238),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_273),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_284),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_1),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_15),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_200),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_306),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_303),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_79),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_171),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_295),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_313),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_170),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_50),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_264),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_100),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_281),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_270),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_294),
.Y(n_431)
);

BUFx8_ASAP7_75t_SL g432 ( 
.A(n_115),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_198),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_145),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_179),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_6),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_283),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_85),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_222),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_11),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_105),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_103),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_151),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_194),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_64),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_99),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_242),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_27),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_14),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_189),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_293),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_40),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_245),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_315),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_14),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_305),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_89),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_163),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_286),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_197),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_77),
.Y(n_461)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_298),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_308),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_220),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_15),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_117),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_104),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_20),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_29),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_183),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_199),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_319),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_82),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_150),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_186),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_113),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_202),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_201),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_33),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_225),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_2),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_49),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_147),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_0),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_301),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_258),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_251),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_282),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_166),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_119),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_195),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_318),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_241),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_86),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_302),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_248),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_177),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_252),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_247),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_304),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_272),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_24),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_254),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_299),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_74),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_5),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_43),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_11),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_18),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_8),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_322),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_277),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_88),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_229),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_45),
.Y(n_515)
);

BUFx5_ASAP7_75t_L g516 ( 
.A(n_108),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_29),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_132),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_263),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_126),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_72),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_149),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_188),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_297),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_175),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_269),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_121),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_237),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_5),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_110),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_209),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_249),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_296),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_255),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_358),
.B(n_36),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_369),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_369),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_353),
.B(n_0),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_479),
.B(n_1),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_360),
.B(n_2),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_369),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_358),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_510),
.Y(n_543)
);

INVxp33_ASAP7_75t_SL g544 ( 
.A(n_345),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_428),
.B(n_471),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_510),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_323),
.B(n_326),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_471),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_328),
.B(n_3),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_486),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_325),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_332),
.B(n_3),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_440),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_4),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_333),
.B(n_4),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_527),
.B(n_6),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_9),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_336),
.B(n_341),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_358),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_425),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_365),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_412),
.B(n_433),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_342),
.B(n_9),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_534),
.B(n_38),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_432),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_425),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_378),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_466),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_346),
.B(n_348),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_466),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_466),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_361),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_465),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_525),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_351),
.B(n_10),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_525),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_502),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_525),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_449),
.B(n_10),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_396),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_368),
.B(n_12),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_450),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_39),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_526),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_517),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_459),
.B(n_12),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_484),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_372),
.B(n_13),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_13),
.Y(n_599)
);

XOR2x2_ASAP7_75t_L g600 ( 
.A(n_383),
.B(n_16),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_330),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_377),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_414),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_355),
.B(n_362),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_381),
.Y(n_606)
);

BUFx12f_ASAP7_75t_L g607 ( 
.A(n_415),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_338),
.B(n_16),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_382),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_370),
.B(n_17),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_435),
.B(n_18),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_334),
.B(n_44),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_386),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_388),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_393),
.B(n_19),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_395),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_373),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_397),
.B(n_19),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_374),
.B(n_21),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_405),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_400),
.B(n_21),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_455),
.B(n_509),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_529),
.B(n_22),
.Y(n_626)
);

BUFx8_ASAP7_75t_L g627 ( 
.A(n_446),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_418),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_421),
.B(n_22),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_423),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_454),
.B(n_23),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_324),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_481),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_430),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_489),
.B(n_23),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_463),
.B(n_24),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_532),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_327),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_437),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_447),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_452),
.B(n_25),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_457),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_470),
.B(n_26),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_387),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

BUFx12f_ASAP7_75t_L g646 ( 
.A(n_329),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_398),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_480),
.B(n_27),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_482),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_483),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_352),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_605),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_546),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_608),
.A2(n_442),
.B1(n_443),
.B2(n_427),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_538),
.A2(n_499),
.B1(n_519),
.B2(n_478),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_547),
.B(n_487),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_625),
.B(n_401),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_613),
.A2(n_495),
.B1(n_501),
.B2(n_488),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_550),
.B(n_462),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_503),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_612),
.A2(n_467),
.B1(n_475),
.B2(n_453),
.Y(n_662)
);

AO22x2_ASAP7_75t_L g663 ( 
.A1(n_540),
.A2(n_514),
.B1(n_520),
.B2(n_504),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_536),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_543),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_556),
.A2(n_512),
.B1(n_402),
.B2(n_404),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_540),
.A2(n_522),
.B1(n_530),
.B2(n_379),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_636),
.A2(n_335),
.B1(n_337),
.B2(n_331),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_559),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_546),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_544),
.A2(n_340),
.B1(n_343),
.B2(n_339),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_539),
.A2(n_626),
.B1(n_633),
.B2(n_624),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_543),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_580),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_558),
.A2(n_347),
.B1(n_349),
.B2(n_344),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_611),
.A2(n_533),
.B1(n_531),
.B2(n_528),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_554),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_586),
.B(n_350),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_639),
.B(n_354),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_621),
.A2(n_524),
.B1(n_523),
.B2(n_521),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_552),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_604),
.B(n_356),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_638),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_621),
.A2(n_518),
.B1(n_359),
.B2(n_515),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_632),
.B(n_357),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_SL g686 ( 
.A1(n_553),
.A2(n_429),
.B1(n_364),
.B2(n_366),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_631),
.A2(n_426),
.B1(n_511),
.B2(n_507),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_631),
.A2(n_635),
.B1(n_554),
.B2(n_599),
.Y(n_688)
);

OA22x2_ASAP7_75t_L g689 ( 
.A1(n_555),
.A2(n_431),
.B1(n_367),
.B2(n_371),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_635),
.A2(n_363),
.B1(n_505),
.B2(n_500),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_580),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_599),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_605),
.B(n_375),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_601),
.A2(n_434),
.B1(n_380),
.B2(n_498),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_581),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_643),
.A2(n_422),
.B1(n_496),
.B2(n_494),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_545),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_376),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_618),
.A2(n_384),
.B1(n_385),
.B2(n_493),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_SL g700 ( 
.A1(n_593),
.A2(n_438),
.B1(n_390),
.B2(n_492),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_581),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_L g703 ( 
.A1(n_647),
.A2(n_389),
.B1(n_392),
.B2(n_491),
.Y(n_703)
);

AND2x2_ASAP7_75t_SL g704 ( 
.A(n_643),
.B(n_394),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_568),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_651),
.B(n_399),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_610),
.A2(n_441),
.B1(n_406),
.B2(n_490),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_591),
.B(n_403),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_641),
.A2(n_439),
.B1(n_485),
.B2(n_477),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_32),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_584),
.Y(n_712)
);

AO22x2_ASAP7_75t_L g713 ( 
.A1(n_583),
.A2(n_560),
.B1(n_572),
.B2(n_549),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_596),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_551),
.A2(n_420),
.B1(n_474),
.B2(n_473),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_576),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_566),
.A2(n_419),
.B1(n_472),
.B2(n_464),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_651),
.B(n_407),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_595),
.B(n_408),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_565),
.A2(n_34),
.B1(n_516),
.B2(n_391),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_585),
.A2(n_417),
.B1(n_461),
.B2(n_456),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_561),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_644),
.B(n_616),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_596),
.B(n_409),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_628),
.A2(n_516),
.B1(n_391),
.B2(n_424),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_628),
.A2(n_516),
.B1(n_391),
.B2(n_424),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_634),
.B(n_410),
.Y(n_727)
);

AO22x2_ASAP7_75t_L g728 ( 
.A1(n_630),
.A2(n_516),
.B1(n_391),
.B2(n_424),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_569),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_644),
.A2(n_411),
.B1(n_451),
.B2(n_445),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_602),
.B(n_413),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_602),
.B(n_416),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_630),
.B(n_444),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_557),
.B(n_391),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_646),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_516),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_598),
.A2(n_424),
.B1(n_48),
.B2(n_51),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_564),
.A2(n_424),
.B1(n_53),
.B2(n_55),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_620),
.A2(n_46),
.B1(n_56),
.B2(n_58),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_590),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_653),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_704),
.B(n_535),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_670),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_657),
.B(n_570),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_674),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_691),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_695),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_702),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_727),
.B(n_542),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_710),
.B(n_607),
.Y(n_751)
);

AOI21x1_ASAP7_75t_L g752 ( 
.A1(n_661),
.A2(n_629),
.B(n_623),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_696),
.B(n_619),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_716),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_741),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_688),
.B(n_606),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_709),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_719),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_686),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_739),
.B(n_535),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_656),
.B(n_600),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_714),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_722),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_711),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_729),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_685),
.B(n_542),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_734),
.B(n_609),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_668),
.B(n_563),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_679),
.B(n_640),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_712),
.Y(n_772)
);

XNOR2xp5_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_648),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_731),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_713),
.B(n_563),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_664),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_665),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_673),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_678),
.B(n_642),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_740),
.B(n_562),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_697),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

XOR2xp5_ASAP7_75t_L g783 ( 
.A(n_662),
.B(n_603),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_681),
.B(n_603),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_724),
.B(n_614),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_732),
.Y(n_786)
);

XNOR2x2_ASAP7_75t_L g787 ( 
.A(n_669),
.B(n_627),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_733),
.B(n_614),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_671),
.B(n_694),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_672),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_683),
.B(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_737),
.B(n_622),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_707),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_682),
.B(n_627),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_622),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_707),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_652),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_725),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_725),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_698),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_726),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_736),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_706),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_726),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_660),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_705),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_680),
.B(n_622),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_723),
.B(n_660),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_728),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_663),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_663),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_718),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_684),
.B(n_637),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_720),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_720),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_666),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_667),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_667),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_687),
.B(n_637),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_677),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_690),
.B(n_615),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_669),
.B(n_617),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_791),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_825),
.B(n_677),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_762),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_772),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_825),
.B(n_692),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_805),
.B(n_717),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_813),
.B(n_617),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_801),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_745),
.B(n_692),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_742),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_790),
.B(n_676),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_788),
.B(n_645),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_801),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_825),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_815),
.B(n_659),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_814),
.B(n_645),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_823),
.B(n_649),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_809),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_774),
.B(n_649),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_744),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_743),
.B(n_738),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_785),
.B(n_650),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_746),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_789),
.B(n_721),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_743),
.B(n_650),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_804),
.B(n_537),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_784),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_747),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_801),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_748),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_802),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_817),
.B(n_541),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_783),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_749),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_770),
.B(n_548),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_824),
.B(n_637),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_752),
.A2(n_715),
.B(n_700),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_768),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_792),
.A2(n_708),
.B(n_675),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_811),
.B(n_779),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_794),
.B(n_730),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_757),
.B(n_569),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_818),
.B(n_535),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_759),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_799),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_820),
.B(n_567),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_800),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_767),
.B(n_766),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_754),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_803),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_755),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_751),
.B(n_699),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_760),
.B(n_571),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_763),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_821),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_753),
.B(n_703),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_767),
.A2(n_567),
.B(n_587),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_765),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_806),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_764),
.B(n_571),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_807),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_769),
.B(n_574),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_776),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_750),
.A2(n_567),
.B(n_587),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_761),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_807),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_773),
.B(n_574),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_758),
.B(n_577),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_808),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_756),
.B(n_655),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_771),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_777),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_778),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_756),
.B(n_587),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_756),
.B(n_577),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_781),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_756),
.B(n_579),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_782),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_807),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_786),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_812),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_793),
.Y(n_907)
);

NAND2x1_ASAP7_75t_SL g908 ( 
.A(n_877),
.B(n_797),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_880),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_848),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_848),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_879),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_892),
.B(n_819),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_832),
.B(n_798),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_865),
.B(n_810),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_879),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_829),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_832),
.B(n_775),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_878),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_836),
.B(n_816),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_856),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_896),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_829),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_843),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_873),
.B(n_760),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_896),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_863),
.B(n_822),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_890),
.B(n_795),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_881),
.B(n_795),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_828),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_884),
.B(n_780),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_839),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_828),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_827),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_878),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_849),
.B(n_831),
.Y(n_937)
);

NAND2x1_ASAP7_75t_SL g938 ( 
.A(n_827),
.B(n_830),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_832),
.B(n_780),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_841),
.B(n_796),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_897),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_897),
.Y(n_942)
);

INVx6_ASAP7_75t_L g943 ( 
.A(n_886),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_841),
.B(n_792),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_841),
.B(n_787),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_866),
.B(n_579),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_898),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_833),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_849),
.B(n_588),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_850),
.B(n_562),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_898),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_862),
.A2(n_846),
.B(n_882),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_895),
.B(n_562),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_886),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_826),
.B(n_573),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_853),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_844),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_833),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_830),
.B(n_842),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_884),
.B(n_588),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_592),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_894),
.B(n_592),
.Y(n_962)
);

BUFx4_ASAP7_75t_SL g963 ( 
.A(n_869),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_852),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_842),
.B(n_891),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_844),
.B(n_573),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_869),
.Y(n_967)
);

BUFx12f_ASAP7_75t_L g968 ( 
.A(n_931),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_934),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_921),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_917),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_967),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_954),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_937),
.B(n_858),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_943),
.Y(n_975)
);

INVx2_ASAP7_75t_R g976 ( 
.A(n_910),
.Y(n_976)
);

INVx5_ASAP7_75t_SL g977 ( 
.A(n_965),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_943),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_964),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_958),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_958),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_911),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_937),
.B(n_930),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_928),
.B(n_844),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_928),
.B(n_850),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_925),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_963),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_919),
.B(n_894),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_912),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_943),
.Y(n_990)
);

BUFx8_ASAP7_75t_L g991 ( 
.A(n_924),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_963),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_945),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_945),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_919),
.B(n_894),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_965),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_929),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_920),
.B(n_842),
.Y(n_998)
);

BUFx6f_ASAP7_75t_SL g999 ( 
.A(n_914),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_965),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_923),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_926),
.B(n_834),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_958),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_939),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_935),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_908),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_939),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_959),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_957),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_938),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_933),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_926),
.B(n_840),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_916),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_970),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_SL g1015 ( 
.A1(n_994),
.A2(n_913),
.B1(n_936),
.B2(n_915),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_982),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_989),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1001),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_SL g1019 ( 
.A1(n_971),
.A2(n_840),
.B1(n_959),
.B2(n_905),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_983),
.B(n_946),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_994),
.A2(n_855),
.B1(n_956),
.B2(n_918),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_993),
.A2(n_855),
.B1(n_918),
.B2(n_947),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_992),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_988),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_985),
.A2(n_936),
.B1(n_846),
.B2(n_950),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_1002),
.A2(n_951),
.B1(n_876),
.B2(n_952),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_1002),
.A2(n_876),
.B1(n_952),
.B2(n_944),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_980),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_989),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_1012),
.A2(n_944),
.B1(n_859),
.B2(n_845),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_980),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_984),
.A2(n_835),
.B1(n_860),
.B2(n_901),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_970),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1013),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1013),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_992),
.Y(n_1036)
);

CKINVDCx11_ASAP7_75t_R g1037 ( 
.A(n_971),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_979),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_974),
.B(n_914),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_972),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_986),
.Y(n_1041)
);

CKINVDCx14_ASAP7_75t_R g1042 ( 
.A(n_986),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1005),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_998),
.A2(n_860),
.B1(n_901),
.B2(n_874),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_997),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1008),
.B(n_959),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1011),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1011),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_973),
.A2(n_933),
.B1(n_940),
.B2(n_904),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_988),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_1005),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_976),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_995),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1019),
.A2(n_997),
.B1(n_999),
.B2(n_1006),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_SL g1055 ( 
.A(n_1047),
.B(n_980),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1020),
.B(n_1009),
.Y(n_1056)
);

INVx5_ASAP7_75t_SL g1057 ( 
.A(n_1028),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1017),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1027),
.B(n_949),
.Y(n_1059)
);

OAI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1039),
.A2(n_972),
.B1(n_995),
.B2(n_1004),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1048),
.B(n_1000),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1030),
.A2(n_949),
.B1(n_977),
.B2(n_1008),
.Y(n_1062)
);

CKINVDCx8_ASAP7_75t_R g1063 ( 
.A(n_1023),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1029),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1015),
.A2(n_999),
.B1(n_1010),
.B2(n_861),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_1033),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1038),
.B(n_1009),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_1027),
.A2(n_861),
.B1(n_1004),
.B2(n_1007),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_1037),
.B(n_991),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_1042),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_1028),
.Y(n_1071)
);

BUFx4f_ASAP7_75t_SL g1072 ( 
.A(n_1041),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1014),
.Y(n_1073)
);

AOI222xp33_ASAP7_75t_L g1074 ( 
.A1(n_1030),
.A2(n_1032),
.B1(n_1044),
.B2(n_1016),
.C1(n_1018),
.C2(n_909),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_1028),
.Y(n_1075)
);

INVx4_ASAP7_75t_SL g1076 ( 
.A(n_1028),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1034),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1029),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1049),
.B(n_975),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1032),
.A2(n_885),
.B(n_955),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1045),
.A2(n_977),
.B1(n_996),
.B2(n_1007),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1044),
.A2(n_977),
.B1(n_996),
.B2(n_987),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_1040),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1025),
.B(n_975),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_1046),
.A2(n_864),
.B1(n_953),
.B2(n_932),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1043),
.B(n_978),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1022),
.A2(n_927),
.B1(n_942),
.B2(n_941),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1022),
.A2(n_922),
.B1(n_953),
.B2(n_847),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1021),
.A2(n_940),
.B1(n_837),
.B2(n_883),
.Y(n_1089)
);

OAI222xp33_ASAP7_75t_L g1090 ( 
.A1(n_1021),
.A2(n_932),
.B1(n_900),
.B2(n_902),
.C1(n_888),
.C2(n_903),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_SL g1091 ( 
.A(n_1031),
.B(n_980),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1026),
.A2(n_864),
.B1(n_966),
.B2(n_857),
.Y(n_1092)
);

OAI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_1074),
.A2(n_1066),
.B(n_1080),
.C(n_1073),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1074),
.A2(n_1026),
.B1(n_857),
.B2(n_1046),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1062),
.A2(n_857),
.B1(n_867),
.B2(n_1051),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1082),
.A2(n_1035),
.B1(n_838),
.B2(n_833),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1062),
.A2(n_1082),
.B1(n_1059),
.B2(n_1079),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1069),
.A2(n_1036),
.B(n_1042),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1059),
.A2(n_1052),
.B(n_1031),
.Y(n_1099)
);

OAI221xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1065),
.A2(n_887),
.B1(n_867),
.B2(n_955),
.C(n_893),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1085),
.A2(n_1053),
.B1(n_1024),
.B2(n_1050),
.C(n_969),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1088),
.A2(n_1035),
.B1(n_838),
.B2(n_833),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1068),
.A2(n_1053),
.B1(n_1050),
.B2(n_1024),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1056),
.B(n_1031),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1061),
.B(n_1031),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1092),
.A2(n_838),
.B1(n_854),
.B2(n_976),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1054),
.A2(n_854),
.B1(n_907),
.B2(n_868),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1084),
.B(n_991),
.C(n_1052),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1089),
.A2(n_854),
.B1(n_907),
.B2(n_868),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1087),
.A2(n_854),
.B1(n_907),
.B2(n_868),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1067),
.A2(n_851),
.B1(n_875),
.B2(n_870),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1058),
.A2(n_948),
.B1(n_871),
.B2(n_899),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1055),
.A2(n_968),
.B1(n_871),
.B2(n_969),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1077),
.A2(n_948),
.B1(n_871),
.B2(n_906),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1060),
.A2(n_906),
.B1(n_875),
.B2(n_870),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_1090),
.A2(n_990),
.B1(n_978),
.B2(n_1003),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1064),
.A2(n_906),
.B1(n_872),
.B2(n_990),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1070),
.A2(n_1003),
.B1(n_962),
.B2(n_961),
.Y(n_1118)
);

AOI222xp33_ASAP7_75t_L g1119 ( 
.A1(n_1072),
.A2(n_889),
.B1(n_872),
.B2(n_961),
.C1(n_960),
.C2(n_962),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1078),
.A2(n_981),
.B1(n_960),
.B2(n_594),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1081),
.A2(n_981),
.B1(n_594),
.B2(n_589),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1086),
.A2(n_594),
.B1(n_589),
.B2(n_582),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1083),
.A2(n_589),
.B1(n_582),
.B2(n_573),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1057),
.A2(n_582),
.B1(n_60),
.B2(n_62),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1057),
.A2(n_1091),
.B1(n_1075),
.B2(n_1071),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1071),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1075),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1057),
.B(n_67),
.Y(n_1128)
);

OAI221xp5_ASAP7_75t_L g1129 ( 
.A1(n_1093),
.A2(n_1100),
.B1(n_1097),
.B2(n_1123),
.C(n_1108),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1094),
.A2(n_1063),
.B1(n_1076),
.B2(n_75),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1094),
.A2(n_1076),
.B1(n_70),
.B2(n_76),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1098),
.A2(n_1076),
.B(n_78),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1119),
.B(n_68),
.C(n_80),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_L g1134 ( 
.A(n_1099),
.B(n_84),
.C(n_92),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1127),
.B(n_93),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1095),
.A2(n_94),
.B(n_95),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1118),
.B(n_321),
.Y(n_1138)
);

OAI221xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1095),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.C(n_102),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1101),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1096),
.B(n_107),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1128),
.B(n_316),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1122),
.B(n_111),
.C(n_112),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_SL g1144 ( 
.A(n_1124),
.B(n_123),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1125),
.B(n_312),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1106),
.B(n_127),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1116),
.B(n_310),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1126),
.A2(n_1115),
.B(n_1111),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1103),
.B(n_1102),
.Y(n_1149)
);

OAI221xp5_ASAP7_75t_L g1150 ( 
.A1(n_1113),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.C(n_142),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1107),
.B(n_1111),
.Y(n_1151)
);

OAI221xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1109),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.C(n_148),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1114),
.B(n_152),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1133),
.B(n_1120),
.C(n_1121),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1135),
.B(n_1110),
.Y(n_1155)
);

OAI211xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1132),
.A2(n_1112),
.B(n_1117),
.C(n_159),
.Y(n_1156)
);

OAI211xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1129),
.A2(n_154),
.B(n_155),
.C(n_160),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1136),
.B(n_161),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1149),
.B(n_162),
.Y(n_1159)
);

NOR4xp75_ASAP7_75t_L g1160 ( 
.A(n_1130),
.B(n_168),
.C(n_169),
.D(n_172),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1142),
.Y(n_1161)
);

AOI211x1_ASAP7_75t_L g1162 ( 
.A1(n_1148),
.A2(n_178),
.B(n_180),
.C(n_184),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_1140),
.B(n_185),
.C(n_190),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1140),
.B(n_191),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_196),
.C(n_203),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1155),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1161),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1165),
.B(n_1151),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1159),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1158),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1164),
.B(n_1145),
.Y(n_1171)
);

NAND4xp75_ASAP7_75t_L g1172 ( 
.A(n_1162),
.B(n_1147),
.C(n_1138),
.D(n_1153),
.Y(n_1172)
);

NAND4xp75_ASAP7_75t_L g1173 ( 
.A(n_1160),
.B(n_1146),
.C(n_1141),
.D(n_1144),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1154),
.B(n_1134),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1163),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1166),
.Y(n_1176)
);

XOR2x2_ASAP7_75t_L g1177 ( 
.A(n_1172),
.B(n_1139),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1170),
.B(n_1156),
.Y(n_1178)
);

XOR2x2_ASAP7_75t_L g1179 ( 
.A(n_1168),
.B(n_1139),
.Y(n_1179)
);

XOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1173),
.B(n_1131),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_SL g1181 ( 
.A(n_1170),
.B(n_1152),
.Y(n_1181)
);

XOR2xp5_ASAP7_75t_L g1182 ( 
.A(n_1174),
.B(n_1143),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1178),
.A2(n_1168),
.B1(n_1175),
.B2(n_1171),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1181),
.A2(n_1175),
.B1(n_1169),
.B2(n_1144),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1182),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1176),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1179),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1180),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1177),
.Y(n_1189)
);

XOR2x2_ASAP7_75t_L g1190 ( 
.A(n_1179),
.B(n_1152),
.Y(n_1190)
);

OA22x2_ASAP7_75t_L g1191 ( 
.A1(n_1182),
.A2(n_1169),
.B1(n_1167),
.B2(n_1157),
.Y(n_1191)
);

AOI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1180),
.A2(n_1150),
.B1(n_207),
.B2(n_208),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1186),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1183),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1185),
.Y(n_1195)
);

INVxp33_ASAP7_75t_SL g1196 ( 
.A(n_1189),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1184),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1187),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1193),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1195),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1194),
.A2(n_1188),
.B(n_1190),
.C(n_1191),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1198),
.Y(n_1202)
);

AOI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1197),
.A2(n_1192),
.B1(n_210),
.B2(n_211),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1196),
.B(n_1192),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1201),
.A2(n_1196),
.B1(n_214),
.B2(n_217),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1201),
.A2(n_206),
.B1(n_218),
.B2(n_221),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1200),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1202),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1205),
.A2(n_1199),
.B1(n_1204),
.B2(n_1203),
.C(n_228),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1207),
.B(n_223),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1208),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1211),
.A2(n_1206),
.B1(n_227),
.B2(n_231),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1210),
.Y(n_1213)
);

INVxp67_ASAP7_75t_L g1214 ( 
.A(n_1209),
.Y(n_1214)
);

NOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1213),
.B(n_226),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1212),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1216),
.Y(n_1217)
);

AO22x2_ASAP7_75t_L g1218 ( 
.A1(n_1217),
.A2(n_1214),
.B1(n_1215),
.B2(n_234),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1217),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.C(n_236),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1218),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1219),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1220),
.A2(n_309),
.B1(n_240),
.B2(n_246),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1221),
.A2(n_239),
.B1(n_253),
.B2(n_256),
.Y(n_1223)
);

AO22x1_ASAP7_75t_L g1224 ( 
.A1(n_1221),
.A2(n_259),
.B1(n_261),
.B2(n_265),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1224),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_1223),
.B1(n_1222),
.B2(n_271),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1226),
.Y(n_1227)
);

AOI221xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_267),
.B1(n_268),
.B2(n_275),
.C(n_276),
.Y(n_1228)
);

AOI211xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_278),
.B(n_279),
.C(n_280),
.Y(n_1229)
);


endmodule