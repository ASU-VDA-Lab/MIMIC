module fake_jpeg_21728_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_49),
.B1(n_42),
.B2(n_48),
.Y(n_73)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_82),
.B1(n_91),
.B2(n_48),
.Y(n_105)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_46),
.B(n_18),
.C(n_17),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_76),
.B(n_102),
.C(n_29),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_18),
.B(n_36),
.C(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx5_ASAP7_75t_SL g113 ( 
.A(n_89),
.Y(n_113)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_28),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_124)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_100),
.C(n_49),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_101),
.B1(n_103),
.B2(n_20),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_27),
.A3(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_34),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_30),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_110),
.B(n_24),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_59),
.C(n_41),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_77),
.C(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_87),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_39),
.B(n_41),
.C(n_43),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_121),
.B(n_131),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_18),
.B1(n_36),
.B2(n_45),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_123),
.B1(n_134),
.B2(n_23),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_36),
.B(n_44),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_27),
.B1(n_29),
.B2(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_10),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NOR4xp25_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_9),
.C(n_16),
.D(n_14),
.Y(n_132)
);

NAND2xp67_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_12),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_23),
.B1(n_22),
.B2(n_30),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_135),
.B(n_138),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_93),
.B1(n_98),
.B2(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_148),
.B1(n_122),
.B2(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_141),
.A2(n_145),
.B1(n_150),
.B2(n_155),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_72),
.B1(n_22),
.B2(n_71),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_159),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_72),
.B1(n_99),
.B2(n_85),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_40),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_107),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_127),
.B1(n_121),
.B2(n_131),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_12),
.C(n_16),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_14),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_160),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_131),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_158),
.C(n_31),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_24),
.B1(n_31),
.B2(n_35),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_35),
.B1(n_31),
.B2(n_10),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_113),
.B1(n_114),
.B2(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_31),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_13),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_179),
.B1(n_187),
.B2(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_107),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_168),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_140),
.B(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_174),
.B1(n_153),
.B2(n_115),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_122),
.B1(n_129),
.B2(n_108),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_166),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_178),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_133),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_114),
.B1(n_130),
.B2(n_118),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_37),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_156),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_85),
.B(n_77),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_188),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_115),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_136),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_13),
.B1(n_11),
.B2(n_8),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_212),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_214),
.B(n_216),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_200),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_159),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_218),
.B(n_226),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_88),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_161),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_0),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_225),
.B1(n_165),
.B2(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_153),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_168),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_177),
.B(n_184),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_115),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_184),
.B1(n_177),
.B2(n_11),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_115),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_244),
.B(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_175),
.C(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_236),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_190),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_235),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_194),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_171),
.C(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_198),
.B1(n_217),
.B2(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_169),
.B(n_193),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_197),
.B(n_220),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_184),
.B(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_171),
.C(n_187),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_184),
.C(n_169),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_207),
.A2(n_11),
.B1(n_8),
.B2(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_253),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_224),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_202),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_254),
.A2(n_264),
.B1(n_236),
.B2(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_255),
.B(n_258),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_206),
.B1(n_203),
.B2(n_210),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_211),
.B(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_205),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_239),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_205),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_243),
.B1(n_245),
.B2(n_203),
.Y(n_289)
);

OR2x6_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_206),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_250),
.C(n_232),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_281),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_250),
.C(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_233),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_285),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_288),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_237),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_259),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_230),
.B1(n_216),
.B2(n_214),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_292),
.B1(n_275),
.B2(n_263),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_240),
.B1(n_237),
.B2(n_225),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_299),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_277),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_263),
.B1(n_256),
.B2(n_271),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_276),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_305),
.C(n_307),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_258),
.B1(n_275),
.B2(n_270),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_306),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_262),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_281),
.A2(n_275),
.B1(n_255),
.B2(n_267),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_308),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_279),
.C(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_317),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_298),
.B(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_285),
.C(n_284),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_288),
.C(n_252),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_310),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_295),
.B1(n_304),
.B2(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_297),
.B1(n_306),
.B2(n_278),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_329),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_325),
.B(n_312),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_300),
.B1(n_253),
.B2(n_5),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_311),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_313),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_6),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_324),
.B(n_320),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_326),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_332),
.Y(n_339)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_338),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_334),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_337),
.B(n_330),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_321),
.C(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_329),
.Y(n_345)
);

FAx1_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_7),
.CI(n_333),
.CON(n_346),
.SN(n_346)
);


endmodule