module real_jpeg_15232_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI21xp33_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_9),
.B(n_10),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_1),
.B(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_2),
.B(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

OR2x4_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_13),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_5),
.B(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NAND5xp2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_28),
.C(n_33),
.D(n_41),
.E(n_44),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

AND2x4_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_45),
.B(n_46),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

AOI22x1_ASAP7_75t_R g41 ( 
.A1(n_34),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);


endmodule