module fake_jpeg_17772_n_155 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_155);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_4),
.B(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_13),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_35),
.B(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_22),
.Y(n_73)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_43),
.B1(n_44),
.B2(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_21),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_21),
.A2(n_8),
.B1(n_10),
.B2(n_19),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_10),
.B(n_30),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_26),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_52),
.B1(n_18),
.B2(n_16),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_63),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_24),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_73),
.B(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_25),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_33),
.B(n_40),
.Y(n_81)
);

OAI22x1_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_99),
.B1(n_96),
.B2(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_63),
.B1(n_64),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_85),
.B1(n_96),
.B2(n_75),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_58),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_53),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_92),
.C(n_75),
.Y(n_104)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_56),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AO21x2_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_50),
.B(n_66),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_54),
.B1(n_73),
.B2(n_58),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_70),
.B1(n_69),
.B2(n_75),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_56),
.B1(n_84),
.B2(n_92),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_114),
.B(n_86),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_87),
.C(n_99),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_100),
.B1(n_90),
.B2(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_115),
.B1(n_102),
.B2(n_108),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_89),
.B1(n_97),
.B2(n_83),
.Y(n_114)
);

NAND2x1_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_91),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_86),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_131),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_136),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_131),
.C(n_133),
.Y(n_144)
);

AO221x1_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_115),
.B1(n_105),
.B2(n_111),
.C(n_112),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_127),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_142),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_101),
.B1(n_126),
.B2(n_117),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_138),
.C(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_126),
.C(n_142),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_130),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_137),
.B(n_112),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_152),
.B(n_149),
.Y(n_155)
);


endmodule