module fake_jpeg_16105_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_19),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_14),
.B1(n_9),
.B2(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_22),
.B1(n_21),
.B2(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_34),
.CI(n_18),
.CON(n_38),
.SN(n_38)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_30),
.C(n_26),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_28),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_38),
.C(n_26),
.Y(n_47)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_42),
.A3(n_38),
.B1(n_39),
.B2(n_33),
.C1(n_20),
.C2(n_17),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_27),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_21),
.C(n_29),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_29),
.Y(n_50)
);


endmodule