module fake_jpeg_4669_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_26),
.B(n_7),
.CON(n_42),
.SN(n_42)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_42),
.B(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_46),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_7),
.B(n_11),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_0),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_20),
.B1(n_34),
.B2(n_35),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_8),
.Y(n_92)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_74),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_76),
.B(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_37),
.B1(n_29),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_28),
.B1(n_30),
.B2(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_61),
.B1(n_58),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_21),
.B1(n_31),
.B2(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_33),
.B1(n_31),
.B2(n_21),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_33),
.B1(n_31),
.B2(n_3),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_105),
.C(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_8),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_8),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_33),
.B1(n_31),
.B2(n_9),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_39),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_47),
.A2(n_33),
.B1(n_6),
.B2(n_4),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_4),
.B1(n_11),
.B2(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_4),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_40),
.B(n_0),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_39),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_89),
.Y(n_147)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_48),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_72),
.B(n_69),
.Y(n_148)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_119),
.Y(n_151)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_71),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_130),
.Y(n_166)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_89),
.Y(n_129)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_48),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_133),
.A2(n_68),
.B1(n_112),
.B2(n_98),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_55),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_138),
.Y(n_173)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_107),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_1),
.C(n_3),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_138),
.C(n_116),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_80),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_148),
.A2(n_174),
.B(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_150),
.Y(n_193)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_152),
.B(n_130),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_155),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_99),
.B1(n_85),
.B2(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_177),
.B1(n_119),
.B2(n_128),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_89),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_175),
.C(n_176),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_149),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_84),
.C(n_78),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_125),
.C(n_144),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_71),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_83),
.B(n_89),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_65),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_77),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_117),
.A2(n_99),
.B1(n_68),
.B2(n_85),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_131),
.B(n_88),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_75),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_123),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_174),
.B(n_175),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_191),
.B(n_208),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_195),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_132),
.B1(n_117),
.B2(n_137),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_197),
.B1(n_198),
.B2(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_136),
.B1(n_139),
.B2(n_115),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_194),
.A2(n_196),
.B1(n_183),
.B2(n_157),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_163),
.B1(n_177),
.B2(n_167),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_136),
.B1(n_115),
.B2(n_73),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_205),
.C(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_204),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_127),
.C(n_97),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_140),
.B1(n_135),
.B2(n_128),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_145),
.B(n_135),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_168),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_120),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_123),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_171),
.B(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_238),
.Y(n_250)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_222),
.Y(n_256)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_224),
.C(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_188),
.B(n_150),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_234),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_162),
.B(n_183),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_202),
.B(n_215),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_205),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_245),
.B1(n_217),
.B2(n_201),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_157),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_184),
.C(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_193),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_185),
.A2(n_194),
.B1(n_190),
.B2(n_208),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_198),
.A2(n_197),
.B1(n_206),
.B2(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_200),
.B1(n_195),
.B2(n_189),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_215),
.B(n_199),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_268),
.B1(n_267),
.B2(n_230),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_268),
.B(n_269),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_242),
.B1(n_229),
.B2(n_223),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_237),
.B1(n_228),
.B2(n_239),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_184),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_265),
.C(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_187),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_192),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_230),
.B(n_232),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_271),
.A2(n_275),
.B(n_263),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_250),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_286),
.C(n_265),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_249),
.A2(n_220),
.B1(n_229),
.B2(n_252),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_285),
.A2(n_260),
.B1(n_248),
.B2(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_251),
.C(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_291),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_251),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_284),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_262),
.CI(n_258),
.CON(n_293),
.SN(n_293)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_293),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_300),
.C(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_298),
.B1(n_275),
.B2(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_248),
.B1(n_247),
.B2(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_255),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_270),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_264),
.C(n_285),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_275),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_303),
.C(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_271),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_308),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_283),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_277),
.C(n_276),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_293),
.B(n_297),
.C(n_298),
.D(n_300),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_273),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_281),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_290),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_304),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_326),
.B(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_306),
.C(n_304),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_293),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.C(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_324),
.B(n_315),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_325),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_322),
.B(n_326),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.C(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_282),
.C(n_289),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_264),
.Y(n_336)
);


endmodule