module fake_netlist_6_1309_n_470 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_470);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_470;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_464;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_26),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_50),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_32),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_35),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_52),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_49),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_34),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_48),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_45),
.B(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_71),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_13),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_23),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_33),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_78),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_39),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_41),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_90),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_55),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_27),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_25),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_44),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_63),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_105),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_66),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_64),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_0),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_0),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_2),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_174),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_151),
.B(n_3),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_11),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_4),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_135),
.B(n_5),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_6),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_7),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_8),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_8),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_9),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_136),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_9),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_10),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_184),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_199),
.B1(n_142),
.B2(n_143),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_184),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_139),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_140),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_179),
.B1(n_149),
.B2(n_180),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_202),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_225),
.B(n_203),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_10),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_163),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

BUFx4f_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_141),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_231),
.B(n_170),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_163),
.C(n_148),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_157),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_215),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_154),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_214),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_221),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_254),
.B(n_207),
.Y(n_291)
);

OR2x6_ASAP7_75t_SL g292 ( 
.A(n_254),
.B(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_243),
.B(n_222),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_243),
.B(n_214),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_265),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_226),
.B(n_232),
.Y(n_297)
);

NAND2x1p5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_144),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_223),
.B(n_241),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_223),
.B1(n_235),
.B2(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_242),
.A2(n_239),
.B1(n_145),
.B2(n_146),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_246),
.B(n_155),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_246),
.B(n_238),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_238),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_239),
.B1(n_178),
.B2(n_147),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_167),
.B1(n_193),
.B2(n_172),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_260),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_291),
.A2(n_269),
.B(n_251),
.C(n_249),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_300),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_SL g327 ( 
.A1(n_295),
.A2(n_189),
.B(n_153),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_286),
.Y(n_328)
);

OAI31xp33_ASAP7_75t_SL g329 ( 
.A1(n_288),
.A2(n_181),
.A3(n_158),
.B(n_159),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_244),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_250),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_293),
.A2(n_152),
.B(n_171),
.C(n_168),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

BUFx2_ASAP7_75t_SL g334 ( 
.A(n_294),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_285),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_245),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_310),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_228),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_301),
.A2(n_188),
.B(n_162),
.C(n_164),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_161),
.Y(n_345)
);

BUFx4f_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_296),
.A2(n_253),
.B(n_191),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_319),
.A2(n_165),
.B(n_166),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_196),
.B1(n_185),
.B2(n_201),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

BUFx8_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_173),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_278),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_294),
.B(n_278),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_294),
.Y(n_358)
);

AOI221xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_320),
.B1(n_307),
.B2(n_200),
.C(n_198),
.Y(n_359)
);

AO21x2_ASAP7_75t_L g360 ( 
.A1(n_337),
.A2(n_304),
.B(n_305),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_326),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_298),
.B(n_284),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_350),
.A2(n_283),
.B(n_314),
.Y(n_363)
);

AO31x2_ASAP7_75t_L g364 ( 
.A1(n_349),
.A2(n_344),
.A3(n_345),
.B(n_352),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_302),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_186),
.B(n_183),
.Y(n_367)
);

CKINVDCx6p67_ASAP7_75t_R g368 ( 
.A(n_334),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_313),
.B(n_306),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_313),
.C(n_306),
.Y(n_370)
);

AO32x2_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_323),
.A3(n_328),
.B1(n_342),
.B2(n_357),
.Y(n_371)
);

OR3x4_ASAP7_75t_SL g372 ( 
.A(n_327),
.B(n_14),
.C(n_17),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_325),
.A2(n_306),
.B(n_302),
.Y(n_373)
);

AO21x2_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_125),
.B(n_20),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_SL g376 ( 
.A1(n_341),
.A2(n_124),
.B(n_21),
.C(n_22),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_336),
.Y(n_378)
);

OAI21x1_ASAP7_75t_SL g379 ( 
.A1(n_348),
.A2(n_18),
.B(n_24),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_354),
.A2(n_31),
.B(n_36),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_37),
.B(n_38),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_331),
.A2(n_40),
.B(n_43),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_346),
.B(n_338),
.C(n_322),
.Y(n_385)
);

OAI221xp5_ASAP7_75t_L g386 ( 
.A1(n_367),
.A2(n_346),
.B1(n_332),
.B2(n_356),
.C(n_323),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_353),
.B1(n_355),
.B2(n_351),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_372),
.A2(n_351),
.B1(n_355),
.B2(n_51),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_384),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_377),
.A2(n_58),
.B1(n_65),
.B2(n_67),
.Y(n_391)
);

OAI211xp5_ASAP7_75t_SL g392 ( 
.A1(n_384),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_358),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_393)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_79),
.B(n_81),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_372),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_87),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_370),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_378),
.A2(n_108),
.B(n_109),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_361),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_398),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

NAND2x1_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_375),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_371),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_371),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_401),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_363),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_364),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_371),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_364),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_360),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_360),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_374),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_374),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_415),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_399),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

OR2x6_ASAP7_75t_SL g431 ( 
.A(n_414),
.B(n_390),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_407),
.A2(n_379),
.B1(n_383),
.B2(n_382),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_420),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_416),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_416),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_410),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_408),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_408),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_410),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_410),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_407),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_415),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_381),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_423),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_422),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_415),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_446),
.B(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_443),
.B(n_447),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_428),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_441),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_446),
.Y(n_452)
);

O2A1O1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_450),
.A2(n_436),
.B(n_440),
.C(n_376),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_434),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_449),
.A2(n_406),
.B(n_365),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_454),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_452),
.Y(n_458)
);

AOI211xp5_ASAP7_75t_L g459 ( 
.A1(n_456),
.A2(n_455),
.B(n_451),
.C(n_445),
.Y(n_459)
);

OAI321xp33_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_439),
.A3(n_442),
.B1(n_437),
.B2(n_438),
.C(n_434),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_444),
.Y(n_461)
);

AOI32xp33_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_438),
.A3(n_435),
.B1(n_432),
.B2(n_444),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_444),
.C(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_464),
.B(n_462),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_465),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

AOI222xp33_ASAP7_75t_SL g468 ( 
.A1(n_467),
.A2(n_112),
.B1(n_113),
.B2(n_121),
.C1(n_122),
.C2(n_123),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_369),
.B(n_373),
.Y(n_470)
);


endmodule