module real_aes_8121_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_364;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_892;
wire n_528;
wire n_578;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_938;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_996;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_922;
wire n_633;
wire n_679;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_719;
wire n_967;
wire n_465;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_968;
wire n_650;
wire n_710;
wire n_646;
wire n_743;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_0), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_1), .A2(n_147), .B1(n_398), .B2(n_402), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_2), .A2(n_152), .B1(n_544), .B2(n_602), .Y(n_936) );
INVx1_ASAP7_75t_L g776 ( .A(n_3), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_4), .A2(n_305), .B1(n_428), .B2(n_432), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_5), .A2(n_118), .B1(n_402), .B2(n_853), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_6), .Y(n_758) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_7), .A2(n_174), .B1(n_265), .B2(n_451), .C1(n_455), .C2(n_504), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_8), .A2(n_85), .B1(n_397), .B2(n_401), .Y(n_396) );
AO22x2_ASAP7_75t_L g358 ( .A1(n_9), .A2(n_199), .B1(n_359), .B2(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g979 ( .A(n_9), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_10), .A2(n_137), .B1(n_417), .B2(n_481), .Y(n_987) );
AOI222xp33_ASAP7_75t_L g877 ( .A1(n_11), .A2(n_286), .B1(n_296), .B2(n_354), .C1(n_454), .C2(n_456), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_12), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_13), .A2(n_42), .B1(n_791), .B2(n_793), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_14), .A2(n_112), .B1(n_498), .B2(n_668), .Y(n_904) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_15), .A2(n_103), .B1(n_476), .B2(n_477), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_16), .A2(n_255), .B1(n_454), .B2(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g963 ( .A(n_17), .Y(n_963) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_18), .A2(n_177), .B1(n_600), .B2(n_602), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_19), .A2(n_233), .B1(n_421), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_20), .A2(n_76), .B1(n_454), .B2(n_456), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_21), .A2(n_188), .B1(n_416), .B2(n_421), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_22), .A2(n_178), .B1(n_458), .B2(n_503), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_23), .A2(n_94), .B1(n_427), .B2(n_470), .C(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_24), .A2(n_140), .B1(n_409), .B2(n_550), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_25), .A2(n_281), .B1(n_793), .B2(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_26), .A2(n_96), .B1(n_486), .B2(n_868), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_27), .A2(n_121), .B1(n_407), .B2(n_412), .Y(n_406) );
AO22x2_ASAP7_75t_L g362 ( .A1(n_28), .A2(n_102), .B1(n_359), .B2(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_29), .A2(n_240), .B1(n_417), .B2(n_549), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g995 ( .A1(n_30), .A2(n_176), .B1(n_264), .B2(n_458), .C1(n_658), .C2(n_775), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_31), .B(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_32), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_33), .A2(n_232), .B1(n_409), .B2(n_767), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_34), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_35), .A2(n_186), .B1(n_584), .B2(n_585), .C(n_586), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_36), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_37), .A2(n_104), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_38), .A2(n_160), .B1(n_430), .B2(n_574), .Y(n_909) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_39), .A2(n_113), .B1(n_658), .B2(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_40), .B(n_379), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_41), .A2(n_81), .B1(n_549), .B2(n_638), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_43), .A2(n_128), .B1(n_486), .B2(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g664 ( .A(n_44), .Y(n_664) );
AOI22x1_ASAP7_75t_L g676 ( .A1(n_45), .A2(n_677), .B1(n_710), .B2(n_711), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_45), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_46), .A2(n_70), .B1(n_416), .B2(n_602), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_47), .A2(n_91), .B1(n_639), .B2(n_808), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_48), .A2(n_250), .B1(n_650), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_49), .A2(n_205), .B1(n_549), .B2(n_671), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_50), .A2(n_78), .B1(n_764), .B2(n_816), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_51), .A2(n_275), .B1(n_573), .B2(n_671), .Y(n_961) );
INVx1_ASAP7_75t_L g581 ( .A(n_52), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_53), .A2(n_170), .B1(n_401), .B2(n_464), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_54), .A2(n_67), .B1(n_462), .B2(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g640 ( .A(n_55), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_56), .B(n_462), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_57), .A2(n_333), .B1(n_427), .B2(n_430), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_58), .A2(n_148), .B1(n_407), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_59), .A2(n_203), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_60), .A2(n_263), .B1(n_638), .B2(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_61), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_62), .A2(n_328), .B1(n_464), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_63), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_64), .A2(n_184), .B1(n_793), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_65), .A2(n_229), .B1(n_470), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_66), .A2(n_248), .B1(n_402), .B2(n_724), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_68), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_69), .A2(n_224), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_71), .A2(n_92), .B1(n_573), .B2(n_574), .C(n_576), .Y(n_572) );
AO22x2_ASAP7_75t_L g368 ( .A1(n_72), .A2(n_231), .B1(n_359), .B2(n_360), .Y(n_368) );
INVx1_ASAP7_75t_L g976 ( .A(n_72), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_73), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_74), .A2(n_88), .B1(n_498), .B2(n_574), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_75), .A2(n_133), .B1(n_397), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_77), .A2(n_194), .B1(n_397), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_79), .A2(n_251), .B1(n_411), .B2(n_671), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_80), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_82), .A2(n_242), .B1(n_398), .B2(n_503), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_83), .A2(n_171), .B1(n_384), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_84), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_86), .A2(n_98), .B1(n_163), .B2(n_451), .C1(n_456), .C2(n_466), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_87), .A2(n_326), .B1(n_455), .B2(n_853), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_89), .Y(n_721) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_90), .A2(n_336), .B(n_344), .C(n_981), .Y(n_335) );
INVx1_ASAP7_75t_L g587 ( .A(n_93), .Y(n_587) );
XOR2x2_ASAP7_75t_L g824 ( .A(n_95), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g614 ( .A(n_97), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_99), .A2(n_247), .B1(n_469), .B2(n_762), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_100), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_101), .A2(n_239), .B1(n_432), .B2(n_437), .Y(n_598) );
INVx1_ASAP7_75t_L g980 ( .A(n_102), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_105), .A2(n_234), .B1(n_605), .B2(n_687), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_106), .A2(n_268), .B1(n_427), .B2(n_605), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_107), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_108), .Y(n_704) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_109), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_110), .B(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_111), .A2(n_245), .B1(n_438), .B2(n_767), .Y(n_766) );
AO22x1_ASAP7_75t_L g802 ( .A1(n_114), .A2(n_803), .B1(n_804), .B2(n_822), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_114), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_115), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_116), .A2(n_135), .B1(n_422), .B2(n_787), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_117), .B(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_119), .A2(n_306), .B1(n_411), .B2(n_428), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_120), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_122), .A2(n_126), .B1(n_469), .B2(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_123), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_124), .A2(n_565), .B1(n_591), .B2(n_592), .Y(n_564) );
INVx1_ASAP7_75t_L g591 ( .A(n_124), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g885 ( .A1(n_125), .A2(n_886), .B1(n_887), .B2(n_910), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_125), .Y(n_910) );
INVx1_ASAP7_75t_L g577 ( .A(n_127), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_129), .A2(n_303), .B1(n_473), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_130), .A2(n_202), .B1(n_479), .B2(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_131), .A2(n_146), .B1(n_683), .B2(n_908), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_132), .A2(n_144), .B1(n_602), .B2(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_134), .A2(n_314), .B1(n_736), .B2(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_136), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_138), .A2(n_270), .B1(n_498), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_139), .A2(n_221), .B1(n_473), .B2(n_764), .Y(n_763) );
AND2x6_ASAP7_75t_L g338 ( .A(n_141), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_141), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_142), .A2(n_254), .B1(n_490), .B2(n_544), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_143), .A2(n_293), .B1(n_455), .B2(n_458), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_145), .A2(n_235), .B1(n_371), .B2(n_379), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_149), .A2(n_284), .B1(n_544), .B2(n_546), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_150), .A2(n_213), .B1(n_230), .B2(n_356), .C1(n_379), .C2(n_455), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_151), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_153), .A2(n_274), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_154), .A2(n_300), .B1(n_435), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g673 ( .A(n_155), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_156), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_157), .A2(n_316), .B1(n_634), .B2(n_787), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_158), .A2(n_278), .B1(n_438), .B2(n_487), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_159), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_161), .A2(n_226), .B1(n_416), .B2(n_421), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_162), .A2(n_219), .B1(n_501), .B2(n_544), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_164), .A2(n_304), .B1(n_762), .B2(n_785), .Y(n_962) );
AO22x2_ASAP7_75t_L g366 ( .A1(n_165), .A2(n_220), .B1(n_359), .B2(n_363), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_165), .B(n_978), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_166), .A2(n_983), .B1(n_984), .B2(n_996), .Y(n_982) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_166), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_167), .A2(n_192), .B1(n_490), .B2(n_684), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_168), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_169), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_172), .A2(n_324), .B1(n_500), .B2(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g369 ( .A(n_173), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_175), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g821 ( .A1(n_179), .A2(n_292), .B1(n_299), .B2(n_451), .C1(n_503), .C2(n_504), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_180), .B(n_524), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_181), .A2(n_223), .B1(n_497), .B2(n_498), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_182), .Y(n_892) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_183), .B(n_849), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_185), .A2(n_272), .B1(n_384), .B2(n_609), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g1003 ( .A(n_187), .Y(n_1003) );
INVx1_ASAP7_75t_L g666 ( .A(n_189), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_190), .A2(n_269), .B1(n_609), .B2(n_628), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_191), .B(n_609), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_193), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_195), .A2(n_238), .B1(n_428), .B2(n_787), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_196), .B(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_197), .A2(n_260), .B1(n_470), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_198), .A2(n_217), .B1(n_401), .B2(n_524), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_200), .A2(n_253), .B1(n_412), .B2(n_634), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_201), .A2(n_261), .B1(n_464), .B2(n_466), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_204), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_206), .A2(n_323), .B1(n_422), .B2(n_432), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_207), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_208), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_209), .Y(n_917) );
INVx1_ASAP7_75t_L g661 ( .A(n_210), .Y(n_661) );
INVx1_ASAP7_75t_L g589 ( .A(n_211), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_212), .A2(n_295), .B1(n_455), .B2(n_853), .Y(n_852) );
AOI222xp33_ASAP7_75t_L g502 ( .A1(n_214), .A2(n_307), .B1(n_318), .B2(n_356), .C1(n_503), .C2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_215), .A2(n_332), .B1(n_493), .B2(n_585), .Y(n_725) );
INVx2_ASAP7_75t_L g343 ( .A(n_216), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_218), .A2(n_249), .B1(n_524), .B2(n_831), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_222), .B(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_225), .A2(n_745), .B1(n_746), .B2(n_769), .Y(n_744) );
CKINVDCx14_ASAP7_75t_R g769 ( .A(n_225), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_227), .A2(n_266), .B1(n_458), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_228), .A2(n_321), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g955 ( .A(n_236), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_237), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_241), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_243), .A2(n_331), .B1(n_479), .B2(n_481), .Y(n_478) );
XOR2x2_ASAP7_75t_L g349 ( .A(n_244), .B(n_350), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_246), .Y(n_525) );
INVx1_ASAP7_75t_L g359 ( .A(n_252), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_252), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_256), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_257), .Y(n_918) );
INVx1_ASAP7_75t_L g571 ( .A(n_258), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_259), .B(n_628), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_262), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_267), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_271), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_273), .B(n_584), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_276), .A2(n_330), .B1(n_386), .B2(n_462), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_277), .A2(n_308), .B1(n_552), .B2(n_554), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_279), .Y(n_542) );
INVx1_ASAP7_75t_L g342 ( .A(n_280), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_282), .Y(n_921) );
INVx1_ASAP7_75t_L g339 ( .A(n_283), .Y(n_339) );
INVx1_ASAP7_75t_L g617 ( .A(n_285), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_287), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_288), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_289), .A2(n_294), .B1(n_432), .B2(n_639), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_290), .Y(n_951) );
INVx1_ASAP7_75t_L g669 ( .A(n_291), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_297), .Y(n_927) );
INVx1_ASAP7_75t_L g568 ( .A(n_298), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_301), .A2(n_317), .B1(n_544), .B2(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_302), .Y(n_691) );
INVx1_ASAP7_75t_L g653 ( .A(n_309), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_310), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_311), .A2(n_327), .B1(n_497), .B2(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_312), .B(n_384), .Y(n_460) );
XOR2x2_ASAP7_75t_L g482 ( .A(n_313), .B(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_315), .A2(n_506), .B1(n_555), .B2(n_556), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_315), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_319), .B(n_656), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_320), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_322), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_325), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_329), .A2(n_914), .B1(n_937), .B2(n_938), .Y(n_913) );
INVx1_ASAP7_75t_L g937 ( .A(n_329), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_334), .Y(n_948) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_338), .B(n_340), .Y(n_337) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_339), .Y(n_972) );
OA21x2_ASAP7_75t_L g1001 ( .A1(n_340), .A2(n_971), .B(n_1002), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_741), .B1(n_966), .B2(n_967), .C(n_968), .Y(n_344) );
INVx1_ASAP7_75t_L g967 ( .A(n_345), .Y(n_967) );
XOR2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_560), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_441), .B1(n_558), .B2(n_559), .Y(n_346) );
INVx1_ASAP7_75t_L g558 ( .A(n_347), .Y(n_558) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND3x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_405), .C(n_425), .Y(n_350) );
NOR2x1_ASAP7_75t_SL g351 ( .A(n_352), .B(n_382), .Y(n_351) );
OAI21xp5_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_369), .B(n_370), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g893 ( .A1(n_353), .A2(n_894), .B1(n_895), .B2(n_896), .C(n_897), .Y(n_893) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g613 ( .A(n_355), .Y(n_613) );
INVx4_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_356), .Y(n_451) );
INVx2_ASAP7_75t_L g622 ( .A(n_356), .Y(n_622) );
BUFx3_ASAP7_75t_L g775 ( .A(n_356), .Y(n_775) );
INVx2_ASAP7_75t_SL g828 ( .A(n_356), .Y(n_828) );
AND2x6_ASAP7_75t_L g356 ( .A(n_357), .B(n_364), .Y(n_356) );
AND2x4_ASAP7_75t_L g402 ( .A(n_357), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g536 ( .A(n_357), .Y(n_536) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_362), .Y(n_357) );
AND2x2_ASAP7_75t_L g378 ( .A(n_358), .B(n_366), .Y(n_378) );
INVx2_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_361), .Y(n_363) );
INVx2_ASAP7_75t_L g377 ( .A(n_362), .Y(n_377) );
AND2x2_ASAP7_75t_L g387 ( .A(n_362), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g395 ( .A(n_362), .B(n_388), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
AND2x6_ASAP7_75t_L g411 ( .A(n_364), .B(n_394), .Y(n_411) );
AND2x2_ASAP7_75t_L g429 ( .A(n_364), .B(n_414), .Y(n_429) );
AND2x4_ASAP7_75t_L g437 ( .A(n_364), .B(n_387), .Y(n_437) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
AND2x2_ASAP7_75t_L g389 ( .A(n_365), .B(n_368), .Y(n_389) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g420 ( .A(n_366), .B(n_404), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_366), .B(n_368), .Y(n_424) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g376 ( .A(n_368), .Y(n_376) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g718 ( .A(n_373), .Y(n_718) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_374), .Y(n_455) );
BUFx4f_ASAP7_75t_SL g503 ( .A(n_374), .Y(n_503) );
BUFx2_ASAP7_75t_L g616 ( .A(n_374), .Y(n_616) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_374), .Y(n_839) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_376), .Y(n_381) );
AND2x2_ASAP7_75t_L g414 ( .A(n_377), .B(n_388), .Y(n_414) );
INVx1_ASAP7_75t_L g531 ( .A(n_377), .Y(n_531) );
AND2x4_ASAP7_75t_L g380 ( .A(n_378), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g398 ( .A(n_378), .B(n_399), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_378), .B(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx12f_ASAP7_75t_L g458 ( .A(n_380), .Y(n_458) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_380), .Y(n_524) );
INVx1_ASAP7_75t_L g720 ( .A(n_380), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .C(n_396), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g585 ( .A(n_385), .Y(n_585) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
BUFx4f_ASAP7_75t_L g628 ( .A(n_386), .Y(n_628) );
BUFx2_ASAP7_75t_L g819 ( .A(n_386), .Y(n_819) );
BUFx2_ASAP7_75t_L g837 ( .A(n_386), .Y(n_837) );
AND2x6_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
AND2x2_ASAP7_75t_L g419 ( .A(n_387), .B(n_420), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_387), .B(n_389), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_387), .B(n_420), .Y(n_570) );
AND2x4_ASAP7_75t_L g393 ( .A(n_389), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g413 ( .A(n_389), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g512 ( .A(n_389), .Y(n_512) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx5_ASAP7_75t_L g462 ( .A(n_392), .Y(n_462) );
INVx2_ASAP7_75t_L g584 ( .A(n_392), .Y(n_584) );
INVx2_ASAP7_75t_L g609 ( .A(n_392), .Y(n_609) );
INVx4_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g511 ( .A(n_395), .B(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g465 ( .A(n_398), .Y(n_465) );
BUFx2_ASAP7_75t_L g724 ( .A(n_398), .Y(n_724) );
BUFx3_ASAP7_75t_L g853 ( .A(n_398), .Y(n_853) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x6_ASAP7_75t_L g423 ( .A(n_400), .B(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_SL g466 ( .A(n_402), .Y(n_466) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_402), .Y(n_611) );
BUFx3_ASAP7_75t_L g658 ( .A(n_402), .Y(n_658) );
INVx1_ASAP7_75t_L g537 ( .A(n_403), .Y(n_537) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_415), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g500 ( .A(n_410), .Y(n_500) );
INVx4_ASAP7_75t_L g573 ( .A(n_410), .Y(n_573) );
INVx2_ASAP7_75t_L g605 ( .A(n_410), .Y(n_605) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_410), .Y(n_814) );
INVx11_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx11_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
INVx4_ASAP7_75t_L g488 ( .A(n_412), .Y(n_488) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g471 ( .A(n_413), .Y(n_471) );
BUFx3_ASAP7_75t_L g684 ( .A(n_413), .Y(n_684) );
BUFx3_ASAP7_75t_L g762 ( .A(n_413), .Y(n_762) );
BUFx3_ASAP7_75t_L g793 ( .A(n_413), .Y(n_793) );
AND2x2_ASAP7_75t_L g433 ( .A(n_414), .B(n_420), .Y(n_433) );
AND2x4_ASAP7_75t_L g439 ( .A(n_414), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_414), .B(n_420), .Y(n_580) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g545 ( .A(n_418), .Y(n_545) );
INVx4_ASAP7_75t_L g601 ( .A(n_418), .Y(n_601) );
INVx2_ASAP7_75t_L g787 ( .A(n_418), .Y(n_787) );
INVx3_ASAP7_75t_L g816 ( .A(n_418), .Y(n_816) );
INVx8_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
BUFx2_ASAP7_75t_L g602 ( .A(n_422), .Y(n_602) );
BUFx2_ASAP7_75t_L g764 ( .A(n_422), .Y(n_764) );
INVx6_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g546 ( .A(n_423), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_423), .A2(n_568), .B1(n_569), .B2(n_571), .Y(n_567) );
INVx1_ASAP7_75t_SL g731 ( .A(n_423), .Y(n_731) );
INVx1_ASAP7_75t_L g440 ( .A(n_424), .Y(n_440) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_434), .Y(n_425) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g680 ( .A(n_428), .Y(n_680) );
BUFx3_ASAP7_75t_L g807 ( .A(n_428), .Y(n_807) );
BUFx3_ASAP7_75t_L g908 ( .A(n_428), .Y(n_908) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_SL g469 ( .A(n_429), .Y(n_469) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_429), .Y(n_486) );
INVx2_ASAP7_75t_L g792 ( .A(n_429), .Y(n_792) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g476 ( .A(n_433), .Y(n_476) );
BUFx3_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
BUFx3_ASAP7_75t_L g868 ( .A(n_433), .Y(n_868) );
INVx2_ASAP7_75t_L g689 ( .A(n_435), .Y(n_689) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
INVx3_ASAP7_75t_L g671 ( .A(n_436), .Y(n_671) );
INVx2_ASAP7_75t_L g933 ( .A(n_436), .Y(n_933) );
INVx6_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
BUFx3_ASAP7_75t_L g550 ( .A(n_437), .Y(n_550) );
BUFx3_ASAP7_75t_L g638 ( .A(n_437), .Y(n_638) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_SL g477 ( .A(n_439), .Y(n_477) );
BUFx3_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
BUFx3_ASAP7_75t_L g554 ( .A(n_439), .Y(n_554) );
BUFx3_ASAP7_75t_L g639 ( .A(n_439), .Y(n_639) );
BUFx3_ASAP7_75t_L g736 ( .A(n_439), .Y(n_736) );
BUFx2_ASAP7_75t_L g785 ( .A(n_439), .Y(n_785) );
INVx1_ASAP7_75t_L g858 ( .A(n_439), .Y(n_858) );
AND2x2_ASAP7_75t_L g634 ( .A(n_440), .B(n_531), .Y(n_634) );
INVx1_ASAP7_75t_L g559 ( .A(n_441), .Y(n_559) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_505), .B2(n_557), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_482), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_467), .C(n_474), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_459), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_452), .B(n_453), .Y(n_449) );
OAI222xp33_ASAP7_75t_L g716 ( .A1(n_450), .A2(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_721), .Y(n_716) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
INVx2_ASAP7_75t_SL g895 ( .A(n_454), .Y(n_895) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_458), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .C(n_463), .Y(n_459) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_462), .Y(n_493) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_462), .Y(n_835) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g553 ( .A(n_476), .Y(n_553) );
BUFx4f_ASAP7_75t_SL g767 ( .A(n_476), .Y(n_767) );
INVx1_ASAP7_75t_SL g582 ( .A(n_477), .Y(n_582) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
INVx3_ASAP7_75t_L g668 ( .A(n_480), .Y(n_668) );
INVx3_ASAP7_75t_L g575 ( .A(n_481), .Y(n_575) );
NAND4xp75_ASAP7_75t_L g483 ( .A(n_484), .B(n_491), .C(n_495), .D(n_502), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
INVx1_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI221xp5_ASAP7_75t_SL g539 ( .A1(n_488), .A2(n_540), .B1(n_541), .B2(n_542), .C(n_543), .Y(n_539) );
INVx3_ASAP7_75t_L g650 ( .A(n_488), .Y(n_650) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_492), .B(n_494), .Y(n_491) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
BUFx2_ASAP7_75t_L g734 ( .A(n_497), .Y(n_734) );
INVx1_ASAP7_75t_L g809 ( .A(n_497), .Y(n_809) );
INVxp67_ASAP7_75t_L g663 ( .A(n_498), .Y(n_663) );
INVx1_ASAP7_75t_L g519 ( .A(n_503), .Y(n_519) );
INVx1_ASAP7_75t_L g702 ( .A(n_503), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_504), .Y(n_705) );
INVx1_ASAP7_75t_L g557 ( .A(n_505), .Y(n_557) );
INVx1_ASAP7_75t_L g556 ( .A(n_506), .Y(n_556) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_538), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .C(n_526), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_513), .B2(n_514), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_510), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g697 ( .A(n_511), .Y(n_697) );
BUFx3_ASAP7_75t_L g947 ( .A(n_511), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_514), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g654 ( .A(n_516), .Y(n_654) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g700 ( .A(n_517), .Y(n_700) );
OAI222xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B1(n_521), .B2(n_522), .C1(n_523), .C2(n_525), .Y(n_518) );
OAI222xp33_ASAP7_75t_L g701 ( .A1(n_521), .A2(n_702), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_532), .B2(n_533), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_528), .A2(n_533), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_SL g926 ( .A(n_529), .Y(n_926) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_530), .Y(n_757) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g901 ( .A(n_534), .Y(n_901) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_535), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_535), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
BUFx2_ASAP7_75t_L g928 ( .A(n_535), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_535), .A2(n_588), .B1(n_954), .B2(n_955), .Y(n_953) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_674), .B1(n_675), .B2(n_740), .Y(n_560) );
INVx1_ASAP7_75t_L g740 ( .A(n_561), .Y(n_740) );
OAI22xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_563), .B1(n_644), .B2(n_645), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OA22x2_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_593), .B1(n_594), .B2(n_643), .Y(n_563) );
INVx1_ASAP7_75t_L g643 ( .A(n_564), .Y(n_643) );
INVx1_ASAP7_75t_L g592 ( .A(n_565), .Y(n_592) );
AND4x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_572), .C(n_583), .D(n_590), .Y(n_565) );
BUFx2_ASAP7_75t_R g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_581), .B2(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g662 ( .A(n_579), .Y(n_662) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g656 ( .A(n_584), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_588), .A2(n_899), .B1(n_900), .B2(n_901), .Y(n_898) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_618), .B1(n_641), .B2(n_642), .Y(n_594) );
INVx2_ASAP7_75t_SL g641 ( .A(n_595), .Y(n_641) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_617), .Y(n_595) );
NOR4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .C(n_607), .D(n_612), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_599), .Y(n_597) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g832 ( .A(n_611), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_614), .B(n_615), .Y(n_612) );
OAI21xp5_ASAP7_75t_SL g752 ( .A1(n_613), .A2(n_753), .B(n_754), .Y(n_752) );
OAI221xp5_ASAP7_75t_SL g920 ( .A1(n_613), .A2(n_702), .B1(n_921), .B2(n_922), .C(n_923), .Y(n_920) );
INVx1_ASAP7_75t_L g642 ( .A(n_618), .Y(n_642) );
OA22x2_ASAP7_75t_SL g712 ( .A1(n_618), .A2(n_642), .B1(n_713), .B2(n_737), .Y(n_712) );
XOR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_640), .Y(n_618) );
NAND2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_630), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B(n_624), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .C(n_629), .Y(n_625) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_639), .Y(n_687) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_673), .Y(n_646) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .C(n_659), .D(n_672), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
OA211x2_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_655), .C(n_657), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_654), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
OA211x2_ASAP7_75t_L g870 ( .A1(n_654), .A2(n_871), .B(n_872), .C(n_873), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_665), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_660) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_662), .A2(n_689), .B1(n_690), .B2(n_691), .C(n_692), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_712), .B1(n_738), .B2(n_739), .Y(n_675) );
INVx1_ASAP7_75t_L g738 ( .A(n_676), .Y(n_738) );
INVx1_ASAP7_75t_L g711 ( .A(n_677), .Y(n_711) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_678), .B(n_693), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_688), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_679) );
INVx2_ASAP7_75t_L g729 ( .A(n_680), .Y(n_729) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_701), .C(n_707), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_699), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g750 ( .A(n_697), .Y(n_750) );
INVx1_ASAP7_75t_SL g891 ( .A(n_697), .Y(n_891) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g919 ( .A(n_700), .Y(n_919) );
INVx1_ASAP7_75t_L g949 ( .A(n_700), .Y(n_949) );
INVx2_ASAP7_75t_L g739 ( .A(n_712), .Y(n_739) );
INVx1_ASAP7_75t_L g737 ( .A(n_713), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_726), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_722), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_732), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g966 ( .A(n_741), .Y(n_966) );
AOI22xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_880), .B1(n_881), .B2(n_965), .Y(n_741) );
INVx1_ASAP7_75t_L g965 ( .A(n_742), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_797), .B1(n_798), .B2(n_879), .Y(n_742) );
INVx2_ASAP7_75t_SL g879 ( .A(n_743), .Y(n_879) );
AO22x1_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_770), .B1(n_795), .B2(n_796), .Y(n_743) );
INVx1_ASAP7_75t_L g796 ( .A(n_744), .Y(n_796) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_759), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .C(n_755), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_765), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx3_ASAP7_75t_SL g795 ( .A(n_770), .Y(n_795) );
AO22x1_ASAP7_75t_L g940 ( .A1(n_770), .A2(n_795), .B1(n_941), .B2(n_942), .Y(n_940) );
XOR2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_794), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_772), .B(n_782), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_778), .Y(n_772) );
OAI21xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_776), .B(n_777), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g950 ( .A1(n_774), .A2(n_951), .B(n_952), .Y(n_950) );
INVx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .C(n_781), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_788), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g844 ( .A(n_792), .Y(n_844) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI22x1_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_863), .B2(n_864), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
XNOR2x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_823), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
NAND4xp75_ASAP7_75t_SL g804 ( .A(n_805), .B(n_811), .C(n_817), .D(n_821), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_815), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_SL g817 ( .A(n_818), .B(n_820), .Y(n_817) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_848), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_826), .B(n_840), .Y(n_825) );
NOR2xp33_ASAP7_75t_SL g826 ( .A(n_827), .B(n_833), .Y(n_826) );
OAI21xp5_ASAP7_75t_SL g827 ( .A1(n_828), .A2(n_829), .B(n_830), .Y(n_827) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .C(n_838), .Y(n_833) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
NAND4xp75_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .C(n_859), .D(n_862), .Y(n_849) );
AND2x2_ASAP7_75t_SL g850 ( .A(n_851), .B(n_852), .Y(n_850) );
AND2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
INVx3_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
XOR2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_878), .Y(n_864) );
NAND4xp75_ASAP7_75t_L g865 ( .A(n_866), .B(n_870), .C(n_874), .D(n_877), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_869), .Y(n_866) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B1(n_911), .B2(n_964), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_SL g886 ( .A(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_902), .Y(n_887) );
NOR3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_893), .C(n_898), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g964 ( .A(n_911), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B1(n_939), .B2(n_940), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g938 ( .A(n_914), .Y(n_938) );
AND2x2_ASAP7_75t_SL g914 ( .A(n_915), .B(n_929), .Y(n_914) );
NOR3xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_920), .C(n_924), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_930), .B(n_934), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx2_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
XOR2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_963), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_956), .Y(n_943) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_950), .C(n_953), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_948), .B2(n_949), .Y(n_945) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_960), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
INVx1_ASAP7_75t_SL g968 ( .A(n_969), .Y(n_968) );
NOR2x1_ASAP7_75t_L g969 ( .A(n_970), .B(n_974), .Y(n_969) );
OR2x2_ASAP7_75t_SL g1007 ( .A(n_970), .B(n_975), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_972), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_972), .B(n_1000), .Y(n_1002) );
CKINVDCx16_ASAP7_75t_R g1000 ( .A(n_973), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_975), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_977), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_979), .B(n_980), .Y(n_978) );
OAI322xp33_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_997), .A3(n_998), .B1(n_1001), .B2(n_1003), .C1(n_1004), .C2(n_1005), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_984), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
XOR2x2_ASAP7_75t_L g1004 ( .A(n_985), .B(n_1003), .Y(n_1004) );
NAND4xp75_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .C(n_992), .D(n_995), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
AND2x2_ASAP7_75t_SL g989 ( .A(n_990), .B(n_991), .Y(n_989) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_1006), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_1007), .Y(n_1006) );
endmodule