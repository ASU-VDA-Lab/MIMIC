module fake_jpeg_18328_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_22),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_27),
.B2(n_19),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_18),
.B1(n_19),
.B2(n_13),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_43),
.B1(n_36),
.B2(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

OA21x2_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_21),
.B(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_16),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_21),
.B1(n_29),
.B2(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_32),
.B1(n_39),
.B2(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_41),
.B1(n_49),
.B2(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_63),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_42),
.B(n_43),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_42),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_70),
.B1(n_60),
.B2(n_59),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_9),
.C(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_9),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_55),
.C(n_58),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_77),
.C(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_34),
.C(n_17),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_17),
.C(n_10),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_62),
.C(n_10),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_87),
.C(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_75),
.B1(n_79),
.B2(n_0),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_13),
.B1(n_6),
.B2(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_15),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_5),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_95),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_5),
.B(n_2),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_7),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_83),
.B1(n_82),
.B2(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_99),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_12),
.C(n_11),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.C(n_92),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_12),
.C(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_4),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_97),
.B(n_3),
.C(n_4),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_104),
.B(n_0),
.Y(n_106)
);

NAND4xp25_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_4),
.C(n_7),
.D(n_11),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.C(n_1),
.Y(n_109)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_108),
.Y(n_111)
);


endmodule