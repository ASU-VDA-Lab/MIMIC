module fake_netlist_1_420_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g11 ( .A(n_4), .B(n_1), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_7), .B(n_3), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_0), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_10), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_10), .B(n_1), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_19), .B(n_13), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_16), .B(n_13), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_16), .B1(n_15), .B2(n_18), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_17), .B1(n_12), .B2(n_11), .C(n_13), .Y(n_24) );
OR2x6_ASAP7_75t_L g25 ( .A(n_23), .B(n_22), .Y(n_25) );
INVxp67_ASAP7_75t_SL g26 ( .A(n_24), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_25), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B1(n_21), .B2(n_5), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_27), .B(n_25), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
CKINVDCx20_ASAP7_75t_R g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
AOI322xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_3), .A3(n_7), .B1(n_8), .B2(n_9), .C1(n_31), .C2(n_13), .Y(n_34) );
endmodule