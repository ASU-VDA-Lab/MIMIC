module real_jpeg_23581_n_26 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_24, n_6, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_158, n_149, n_16, n_15, n_13, n_155, n_26);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_24;
input n_6;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_158;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_26;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_3),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_3),
.B(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.C(n_124),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_5),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_7),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_9),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_129),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_11),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_12),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_13),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_15),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_16),
.B(n_78),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_18),
.B(n_47),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_19),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_20),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_40),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_25),
.B(n_96),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_142),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_139),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_32),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_33),
.Y(n_127)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_36),
.B(n_135),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_138),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_132),
.B(n_137),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_128),
.B(n_131),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_123),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_118),
.B(n_122),
.Y(n_49)
);

OAI321xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_108),
.A3(n_113),
.B1(n_116),
.B2(n_117),
.C(n_148),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_100),
.B(n_107),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_95),
.B(n_99),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_89),
.B(n_94),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_88),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_81),
.B(n_87),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_77),
.B(n_80),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_70),
.B(n_76),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_145),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_136),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_149),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_150),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_151),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_152),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_153),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_154),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_155),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_156),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_157),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_158),
.Y(n_115)
);


endmodule