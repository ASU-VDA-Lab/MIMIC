module fake_jpeg_4780_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_15),
.B(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_46),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_52),
.B1(n_55),
.B2(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_24),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_25),
.B1(n_30),
.B2(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_30),
.B1(n_15),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_62),
.B1(n_19),
.B2(n_21),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_33),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_69),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_20),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_38),
.B(n_33),
.C(n_35),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_94)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_49),
.B1(n_54),
.B2(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_115)
);

NOR2x1p5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_49),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_76),
.B(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_54),
.C(n_49),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_58),
.B1(n_64),
.B2(n_57),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_83),
.B1(n_77),
.B2(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_58),
.B1(n_57),
.B2(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_60),
.B1(n_41),
.B2(n_27),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_66),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_110),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_81),
.B(n_73),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_113),
.B(n_124),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_36),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_70),
.B(n_35),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_120),
.C(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_119),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_71),
.B1(n_66),
.B2(n_19),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_127),
.B1(n_107),
.B2(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_23),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_48),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_0),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_84),
.B(n_36),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_48),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_84),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_139),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_106),
.B(n_99),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_141),
.B(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_146),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_92),
.B(n_87),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_100),
.B1(n_105),
.B2(n_101),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_129),
.B1(n_115),
.B2(n_130),
.Y(n_155)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_101),
.B1(n_36),
.B2(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_68),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_114),
.C(n_120),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_162),
.C(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_122),
.C(n_109),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_112),
.C(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_65),
.C(n_29),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_165),
.C(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_29),
.C(n_22),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_29),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_29),
.B(n_22),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_147),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_151),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_172),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_131),
.Y(n_172)
);

BUFx12f_ASAP7_75t_SL g175 ( 
.A(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_165),
.B(n_158),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_131),
.C(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_181),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_1),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_139),
.C(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_143),
.B1(n_135),
.B2(n_138),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_22),
.B1(n_29),
.B2(n_3),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_134),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_176),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_153),
.B(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_191),
.B1(n_195),
.B2(n_181),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_154),
.C(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_194),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_157),
.B(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_192),
.Y(n_198)
);

AOI321xp33_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_149),
.A3(n_159),
.B1(n_135),
.B2(n_146),
.C(n_29),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_177),
.C(n_176),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_203),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_204),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_182),
.B1(n_174),
.B2(n_186),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_186),
.B1(n_2),
.B2(n_3),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_1),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_203),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_216),
.B(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_198),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_208),
.C(n_198),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_220),
.B(n_221),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_10),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_2),
.C(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_214),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_224),
.A3(n_4),
.B1(n_7),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

OAI311xp33_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.C1(n_204),
.Y(n_226)
);


endmodule