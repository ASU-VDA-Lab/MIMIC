module fake_jpeg_6101_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_26),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_55),
.B1(n_29),
.B2(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_59),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_15),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_21),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_70),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_61),
.B(n_40),
.C(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_41),
.B1(n_15),
.B2(n_29),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_15),
.B1(n_29),
.B2(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_81),
.B1(n_45),
.B2(n_61),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_78),
.B(n_60),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_52),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_89),
.B1(n_27),
.B2(n_17),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_21),
.B1(n_17),
.B2(n_28),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_93),
.B1(n_100),
.B2(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_50),
.C(n_57),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_105),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_107),
.C(n_110),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_49),
.B1(n_43),
.B2(n_46),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_51),
.B1(n_61),
.B2(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_52),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_64),
.C(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_86),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_48),
.B(n_27),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_51),
.B(n_63),
.C(n_16),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_77),
.B1(n_66),
.B2(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_62),
.B1(n_63),
.B2(n_16),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_73),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_125),
.B1(n_99),
.B2(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_123),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_75),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_82),
.B1(n_83),
.B2(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_132),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_130),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_111),
.B1(n_93),
.B2(n_90),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_R g129 ( 
.A(n_110),
.B(n_32),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_137),
.B(n_123),
.Y(n_144)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_85),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_139),
.Y(n_165)
);

NOR2x1_ASAP7_75t_R g137 ( 
.A(n_110),
.B(n_32),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_99),
.B(n_90),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_56),
.C(n_31),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_107),
.B1(n_62),
.B2(n_69),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_118),
.B1(n_121),
.B2(n_119),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_149),
.B(n_166),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_106),
.B1(n_100),
.B2(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_69),
.B1(n_84),
.B2(n_70),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_105),
.C(n_98),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_105),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_161),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_92),
.C(n_103),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_108),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_20),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_128),
.B1(n_134),
.B2(n_130),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_115),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_107),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_160),
.B(n_167),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_107),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_56),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_138),
.C(n_118),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_56),
.C(n_20),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_155),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_113),
.B(n_111),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_151),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_135),
.C(n_122),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_185),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_116),
.B1(n_133),
.B2(n_134),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_167),
.B1(n_160),
.B2(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_187),
.C(n_194),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_186),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_70),
.B1(n_63),
.B2(n_73),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_150),
.B1(n_155),
.B2(n_163),
.Y(n_199)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_23),
.B1(n_16),
.B2(n_127),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_149),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_20),
.B(n_23),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_1),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_56),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_146),
.C(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_204),
.C(n_213),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_179),
.B1(n_209),
.B2(n_191),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_210),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_154),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_209),
.B1(n_172),
.B2(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_144),
.B1(n_164),
.B2(n_150),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_156),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_174),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_127),
.B(n_23),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_181),
.B1(n_180),
.B2(n_171),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_16),
.C(n_23),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_232),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_187),
.C(n_192),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_229),
.C(n_235),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_184),
.C(n_182),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_240),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_182),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_217),
.B(n_218),
.C(n_3),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_183),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_183),
.C(n_173),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_210),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_12),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_1),
.C(n_2),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_214),
.C(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_202),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_251),
.C(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_195),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_207),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_206),
.B(n_229),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_220),
.B1(n_237),
.B2(n_222),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_198),
.C(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_210),
.C(n_201),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_1),
.C(n_2),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_224),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_217),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_12),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_269),
.B(n_270),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_243),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_273),
.Y(n_283)
);

XOR2x1_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_3),
.C(n_4),
.Y(n_275)
);

BUFx4f_ASAP7_75t_SL g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

AOI321xp33_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_264),
.A3(n_273),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_251),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_285),
.B(n_10),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_286),
.C(n_4),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_242),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_243),
.B1(n_242),
.B2(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_11),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_4),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_290),
.B(n_292),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_267),
.B(n_265),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_293),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_3),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_6),
.C(n_7),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_281),
.C(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_8),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_8),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_303),
.B(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_287),
.B1(n_278),
.B2(n_283),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_280),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

NAND2x1_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_10),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_312),
.B(n_309),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.C(n_304),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_10),
.Y(n_317)
);


endmodule