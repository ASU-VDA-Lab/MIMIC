module fake_jpeg_16709_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_37),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_56),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_52),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_52),
.B1(n_43),
.B2(n_47),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_1),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_79),
.Y(n_96)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_2),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_85),
.B(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_3),
.B(n_4),
.C(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_99),
.Y(n_100)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_10),
.C(n_11),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_15),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_81),
.B1(n_86),
.B2(n_76),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_106),
.C(n_100),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_114),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

OAI322xp33_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_103),
.A3(n_110),
.B1(n_20),
.B2(n_21),
.C1(n_22),
.C2(n_23),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_92),
.B1(n_90),
.B2(n_24),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_119),
.C(n_90),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_17),
.CI(n_19),
.CON(n_124),
.SN(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_26),
.Y(n_125)
);

OAI21x1_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_30),
.B(n_31),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_32),
.B(n_35),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_36),
.Y(n_128)
);


endmodule