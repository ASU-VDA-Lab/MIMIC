module fake_jpeg_23275_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_1),
.C(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_47),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_19),
.B1(n_28),
.B2(n_20),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_51),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_34),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_28),
.B1(n_22),
.B2(n_26),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_16),
.B1(n_20),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_34),
.B1(n_33),
.B2(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_59),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_62),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_37),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_52),
.C(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_34),
.B1(n_38),
.B2(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_35),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_79),
.B1(n_85),
.B2(n_22),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_78),
.B1(n_17),
.B2(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_51),
.B1(n_38),
.B2(n_33),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_52),
.B1(n_49),
.B2(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_109),
.B1(n_75),
.B2(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_95),
.Y(n_116)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_108),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_70),
.B(n_77),
.C(n_80),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_69),
.B1(n_63),
.B2(n_81),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_11),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_17),
.B1(n_32),
.B2(n_54),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_65),
.B1(n_79),
.B2(n_62),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_29),
.A3(n_25),
.B1(n_48),
.B2(n_18),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_71),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_120),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_60),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_118),
.B(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_123),
.Y(n_151)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_136),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_134),
.B(n_84),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_81),
.B(n_72),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_61),
.B(n_70),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_61),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_73),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_89),
.B(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_85),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_146),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_104),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_25),
.B(n_29),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_104),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_153),
.C(n_155),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_73),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_127),
.B1(n_114),
.B2(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_161),
.B1(n_132),
.B2(n_130),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_87),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_105),
.B1(n_18),
.B2(n_21),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_87),
.C(n_110),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_160),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_101),
.C(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_118),
.C(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_88),
.C(n_86),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_169),
.B1(n_185),
.B2(n_150),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_120),
.B1(n_115),
.B2(n_69),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_184),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_88),
.C(n_30),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_69),
.B1(n_83),
.B2(n_100),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_174),
.B1(n_178),
.B2(n_161),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_142),
.B1(n_158),
.B2(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_105),
.B1(n_30),
.B2(n_21),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_179),
.A2(n_186),
.B(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_48),
.B1(n_54),
.B2(n_29),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_167),
.B(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_194),
.B(n_195),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_155),
.C(n_145),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_202),
.C(n_181),
.Y(n_212)
);

OAI322xp33_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_162),
.A3(n_148),
.B1(n_141),
.B2(n_153),
.C1(n_159),
.C2(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_198),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_148),
.B(n_146),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_141),
.B(n_156),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_185),
.B1(n_169),
.B2(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_147),
.B1(n_48),
.B2(n_25),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_1),
.C(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_204),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_172),
.C(n_180),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_170),
.B1(n_179),
.B2(n_183),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_197),
.B1(n_196),
.B2(n_199),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_202),
.CI(n_193),
.CON(n_216),
.SN(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_189),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_218),
.A2(n_188),
.B(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_227),
.B1(n_221),
.B2(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_211),
.A2(n_200),
.B1(n_188),
.B2(n_189),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_228),
.B1(n_216),
.B2(n_3),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_200),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_6),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_207),
.B(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_218),
.B1(n_210),
.B2(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_214),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_235),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_232),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_212),
.C(n_213),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_6),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_238),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_243),
.B(n_244),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_224),
.B(n_9),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_11),
.B(n_12),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_224),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_231),
.B(n_235),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_237),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_11),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_245),
.C(n_14),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_253),
.B(n_13),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_13),
.C(n_14),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_13),
.B(n_14),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.C(n_15),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_15),
.Y(n_257)
);


endmodule