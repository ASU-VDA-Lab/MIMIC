module fake_jpeg_18595_n_166 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_21),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_9),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_0),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_65),
.B1(n_49),
.B2(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_93),
.B1(n_75),
.B2(n_67),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_49),
.B1(n_65),
.B2(n_76),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_76),
.B1(n_73),
.B2(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_52),
.B1(n_51),
.B2(n_62),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_57),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_73),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_55),
.B(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_107),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_77),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_90),
.B(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_115),
.B1(n_119),
.B2(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_89),
.B1(n_91),
.B2(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_113),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_89),
.B1(n_53),
.B2(n_61),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_70),
.B1(n_71),
.B2(n_5),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_70),
.A3(n_71),
.B1(n_27),
.B2(n_44),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_28),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_72),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_68),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_124),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_8),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_142),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_127),
.B1(n_138),
.B2(n_109),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.C(n_145),
.Y(n_153)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_154),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_148),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_144),
.B1(n_152),
.B2(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_140),
.B(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_138),
.B(n_10),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_34),
.B(n_12),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_35),
.C(n_13),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_36),
.A3(n_16),
.B1(n_18),
.B2(n_25),
.C1(n_26),
.C2(n_42),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_166)
);


endmodule