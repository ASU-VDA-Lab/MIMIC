module fake_jpeg_30656_n_217 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_12),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_43)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_1),
.Y(n_89)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_57),
.Y(n_66)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_11),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_21),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_76),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_36),
.B1(n_20),
.B2(n_37),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_78),
.B1(n_83),
.B2(n_45),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_25),
.B1(n_35),
.B2(n_19),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_40),
.B1(n_23),
.B2(n_42),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_23),
.B1(n_21),
.B2(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_48),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_23),
.B(n_5),
.C(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_88),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_41),
.C(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_108),
.Y(n_139)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_102),
.B1(n_93),
.B2(n_69),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_38),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_7),
.A3(n_39),
.B1(n_83),
.B2(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_70),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_64),
.A2(n_71),
.B(n_86),
.C(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_120),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_69),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_107),
.B1(n_108),
.B2(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_144),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_81),
.B(n_65),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_101),
.B(n_114),
.C(n_113),
.D(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_72),
.B1(n_74),
.B2(n_81),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_120),
.B1(n_106),
.B2(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_65),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_147),
.B1(n_149),
.B2(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_97),
.C(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_135),
.C(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_107),
.B1(n_103),
.B2(n_111),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_130),
.B1(n_128),
.B2(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_96),
.B1(n_119),
.B2(n_98),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_155),
.B(n_163),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_126),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_131),
.B(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_113),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_123),
.B1(n_133),
.B2(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_146),
.C(n_154),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_135),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_177),
.B1(n_149),
.B2(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_138),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_141),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_182),
.B1(n_189),
.B2(n_175),
.C(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_184),
.C(n_183),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_151),
.B(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_154),
.C(n_151),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_153),
.B(n_145),
.C(n_162),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_171),
.B1(n_164),
.B2(n_172),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_166),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_153),
.A3(n_123),
.B1(n_127),
.B2(n_148),
.C1(n_150),
.C2(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_170),
.B1(n_174),
.B2(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_183),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_178),
.B1(n_173),
.B2(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_185),
.B(n_186),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_184),
.C(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_202),
.B(n_199),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_195),
.B(n_186),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_194),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_200),
.C(n_202),
.Y(n_210)
);

AOI31xp33_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_186),
.A3(n_198),
.B(n_133),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_142),
.B1(n_129),
.B2(n_122),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_205),
.B(n_125),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_206),
.B1(n_134),
.B2(n_125),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_212),
.C(n_214),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_85),
.Y(n_217)
);


endmodule