module fake_jpeg_2710_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_36),
.B(n_39),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_40),
.B1(n_46),
.B2(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_74),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_47),
.C(n_37),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_82),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_64),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_35),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_55),
.B1(n_54),
.B2(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_61),
.B1(n_64),
.B2(n_35),
.Y(n_86)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_70),
.B(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_1),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_96),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_84),
.C(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_2),
.B(n_5),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_102),
.B(n_86),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_6),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_89),
.C(n_83),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_109),
.C(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_93),
.B1(n_98),
.B2(n_23),
.Y(n_114)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_21),
.C(n_30),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_20),
.C(n_29),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_116)
);

OAI321xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_31),
.A3(n_12),
.B1(n_17),
.B2(n_18),
.C(n_11),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_108),
.C(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_122),
.B(n_123),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_110),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_115),
.CI(n_116),
.CON(n_124),
.SN(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_121),
.B(n_107),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_24),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_28),
.C(n_25),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_26),
.Y(n_131)
);


endmodule