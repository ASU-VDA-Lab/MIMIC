module fake_jpeg_30203_n_72 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx11_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_38),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_1),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_6),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_15),
.B(n_25),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_11),
.C(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_31),
.B1(n_30),
.B2(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_12),
.B1(n_22),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_10),
.B1(n_20),
.B2(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_53),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_41),
.C(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.C(n_62),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.C(n_60),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_62),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_54),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_65),
.Y(n_70)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_3),
.B(n_4),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_4),
.B(n_5),
.Y(n_72)
);


endmodule