module fake_jpeg_16086_n_166 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_38),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_30),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_25),
.B1(n_23),
.B2(n_16),
.Y(n_70)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_29),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_25),
.B1(n_37),
.B2(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_73),
.B1(n_74),
.B2(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_51),
.B1(n_31),
.B2(n_20),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_76),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_1),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_1),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_43),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_21),
.B(n_28),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_31),
.C(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_18),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_79),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_78),
.C(n_84),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_105),
.B(n_65),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_43),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_31),
.B1(n_19),
.B2(n_43),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_86),
.B1(n_71),
.B2(n_64),
.Y(n_114)
);

NAND2x1_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_26),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_106),
.B(n_80),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_2),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_117),
.C(n_120),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_124),
.B(n_104),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_113),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_69),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_85),
.C(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_127),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_67),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_87),
.C(n_75),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_105),
.C(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_86),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_134),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_124),
.B(n_113),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_106),
.B(n_96),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_93),
.B(n_95),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_121),
.C(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_141),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_128),
.Y(n_141)
);

NAND4xp25_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_99),
.C(n_109),
.D(n_138),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_118),
.B(n_120),
.C(n_110),
.D(n_117),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_145),
.C(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_R g145 ( 
.A(n_137),
.B(n_102),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_140),
.C(n_141),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_136),
.B(n_135),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_150),
.B(n_132),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_136),
.B(n_135),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_114),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.C(n_87),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_119),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_147),
.B(n_12),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_4),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_155),
.C(n_154),
.Y(n_163)
);

OAI31xp33_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_14),
.A3(n_6),
.B(n_7),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_159),
.B1(n_4),
.B2(n_8),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_163),
.C(n_26),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_26),
.B1(n_162),
.B2(n_146),
.C(n_96),
.Y(n_166)
);


endmodule