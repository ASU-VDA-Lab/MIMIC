module fake_jpeg_28032_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

OR2x2_ASAP7_75t_L g6 ( 
.A(n_5),
.B(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_1),
.C(n_7),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_20),
.B(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_1),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_22),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_9),
.B1(n_19),
.B2(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_15),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_9),
.B1(n_25),
.B2(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_26),
.C(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_36),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_38),
.Y(n_40)
);


endmodule