module real_jpeg_31874_n_19 (n_17, n_8, n_0, n_141, n_2, n_142, n_143, n_10, n_9, n_12, n_152, n_147, n_146, n_6, n_151, n_11, n_14, n_7, n_18, n_3, n_145, n_144, n_5, n_4, n_150, n_1, n_148, n_149, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_141;
input n_2;
input n_142;
input n_143;
input n_10;
input n_9;
input n_12;
input n_152;
input n_147;
input n_146;
input n_6;
input n_151;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_150;
input n_1;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_0),
.B(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_89),
.A3(n_91),
.B1(n_96),
.B2(n_121),
.C1(n_123),
.C2(n_152),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_18),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_49),
.C(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_5),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_6),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_109),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_10),
.B(n_37),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_98),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_15),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_15),
.Y(n_135)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_17),
.B(n_132),
.Y(n_131)
);

OAI31xp33_ASAP7_75t_L g48 ( 
.A1(n_18),
.A2(n_49),
.A3(n_51),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_137),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_129),
.B(n_134),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_33),
.B(n_127),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_24),
.B(n_32),
.Y(n_128)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_31),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_43),
.B(n_126),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_42),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI31xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_82),
.A3(n_107),
.B(n_115),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_76),
.C(n_77),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_66),
.B(n_75),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_47)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_141),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_143),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_74),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_95),
.C(n_102),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_116),
.B(n_120),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_102),
.C(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_148),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_117),
.B(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_142),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_144),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_145),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_146),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_147),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_149),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_150),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_151),
.Y(n_110)
);


endmodule