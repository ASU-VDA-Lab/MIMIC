module fake_netlist_1_12273_n_586 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_586);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_586;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_169;
wire n_424;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g167 ( .A(n_71), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_35), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_68), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_34), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_11), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_30), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_3), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_32), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_84), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_110), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_69), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_86), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_54), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_124), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_59), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_91), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_19), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_123), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_28), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_107), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_58), .Y(n_187) );
NOR2xp67_ASAP7_75t_L g188 ( .A(n_50), .B(n_136), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_131), .Y(n_189) );
INVx1_ASAP7_75t_SL g190 ( .A(n_153), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_3), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_126), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_96), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_45), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_122), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_97), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_164), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_83), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_13), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_21), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_1), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_85), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_72), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_154), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_108), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_16), .Y(n_208) );
BUFx10_ASAP7_75t_L g209 ( .A(n_6), .Y(n_209) );
INVx1_ASAP7_75t_SL g210 ( .A(n_89), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_15), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_88), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_51), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_155), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_20), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_2), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_57), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_127), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_2), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_144), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_13), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_12), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_79), .Y(n_224) );
BUFx5_ASAP7_75t_L g225 ( .A(n_76), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_44), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_111), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_104), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_132), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_80), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_116), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_39), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_7), .Y(n_233) );
INVxp33_ASAP7_75t_L g234 ( .A(n_103), .Y(n_234) );
XOR2xp5_ASAP7_75t_L g235 ( .A(n_160), .B(n_163), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_67), .Y(n_236) );
INVxp67_ASAP7_75t_L g237 ( .A(n_42), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_48), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_113), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_106), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_92), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_112), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_125), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_129), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_90), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_77), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_82), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_81), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_52), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_47), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_5), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_46), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_156), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_247), .B(n_0), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_216), .B(n_1), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_196), .B(n_4), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_168), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_168), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g262 ( .A(n_225), .B(n_166), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_168), .Y(n_263) );
OAI22x1_ASAP7_75t_R g264 ( .A1(n_173), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_183), .B(n_7), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_189), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_184), .B(n_8), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
AND2x6_ASAP7_75t_L g269 ( .A(n_172), .B(n_17), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_231), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_187), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_209), .Y(n_272) );
BUFx8_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_171), .B(n_8), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_214), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_174), .A2(n_95), .B(n_165), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
INVx4_ASAP7_75t_L g278 ( .A(n_169), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_274), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_274), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_259), .B(n_225), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_270), .A2(n_243), .B1(n_254), .B2(n_219), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_271), .B(n_225), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_258), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_269), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_271), .B(n_225), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
NAND2xp33_ASAP7_75t_L g291 ( .A(n_269), .B(n_191), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_260), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_271), .B(n_185), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_256), .A2(n_176), .B(n_175), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_256), .A2(n_235), .B1(n_201), .B2(n_203), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_273), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g302 ( .A(n_282), .B(n_271), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_283), .B(n_278), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_267), .B(n_262), .C(n_217), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_295), .B(n_288), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_294), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_280), .B(n_278), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_301), .B(n_277), .Y(n_312) );
INVx5_ASAP7_75t_L g313 ( .A(n_295), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_301), .B(n_257), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_298), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_281), .B(n_177), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_293), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_272), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_293), .B(n_268), .Y(n_323) );
AND2x6_ASAP7_75t_SL g324 ( .A(n_297), .B(n_264), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_291), .B(n_273), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_308), .A2(n_291), .B(n_276), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_309), .A2(n_276), .B(n_238), .Y(n_327) );
NOR2xp33_ASAP7_75t_SL g328 ( .A(n_315), .B(n_275), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_313), .B(n_170), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_305), .A2(n_220), .B(n_223), .C(n_192), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_307), .A2(n_193), .B(n_182), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_305), .A2(n_252), .B(n_233), .C(n_186), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_310), .A2(n_266), .B1(n_232), .B2(n_248), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_316), .A2(n_266), .B1(n_234), .B2(n_222), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_318), .Y(n_335) );
AOI21x1_ASAP7_75t_L g336 ( .A1(n_319), .A2(n_296), .B(n_290), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_306), .B(n_228), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_306), .A2(n_228), .B1(n_237), .B2(n_210), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_311), .B(n_237), .Y(n_339) );
NOR3xp33_ASAP7_75t_L g340 ( .A(n_322), .B(n_195), .C(n_194), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_312), .B(n_167), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_323), .B(n_167), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_319), .A2(n_204), .B(n_198), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_323), .B(n_321), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_321), .B(n_190), .Y(n_347) );
AOI21x1_ASAP7_75t_SL g348 ( .A1(n_337), .A2(n_325), .B(n_302), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_188), .B(n_206), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_335), .Y(n_350) );
BUFx8_ASAP7_75t_L g351 ( .A(n_344), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_320), .B(n_317), .Y(n_352) );
AO31x2_ASAP7_75t_L g353 ( .A1(n_338), .A2(n_246), .A3(n_226), .B(n_227), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_330), .B(n_324), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_334), .A2(n_222), .B1(n_239), .B2(n_255), .C(n_230), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_346), .A2(n_313), .B(n_304), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_335), .Y(n_357) );
NAND3x1_ASAP7_75t_L g358 ( .A(n_328), .B(n_212), .C(n_208), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_336), .A2(n_218), .B(n_213), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_345), .A2(n_303), .B(n_250), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_341), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_340), .A2(n_251), .B(n_253), .C(n_244), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_SL g364 ( .A1(n_332), .A2(n_190), .B(n_210), .C(n_241), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_340), .B(n_222), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_342), .A2(n_202), .B(n_197), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_SL g369 ( .A1(n_329), .A2(n_241), .B(n_224), .C(n_229), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
AO31x2_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_205), .A3(n_292), .B(n_287), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_339), .A2(n_300), .B(n_299), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_351), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_350), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_370), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_370), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_349), .A2(n_240), .B(n_236), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_360), .B(n_9), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_366), .A2(n_249), .B1(n_245), .B2(n_242), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_372), .A2(n_22), .B(n_18), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_24), .B(n_23), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_26), .B(n_25), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_368), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_371), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_371), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_357), .B(n_10), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_109), .B(n_162), .Y(n_388) );
AOI21x1_ASAP7_75t_L g389 ( .A1(n_365), .A2(n_367), .B(n_361), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_354), .B(n_11), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_371), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_221), .B(n_215), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_364), .A2(n_105), .B(n_161), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_353), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_353), .B(n_14), .Y(n_397) );
AO31x2_ASAP7_75t_L g398 ( .A1(n_370), .A2(n_15), .A3(n_27), .B(n_29), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_362), .B(n_178), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_31), .B(n_33), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_200), .B(n_199), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_359), .A2(n_181), .B(n_180), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_363), .A2(n_179), .B(n_37), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g404 ( .A(n_355), .B(n_36), .C(n_38), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_368), .B(n_40), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_352), .A2(n_41), .B(n_43), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_384), .B(n_49), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_395), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
OAI21x1_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_406), .B(n_400), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_53), .B(n_55), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx5_ASAP7_75t_SL g415 ( .A(n_375), .Y(n_415) );
INVx5_ASAP7_75t_L g416 ( .A(n_375), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_56), .B(n_60), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_392), .B(n_61), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_390), .B(n_159), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_377), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_399), .B(n_62), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_391), .A2(n_63), .B(n_64), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_403), .A2(n_65), .B(n_66), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_378), .A2(n_70), .B(n_73), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_397), .A2(n_74), .B1(n_75), .B2(n_78), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_375), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_373), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_380), .B(n_87), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
BUFx2_ASAP7_75t_SL g443 ( .A(n_401), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_402), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_393), .A2(n_93), .B1(n_94), .B2(n_98), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_392), .B(n_99), .Y(n_448) );
INVxp33_ASAP7_75t_SL g449 ( .A(n_374), .Y(n_449) );
INVxp33_ASAP7_75t_L g450 ( .A(n_375), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_376), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_384), .B(n_100), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_375), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_376), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_384), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_409), .B(n_101), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_455), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_409), .B(n_102), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_448), .B(n_432), .Y(n_459) );
NOR2x1_ASAP7_75t_SL g460 ( .A(n_421), .B(n_114), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_414), .B(n_158), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_449), .B(n_115), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_423), .B(n_117), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_449), .B(n_118), .Y(n_466) );
BUFx2_ASAP7_75t_SL g467 ( .A(n_434), .Y(n_467) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_440), .A2(n_119), .B(n_120), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_451), .B(n_121), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_451), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_454), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_416), .Y(n_473) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_410), .A2(n_128), .B(n_130), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_424), .B(n_133), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_408), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_413), .B(n_157), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_416), .B(n_134), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_407), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_452), .B(n_135), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_436), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_432), .B(n_137), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_450), .B(n_138), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_416), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_427), .A2(n_140), .B1(n_143), .B2(n_145), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_450), .B(n_146), .Y(n_493) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_453), .B(n_147), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_415), .B(n_149), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_419), .B(n_150), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_444), .B(n_152), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_445), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_446), .A2(n_422), .B1(n_442), .B2(n_429), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_442), .B(n_443), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_470), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_477), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_481), .B(n_428), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_462), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_477), .B(n_467), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_487), .B(n_446), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_471), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_472), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_499), .Y(n_513) );
OAI222xp33_ASAP7_75t_L g514 ( .A1(n_500), .A2(n_429), .B1(n_439), .B2(n_446), .C1(n_438), .C2(n_435), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_412), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_490), .B(n_417), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_492), .B(n_417), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_489), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_484), .B(n_426), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_478), .B(n_426), .Y(n_526) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_502), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_501), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_459), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_464), .B(n_437), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_461), .B(n_437), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_494), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_494), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_528), .B(n_459), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_509), .B(n_469), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_515), .B(n_476), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_522), .B(n_465), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_503), .B(n_479), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_513), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_504), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_505), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_507), .B(n_465), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_505), .B(n_458), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_508), .B(n_456), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_521), .B(n_456), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_523), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_503), .B(n_479), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_521), .B(n_493), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_516), .B(n_494), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_506), .B(n_486), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g552 ( .A(n_529), .B(n_466), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_524), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_541), .B(n_529), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_540), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_535), .B(n_551), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_546), .B(n_512), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_539), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_547), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_552), .A2(n_526), .B1(n_520), .B2(n_510), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_553), .B(n_511), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_534), .B(n_520), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_560), .A2(n_538), .B(n_548), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_559), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
NAND2x1_ASAP7_75t_L g567 ( .A(n_562), .B(n_550), .Y(n_567) );
AOI222xp33_ASAP7_75t_L g568 ( .A1(n_565), .A2(n_561), .B1(n_557), .B2(n_560), .C1(n_556), .C2(n_514), .Y(n_568) );
XNOR2x1_ASAP7_75t_L g569 ( .A(n_567), .B(n_549), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_564), .B(n_558), .Y(n_570) );
AOI221x1_ASAP7_75t_L g571 ( .A1(n_563), .A2(n_537), .B1(n_536), .B2(n_542), .C(n_544), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_568), .B(n_566), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_571), .B(n_530), .C(n_543), .D(n_545), .Y(n_573) );
OAI211xp5_ASAP7_75t_SL g574 ( .A1(n_572), .A2(n_570), .B(n_569), .C(n_496), .Y(n_574) );
OAI21xp33_ASAP7_75t_SL g575 ( .A1(n_573), .A2(n_525), .B(n_527), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_575), .A2(n_491), .B(n_497), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_574), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_577), .B(n_460), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_578), .B(n_576), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_579), .B(n_527), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_485), .B(n_495), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_581), .A2(n_482), .B1(n_533), .B2(n_531), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_447), .B(n_474), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_532), .B1(n_498), .B2(n_517), .C1(n_519), .C2(n_518), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_584), .B(n_468), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_447), .B(n_468), .Y(n_586) );
endmodule