module fake_jpeg_1748_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_54),
.Y(n_96)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_22),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_63),
.Y(n_95)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_3),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_87),
.Y(n_137)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_3),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_69),
.Y(n_119)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_79),
.Y(n_100)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_27),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_76),
.Y(n_124)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_23),
.B(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_6),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_36),
.B1(n_34),
.B2(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_97),
.A2(n_121),
.B1(n_138),
.B2(n_140),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_36),
.B1(n_43),
.B2(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_101),
.A2(n_103),
.B1(n_111),
.B2(n_118),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_87),
.B1(n_84),
.B2(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_48),
.A2(n_59),
.B1(n_41),
.B2(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_49),
.B(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_8),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_24),
.B1(n_41),
.B2(n_39),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_54),
.A2(n_74),
.B1(n_62),
.B2(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_35),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_43),
.B1(n_26),
.B2(n_39),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_40),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_38),
.B1(n_32),
.B2(n_30),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_111),
.B1(n_101),
.B2(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_38),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_52),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_46),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_72),
.A2(n_40),
.B1(n_20),
.B2(n_21),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_98),
.B1(n_119),
.B2(n_93),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_51),
.A2(n_40),
.B1(n_20),
.B2(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_58),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_153),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_7),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_149),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_148),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_40),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_47),
.B(n_40),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_125),
.C(n_114),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_8),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_20),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_165),
.B1(n_175),
.B2(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_9),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_11),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_163),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_167),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_13),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_14),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_15),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_176),
.Y(n_211)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_20),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_173),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_108),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_129),
.B(n_117),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_106),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_134),
.B1(n_93),
.B2(n_108),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_193),
.B1(n_202),
.B2(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_132),
.B1(n_125),
.B2(n_109),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_109),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_213),
.C(n_151),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_161),
.B(n_166),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_162),
.B1(n_147),
.B2(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_200),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_123),
.B1(n_141),
.B2(n_132),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_122),
.B1(n_114),
.B2(n_123),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_154),
.B1(n_165),
.B2(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_184),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_122),
.B1(n_141),
.B2(n_153),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_144),
.B(n_168),
.C(n_170),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_223),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_180),
.B(n_181),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_226),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_176),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_235),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_160),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_231),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_229),
.B(n_236),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_177),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_159),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_175),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

XOR2x1_ASAP7_75t_SL g236 ( 
.A(n_204),
.B(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_186),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_239),
.A2(n_194),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_199),
.B1(n_207),
.B2(n_197),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_195),
.C(n_190),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_255),
.C(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_251),
.B(n_223),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_203),
.C(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_215),
.C(n_206),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_200),
.B1(n_193),
.B2(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_220),
.B1(n_229),
.B2(n_228),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_211),
.B(n_188),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_229),
.B(n_226),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_221),
.B1(n_227),
.B2(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_266),
.B1(n_270),
.B2(n_249),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_247),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

OAI322xp33_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_224),
.A3(n_219),
.B1(n_225),
.B2(n_232),
.C1(n_236),
.C2(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_259),
.C(n_268),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_239),
.C(n_229),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_269),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_228),
.B1(n_234),
.B2(n_220),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_257),
.B1(n_243),
.B2(n_241),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_274),
.B(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_238),
.B1(n_237),
.B2(n_233),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_218),
.B1(n_217),
.B2(n_240),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_252),
.B1(n_254),
.B2(n_253),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_279),
.B(n_281),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_245),
.B1(n_244),
.B2(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_257),
.B1(n_256),
.B2(n_254),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_265),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_248),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_277),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_265),
.C(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.C(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_260),
.C(n_273),
.Y(n_288)
);

AOI321xp33_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_274),
.A3(n_269),
.B1(n_270),
.B2(n_264),
.C(n_248),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_278),
.B1(n_276),
.B2(n_283),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.C(n_288),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_280),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_298),
.C(n_300),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_302),
.A2(n_214),
.B(n_209),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_209),
.Y(n_304)
);


endmodule