module fake_jpeg_12226_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_7),
.B1(n_2),
.B2(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_11),
.B1(n_13),
.B2(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_8),
.B1(n_11),
.B2(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_5),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_21),
.B1(n_10),
.B2(n_23),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_37),
.B1(n_28),
.B2(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_15),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_28),
.B(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_32),
.B(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_37),
.B1(n_36),
.B2(n_26),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_31),
.C(n_33),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_46),
.C(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_39),
.B1(n_40),
.B2(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_47),
.A3(n_45),
.B1(n_46),
.B2(n_6),
.C1(n_5),
.C2(n_15),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_51),
.B1(n_5),
.B2(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);


endmodule