module fake_jpeg_11465_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_23),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_45),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_9),
.B(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_34),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_1),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_72),
.Y(n_95)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_64),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_74),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_103),
.C(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_55),
.B1(n_52),
.B2(n_56),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_108),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_90),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_85),
.B1(n_52),
.B2(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_20),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_53),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_85),
.B1(n_62),
.B2(n_63),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_119),
.Y(n_135)
);

BUFx2_ASAP7_75t_SL g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_63),
.B1(n_75),
.B2(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_57),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_61),
.Y(n_136)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_76),
.B1(n_65),
.B2(n_60),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_79),
.B1(n_78),
.B2(n_26),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_75),
.B1(n_70),
.B2(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_143),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_36),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_71),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_141),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_68),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_145),
.B1(n_8),
.B2(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_3),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_22),
.C(n_49),
.Y(n_144)
);

XOR2x1_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_32),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_28),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_161),
.C(n_162),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_164),
.C(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_128),
.B1(n_133),
.B2(n_148),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_12),
.B(n_13),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_157),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_33),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_131),
.C(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_131),
.C(n_140),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_158),
.B1(n_159),
.B2(n_151),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_152),
.C(n_157),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_173),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_172),
.C(n_175),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_158),
.C(n_170),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_163),
.B(n_159),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_137),
.B1(n_41),
.B2(n_43),
.C(n_44),
.Y(n_182)
);


endmodule