module fake_jpeg_14080_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_15),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_19),
.B1(n_27),
.B2(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_73),
.B1(n_44),
.B2(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_46),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_63),
.B1(n_66),
.B2(n_22),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_75),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_70),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_28),
.B1(n_35),
.B2(n_17),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_33),
.B1(n_24),
.B2(n_40),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_17),
.B1(n_35),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_69),
.B1(n_71),
.B2(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_17),
.B1(n_35),
.B2(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_36),
.B(n_34),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_17),
.B1(n_35),
.B2(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_45),
.B1(n_41),
.B2(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_22),
.B1(n_20),
.B2(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_24),
.B1(n_23),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_90),
.B1(n_69),
.B2(n_71),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_45),
.B(n_18),
.C(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_39),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_108),
.C(n_56),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_83),
.A2(n_72),
.B1(n_64),
.B2(n_50),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_75),
.B1(n_48),
.B2(n_64),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_92),
.B1(n_57),
.B2(n_50),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_26),
.B1(n_22),
.B2(n_34),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_74),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_9),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_104),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_74),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_0),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_9),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_48),
.B(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_0),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_30),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_82),
.Y(n_159)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_125),
.B1(n_128),
.B2(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_87),
.A2(n_71),
.B1(n_49),
.B2(n_75),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_50),
.B1(n_93),
.B2(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_137),
.B(n_110),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_89),
.B(n_57),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_105),
.B(n_80),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_142),
.B(n_21),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_131),
.B(n_138),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_119),
.B(n_139),
.Y(n_178)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_81),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_78),
.B1(n_106),
.B2(n_97),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_165),
.B1(n_122),
.B2(n_125),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_152),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_85),
.B(n_107),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_121),
.B(n_133),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_78),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_89),
.C(n_107),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_158),
.B(n_160),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_95),
.C(n_82),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_13),
.C(n_12),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_84),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_109),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_120),
.B1(n_103),
.B2(n_93),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_104),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_116),
.B(n_91),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_174),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_133),
.B1(n_101),
.B2(n_77),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_79),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_116),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_202),
.C(n_162),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_113),
.CI(n_127),
.CON(n_176),
.SN(n_176)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_176),
.B(n_161),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_183),
.B(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_192),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_112),
.B(n_126),
.C(n_121),
.D(n_101),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_121),
.B(n_133),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_201),
.B(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_169),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_31),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_154),
.B(n_159),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_199),
.B1(n_204),
.B2(n_159),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_142),
.B(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_120),
.B1(n_21),
.B2(n_13),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_0),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_31),
.B(n_30),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_145),
.B1(n_156),
.B2(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_12),
.B1(n_11),
.B2(n_30),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_205),
.A2(n_172),
.B1(n_161),
.B2(n_152),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_1),
.B(n_2),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_209),
.Y(n_258)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_172),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_224),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_213),
.B(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_236),
.B1(n_182),
.B2(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_174),
.C(n_164),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_222),
.C(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_189),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g221 ( 
.A1(n_178),
.A2(n_146),
.B(n_157),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_157),
.C(n_143),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_196),
.C(n_187),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_143),
.C(n_2),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_235),
.C(n_193),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

AOI22x1_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_205),
.B1(n_183),
.B2(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_1),
.C(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_180),
.B(n_1),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_255),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_176),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_244),
.C(n_253),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_211),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_197),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_252),
.B(n_235),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_182),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_216),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_193),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_260),
.C(n_226),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_217),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_194),
.B1(n_214),
.B2(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_219),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_246),
.A2(n_229),
.B1(n_234),
.B2(n_211),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_267),
.A2(n_230),
.B1(n_177),
.B2(n_5),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_276),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_274),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_258),
.B1(n_237),
.B2(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_223),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_210),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_203),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_229),
.C(n_227),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.C(n_244),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_227),
.C(n_201),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_243),
.B(n_259),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_293),
.B(n_272),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_245),
.B1(n_238),
.B2(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_250),
.C(n_240),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_253),
.C(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_245),
.C(n_203),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_230),
.B(n_245),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_292),
.C(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_291),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_265),
.C(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_264),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_262),
.C(n_267),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_309),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_177),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_287),
.B(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_282),
.C(n_284),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_301),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_266),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_312),
.Y(n_324)
);

AOI221xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_275),
.B1(n_273),
.B2(n_296),
.C(n_274),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_4),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_3),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_306),
.C(n_303),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_325),
.B(n_313),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_4),
.C(n_5),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_326),
.Y(n_328)
);

AO221x1_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_325),
.B1(n_330),
.B2(n_328),
.C(n_317),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_315),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_321),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_316),
.C(n_6),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_5),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_7),
.Y(n_337)
);


endmodule