module fake_aes_8780_n_1059 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1059);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1059;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_844;
wire n_818;
wire n_230;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_235;
wire n_482;
wire n_243;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_947;
wire n_912;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
AND2x2_ASAP7_75t_L g227 ( .A(n_50), .B(n_208), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_41), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_141), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_133), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_60), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_63), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_9), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_114), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_84), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_107), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_126), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_85), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_45), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_66), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_12), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_151), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_213), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_136), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_172), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_42), .B(n_105), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_94), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_16), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_135), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_97), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_24), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_137), .Y(n_258) );
INVx4_ASAP7_75t_R g259 ( .A(n_7), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_80), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_164), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_71), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_26), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_155), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_4), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_54), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_166), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_142), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_72), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_150), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_50), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_99), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_104), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_113), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_15), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_196), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g279 ( .A(n_122), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_132), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_206), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_214), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_5), .Y(n_283) );
CKINVDCx14_ASAP7_75t_R g284 ( .A(n_17), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_74), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_144), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_40), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_111), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_118), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_69), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_188), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_65), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_58), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_31), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_129), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_218), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_224), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_6), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_64), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_158), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_162), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_153), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_109), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_19), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_156), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_53), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_186), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_199), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_217), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_226), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_22), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_167), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_91), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_182), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_75), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_55), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_194), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_21), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_2), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_47), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_154), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_101), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_79), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_203), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_205), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_215), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_98), .Y(n_328) );
INVxp33_ASAP7_75t_SL g329 ( .A(n_148), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_124), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_121), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_48), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_47), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_170), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_180), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_225), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_8), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_139), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_20), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_42), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_56), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_125), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_168), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_312), .B(n_0), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_248), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_337), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_337), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_337), .B(n_0), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_284), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_228), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_228), .Y(n_351) );
INVx6_ASAP7_75t_L g352 ( .A(n_248), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_245), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_284), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_257), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_245), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_266), .B(n_1), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_301), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_305), .Y(n_360) );
AND2x6_ASAP7_75t_L g361 ( .A(n_311), .B(n_59), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_266), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_230), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_300), .B(n_3), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_248), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_229), .B(n_4), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_233), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_238), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_227), .B(n_61), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_291), .B(n_5), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_238), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_240), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_267), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_240), .Y(n_375) );
CKINVDCx6p67_ASAP7_75t_R g376 ( .A(n_313), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_345), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_364), .B(n_315), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_346), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_364), .B(n_236), .Y(n_381) );
BUFx4f_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_361), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_361), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_376), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_371), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_345), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_364), .B(n_242), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_346), .B(n_246), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_376), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_358), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_348), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_363), .B(n_261), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_363), .B(n_296), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_347), .B(n_246), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_347), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_279), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_279), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_361), .B(n_232), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_371), .Y(n_408) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_354), .A2(n_319), .B1(n_317), .B2(n_268), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_367), .B(n_252), .Y(n_411) );
BUFx10_ASAP7_75t_L g412 ( .A(n_361), .Y(n_412) );
INVx4_ASAP7_75t_L g413 ( .A(n_361), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_351), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_345), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_357), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_351), .B(n_231), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_351), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_345), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_378), .A2(n_371), .B1(n_357), .B2(n_366), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_416), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_379), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_412), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_380), .B(n_357), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_380), .B(n_370), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_417), .B(n_370), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_384), .B(n_231), .Y(n_429) );
INVx5_ASAP7_75t_L g430 ( .A(n_416), .Y(n_430) );
BUFx4f_ASAP7_75t_L g431 ( .A(n_408), .Y(n_431) );
NOR3xp33_ASAP7_75t_SL g432 ( .A(n_392), .B(n_339), .C(n_344), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_416), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_378), .B(n_371), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_384), .B(n_232), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_417), .B(n_368), .Y(n_436) );
AND2x6_ASAP7_75t_L g437 ( .A(n_385), .B(n_342), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_404), .B(n_368), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_404), .B(n_368), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_387), .A2(n_237), .B1(n_270), .B2(n_265), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
NAND2xp33_ASAP7_75t_SL g453 ( .A(n_386), .B(n_237), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_393), .B(n_368), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
NOR2xp33_ASAP7_75t_SL g456 ( .A(n_395), .B(n_265), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_396), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_406), .A2(n_270), .B1(n_298), .B2(n_290), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_393), .B(n_362), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_397), .B(n_355), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_381), .B(n_290), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_391), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_381), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_409), .A2(n_374), .B1(n_267), .B2(n_307), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_410), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_381), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_389), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_382), .A2(n_373), .B(n_372), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_394), .B(n_369), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_418), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_394), .B(n_369), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_398), .B(n_307), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_396), .B(n_369), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_396), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_389), .B(n_310), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_411), .Y(n_481) );
NOR2xp33_ASAP7_75t_R g482 ( .A(n_399), .B(n_318), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
NOR3xp33_ASAP7_75t_SL g484 ( .A(n_411), .B(n_263), .C(n_249), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_399), .A2(n_372), .B(n_375), .C(n_373), .Y(n_485) );
O2A1O1Ixp5_ASAP7_75t_L g486 ( .A1(n_382), .A2(n_322), .B(n_235), .C(n_239), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_399), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_423), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_434), .A2(n_382), .B1(n_413), .B2(n_395), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_443), .A2(n_382), .B(n_400), .C(n_390), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_458), .A2(n_390), .B1(n_400), .B2(n_413), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_427), .B(n_409), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_462), .B(n_409), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g496 ( .A1(n_465), .A2(n_329), .B1(n_254), .B2(n_264), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_445), .A2(n_385), .B(n_369), .C(n_375), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_422), .Y(n_498) );
NAND2xp33_ASAP7_75t_L g499 ( .A(n_424), .B(n_413), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_434), .B(n_412), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_482), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_462), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_430), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_447), .A2(n_277), .B(n_283), .C(n_272), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_478), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_421), .A2(n_295), .B(n_299), .C(n_288), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_448), .B(n_263), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_449), .A2(n_321), .B1(n_332), .B2(n_320), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_449), .B(n_353), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_460), .B(n_333), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_430), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g515 ( .A(n_420), .B(n_62), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_424), .Y(n_516) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_480), .B(n_340), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_426), .B(n_294), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_426), .B(n_306), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_463), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_428), .A2(n_341), .B1(n_241), .B2(n_243), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_425), .A2(n_244), .B(n_234), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_474), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_477), .B(n_323), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_436), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_464), .A2(n_356), .B1(n_359), .B2(n_353), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_439), .A2(n_359), .B(n_360), .C(n_356), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_450), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_467), .B(n_360), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_453), .Y(n_532) );
AOI221x1_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_303), .B1(n_253), .B2(n_255), .C(n_256), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_431), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_476), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_450), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_424), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_437), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_431), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_440), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_425), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_432), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_457), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_479), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_479), .B(n_314), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_438), .A2(n_258), .B(n_247), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_446), .Y(n_549) );
INVx4_ASAP7_75t_L g550 ( .A(n_437), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_483), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_435), .A2(n_262), .B1(n_269), .B2(n_260), .Y(n_552) );
AO22x1_ASAP7_75t_L g553 ( .A1(n_435), .A2(n_278), .B1(n_259), .B2(n_343), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_455), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_456), .A2(n_273), .B1(n_274), .B2(n_271), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_436), .A2(n_280), .B(n_281), .C(n_276), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_442), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_451), .Y(n_560) );
NAND2x2_ASAP7_75t_L g561 ( .A(n_456), .B(n_342), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_452), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_438), .B(n_282), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_437), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_429), .B(n_285), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_459), .A2(n_454), .B(n_444), .C(n_486), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_444), .A2(n_289), .B(n_287), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_459), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_466), .B(n_468), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_470), .Y(n_570) );
CKINVDCx6p67_ASAP7_75t_R g571 ( .A(n_437), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_472), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_440), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_454), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_475), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_471), .B(n_292), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_461), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_461), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_461), .A2(n_297), .B(n_293), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_481), .B(n_302), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_430), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_SL g583 ( .A1(n_491), .A2(n_308), .B(n_309), .C(n_304), .Y(n_583) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_515), .A2(n_268), .B(n_252), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_507), .A2(n_275), .B(n_316), .C(n_286), .Y(n_585) );
BUFx10_ASAP7_75t_L g586 ( .A(n_489), .Y(n_586) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_566), .A2(n_316), .B(n_324), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_558), .Y(n_588) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_569), .A2(n_326), .B(n_325), .Y(n_589) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_572), .A2(n_328), .B(n_327), .Y(n_590) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_533), .A2(n_338), .A3(n_331), .B(n_334), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_504), .B(n_335), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_534), .B(n_336), .Y(n_593) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_572), .A2(n_383), .B(n_377), .Y(n_594) );
OAI21x1_ASAP7_75t_SL g595 ( .A1(n_550), .A2(n_8), .B(n_9), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_543), .B(n_250), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_488), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_557), .A2(n_248), .B(n_251), .C(n_330), .Y(n_598) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_578), .A2(n_383), .B(n_377), .Y(n_599) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_578), .A2(n_401), .B(n_388), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_531), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_540), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_503), .B(n_10), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_568), .B(n_11), .Y(n_605) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_488), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_531), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_504), .Y(n_608) );
AO31x2_ASAP7_75t_L g609 ( .A1(n_497), .A2(n_415), .A3(n_401), .B(n_388), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_524), .B(n_11), .Y(n_610) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_580), .A2(n_415), .B(n_330), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_513), .B(n_12), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_570), .Y(n_614) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_549), .A2(n_415), .B(n_330), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_522), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_496), .A2(n_352), .B1(n_330), .B2(n_251), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_510), .A2(n_251), .B1(n_352), .B2(n_365), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_548), .A2(n_419), .B(n_251), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_488), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_494), .B(n_13), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_492), .Y(n_623) );
CKINVDCx9p33_ASAP7_75t_R g624 ( .A(n_559), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_567), .A2(n_419), .B(n_365), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
OAI21x1_ASAP7_75t_SL g628 ( .A1(n_550), .A2(n_13), .B(n_14), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_552), .B(n_365), .C(n_419), .Y(n_629) );
OAI21x1_ASAP7_75t_L g630 ( .A1(n_554), .A2(n_68), .B(n_67), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_523), .A2(n_352), .B(n_14), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_492), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_492), .Y(n_633) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_551), .A2(n_73), .B(n_70), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_530), .B(n_17), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_535), .A2(n_352), .B(n_18), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_498), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_536), .B(n_18), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_552), .B(n_419), .C(n_19), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_520), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_528), .Y(n_641) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_556), .A2(n_419), .B(n_77), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_512), .A2(n_20), .B(n_21), .Y(n_643) );
AO32x2_ASAP7_75t_L g644 ( .A1(n_496), .A2(n_22), .A3(n_23), .B1(n_24), .B2(n_25), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_506), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_495), .B(n_27), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_514), .A2(n_27), .B(n_28), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_555), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_502), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_582), .Y(n_650) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_579), .A2(n_78), .B(n_76), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_501), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_526), .B(n_28), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_563), .A2(n_82), .B(n_81), .Y(n_654) );
CKINVDCx6p67_ASAP7_75t_R g655 ( .A(n_544), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_582), .A2(n_86), .B(n_83), .Y(n_656) );
BUFx2_ASAP7_75t_SL g657 ( .A(n_539), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_511), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_509), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_517), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_529), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_516), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_577), .Y(n_663) );
OA21x2_ASAP7_75t_L g664 ( .A1(n_515), .A2(n_88), .B(n_87), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_505), .A2(n_29), .B(n_30), .C(n_32), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_490), .A2(n_145), .B(n_223), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_525), .B(n_32), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_546), .Y(n_668) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_493), .A2(n_577), .B(n_521), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_527), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_526), .B(n_33), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_575), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_553), .B(n_33), .Y(n_673) );
OAI21x1_ASAP7_75t_L g674 ( .A1(n_537), .A2(n_146), .B(n_222), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_532), .B(n_34), .Y(n_675) );
OA21x2_ASAP7_75t_L g676 ( .A1(n_521), .A2(n_143), .B(n_221), .Y(n_676) );
AO31x2_ASAP7_75t_L g677 ( .A1(n_565), .A2(n_35), .A3(n_36), .B(n_37), .Y(n_677) );
NAND3xp33_ASAP7_75t_SL g678 ( .A(n_508), .B(n_35), .C(n_36), .Y(n_678) );
OR2x6_ASAP7_75t_L g679 ( .A(n_564), .B(n_37), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_541), .A2(n_149), .B(n_220), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_518), .A2(n_147), .B(n_219), .Y(n_681) );
OR2x6_ASAP7_75t_L g682 ( .A(n_500), .B(n_38), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_519), .A2(n_140), .B(n_216), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_561), .A2(n_39), .B1(n_41), .B2(n_43), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_545), .Y(n_685) );
BUFx4f_ASAP7_75t_SL g686 ( .A(n_655), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_645), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_649), .Y(n_688) );
CKINVDCx12_ASAP7_75t_R g689 ( .A(n_679), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_588), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_616), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_658), .A2(n_547), .B1(n_571), .B2(n_539), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_672), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_617), .A2(n_573), .B(n_542), .C(n_538), .Y(n_694) );
AO21x2_ASAP7_75t_L g695 ( .A1(n_587), .A2(n_499), .B(n_542), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_622), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_667), .A2(n_573), .B(n_538), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_604), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_626), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_613), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_669), .A2(n_39), .B(n_43), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_672), .B(n_44), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_605), .A2(n_45), .B1(n_46), .B2(n_48), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_606), .Y(n_704) );
CKINVDCx8_ASAP7_75t_R g705 ( .A(n_673), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_627), .A2(n_49), .B(n_51), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_614), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_648), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_625), .A2(n_159), .B(n_211), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_679), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_625), .A2(n_160), .B(n_210), .Y(n_711) );
OR2x6_ASAP7_75t_L g712 ( .A(n_682), .B(n_56), .Y(n_712) );
OR2x6_ASAP7_75t_L g713 ( .A(n_682), .B(n_57), .Y(n_713) );
AOI221xp5_ASAP7_75t_SL g714 ( .A1(n_585), .A2(n_89), .B1(n_90), .B2(n_92), .C(n_93), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_640), .B(n_95), .Y(n_715) );
BUFx8_ASAP7_75t_L g716 ( .A(n_644), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_605), .A2(n_96), .B1(n_100), .B2(n_102), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_682), .A2(n_103), .B1(n_106), .B2(n_108), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_670), .A2(n_110), .B1(n_112), .B2(n_115), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_603), .A2(n_671), .B1(n_621), .B2(n_646), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_617), .A2(n_116), .B1(n_117), .B2(n_119), .C(n_120), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_643), .A2(n_123), .B1(n_127), .B2(n_128), .C(n_130), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_597), .B(n_131), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_684), .A2(n_134), .B1(n_138), .B2(n_152), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_602), .B(n_157), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_610), .Y(n_726) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_606), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_619), .A2(n_161), .B(n_163), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_663), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_601), .B(n_607), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_596), .A2(n_178), .B1(n_183), .B2(n_184), .C(n_185), .Y(n_731) );
NAND2x1_ASAP7_75t_L g732 ( .A(n_597), .B(n_187), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_643), .A2(n_189), .B1(n_190), .B2(n_191), .C(n_192), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_637), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_673), .A2(n_193), .B1(n_195), .B2(n_197), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_678), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_610), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_684), .A2(n_204), .B1(n_207), .B2(n_209), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_659), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_635), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_586), .B(n_592), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_596), .A2(n_636), .B1(n_618), .B2(n_631), .C(n_639), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_652), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_653), .A2(n_635), .B1(n_638), .B2(n_592), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_665), .A2(n_641), .B1(n_593), .B2(n_647), .C(n_631), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_638), .B(n_685), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_612), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_675), .A2(n_647), .B1(n_660), .B2(n_608), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_620), .B(n_623), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_608), .B(n_661), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_677), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_636), .A2(n_650), .B1(n_629), .B2(n_628), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_665), .A2(n_589), .B(n_598), .C(n_629), .Y(n_753) );
BUFx6f_ASAP7_75t_L g754 ( .A(n_662), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_644), .B(n_677), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_650), .A2(n_595), .B1(n_668), .B2(n_633), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_632), .A2(n_633), .B1(n_657), .B2(n_590), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_583), .A2(n_683), .B1(n_681), .B2(n_619), .C(n_654), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_677), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_676), .A2(n_664), .B1(n_632), .B2(n_683), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_609), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_676), .A2(n_664), .B1(n_642), .B2(n_666), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_662), .B(n_681), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_L g764 ( .A1(n_654), .A2(n_642), .B(n_624), .C(n_644), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_591), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_591), .B(n_584), .Y(n_766) );
OR2x6_ASAP7_75t_L g767 ( .A(n_656), .B(n_630), .Y(n_767) );
AOI222xp33_ASAP7_75t_L g768 ( .A1(n_634), .A2(n_680), .B1(n_674), .B2(n_651), .C1(n_591), .C2(n_611), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_609), .B(n_599), .Y(n_769) );
AO21x2_ASAP7_75t_L g770 ( .A1(n_615), .A2(n_594), .B(n_600), .Y(n_770) );
INVx4_ASAP7_75t_L g771 ( .A(n_609), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_616), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_616), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_712), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_761), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_751), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_690), .B(n_698), .Y(n_777) );
AND2x4_ASAP7_75t_L g778 ( .A(n_763), .B(n_747), .Y(n_778) );
BUFx2_ASAP7_75t_L g779 ( .A(n_712), .Y(n_779) );
OR2x2_ASAP7_75t_SL g780 ( .A(n_705), .B(n_689), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_700), .B(n_707), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_734), .B(n_739), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_743), .B(n_687), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_759), .Y(n_784) );
BUFx3_ASAP7_75t_L g785 ( .A(n_704), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_765), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_763), .B(n_769), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_696), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_693), .B(n_726), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_754), .B(n_737), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_699), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_740), .B(n_746), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_713), .B(n_708), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_754), .B(n_767), .Y(n_794) );
NOR2x1_ASAP7_75t_SL g795 ( .A(n_713), .B(n_694), .Y(n_795) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_744), .A2(n_742), .B(n_745), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_713), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_691), .B(n_772), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_755), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_773), .B(n_706), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_720), .B(n_741), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_766), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_771), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_749), .B(n_730), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_771), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_770), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_704), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_750), .Y(n_808) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_704), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_716), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_716), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_767), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_767), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_695), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_703), .B(n_723), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_764), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_723), .Y(n_817) );
BUFx3_ASAP7_75t_L g818 ( .A(n_727), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_748), .B(n_701), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_760), .Y(n_820) );
AOI211xp5_ASAP7_75t_SL g821 ( .A1(n_710), .A2(n_735), .B(n_686), .C(n_738), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_760), .Y(n_822) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_727), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_732), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_702), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_727), .B(n_752), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_725), .B(n_738), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_756), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_768), .Y(n_829) );
INVx3_ASAP7_75t_L g830 ( .A(n_715), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_722), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_733), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_753), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_692), .B(n_697), .Y(n_834) );
BUFx6f_ASAP7_75t_L g835 ( .A(n_757), .Y(n_835) );
NAND2x1p5_ASAP7_75t_L g836 ( .A(n_736), .B(n_709), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_762), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_711), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_724), .B(n_717), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_718), .B(n_714), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_728), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_758), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_721), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_688), .B(n_719), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_731), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_729), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_763), .B(n_747), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_775), .Y(n_848) );
AND2x4_ASAP7_75t_SL g849 ( .A(n_815), .B(n_807), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_799), .B(n_802), .Y(n_850) );
AOI211xp5_ASAP7_75t_L g851 ( .A1(n_774), .A2(n_797), .B(n_779), .C(n_796), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_799), .B(n_802), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_829), .B(n_787), .Y(n_853) );
BUFx2_ASAP7_75t_L g854 ( .A(n_794), .Y(n_854) );
INVx4_ASAP7_75t_L g855 ( .A(n_779), .Y(n_855) );
INVx2_ASAP7_75t_SL g856 ( .A(n_794), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_829), .B(n_787), .Y(n_857) );
AOI22x1_ASAP7_75t_L g858 ( .A1(n_821), .A2(n_839), .B1(n_824), .B2(n_844), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_775), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_793), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_798), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_778), .B(n_847), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_776), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_787), .B(n_786), .Y(n_864) );
AOI33xp33_ASAP7_75t_L g865 ( .A1(n_801), .A2(n_788), .A3(n_791), .B1(n_798), .B2(n_825), .B3(n_811), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_783), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_787), .B(n_786), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_810), .B(n_789), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_776), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_783), .B(n_784), .Y(n_870) );
AND2x4_ASAP7_75t_L g871 ( .A(n_778), .B(n_847), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_789), .Y(n_872) );
INVx1_ASAP7_75t_SL g873 ( .A(n_780), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_784), .B(n_847), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_806), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_806), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_777), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_827), .A2(n_830), .B1(n_817), .B2(n_845), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_778), .B(n_847), .Y(n_879) );
INVx4_ASAP7_75t_L g880 ( .A(n_830), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_792), .B(n_804), .Y(n_881) );
OR2x6_ASAP7_75t_L g882 ( .A(n_817), .B(n_813), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_804), .B(n_792), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_827), .A2(n_830), .B1(n_845), .B2(n_843), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_777), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_781), .B(n_782), .Y(n_886) );
AOI221x1_ASAP7_75t_L g887 ( .A1(n_842), .A2(n_816), .B1(n_833), .B2(n_837), .C(n_838), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_778), .B(n_781), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_782), .B(n_833), .Y(n_889) );
INVx5_ASAP7_75t_SL g890 ( .A(n_794), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_828), .A2(n_819), .B1(n_800), .B2(n_808), .C(n_837), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_809), .B(n_823), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_845), .A2(n_843), .B1(n_808), .B2(n_846), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_800), .B(n_819), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_828), .B(n_816), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_803), .Y(n_896) );
AND2x4_ASAP7_75t_SL g897 ( .A(n_790), .B(n_794), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_812), .B(n_803), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_812), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_805), .B(n_813), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_805), .Y(n_901) );
BUFx2_ASAP7_75t_L g902 ( .A(n_814), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_814), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_820), .B(n_822), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_826), .Y(n_905) );
OR2x2_ASAP7_75t_L g906 ( .A(n_834), .B(n_835), .Y(n_906) );
AO21x2_ASAP7_75t_L g907 ( .A1(n_841), .A2(n_840), .B(n_832), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_785), .B(n_818), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_795), .Y(n_909) );
INVx3_ASAP7_75t_L g910 ( .A(n_909), .Y(n_910) );
INVxp33_ASAP7_75t_L g911 ( .A(n_866), .Y(n_911) );
BUFx2_ASAP7_75t_L g912 ( .A(n_855), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_853), .B(n_835), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_894), .B(n_835), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_905), .B(n_835), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_863), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_861), .B(n_835), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_853), .B(n_840), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_870), .B(n_818), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_857), .B(n_836), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_863), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_869), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_857), .B(n_836), .Y(n_923) );
INVx1_ASAP7_75t_SL g924 ( .A(n_883), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_869), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_864), .B(n_831), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_899), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_867), .B(n_850), .Y(n_928) );
AOI211xp5_ASAP7_75t_L g929 ( .A1(n_851), .A2(n_873), .B(n_893), .C(n_884), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_899), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_850), .Y(n_931) );
INVx3_ASAP7_75t_L g932 ( .A(n_880), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_883), .B(n_868), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_852), .Y(n_934) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_896), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_868), .B(n_872), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_875), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_877), .B(n_885), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_881), .B(n_886), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_874), .B(n_888), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_900), .B(n_898), .Y(n_941) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_858), .B(n_887), .C(n_865), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_849), .B(n_855), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_848), .Y(n_944) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_896), .Y(n_945) );
OR2x2_ASAP7_75t_L g946 ( .A(n_895), .B(n_906), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_848), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_895), .B(n_906), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_859), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_889), .B(n_891), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_875), .Y(n_951) );
BUFx2_ASAP7_75t_L g952 ( .A(n_880), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_879), .B(n_901), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_879), .B(n_901), .Y(n_954) );
OAI31xp33_ASAP7_75t_L g955 ( .A1(n_849), .A2(n_878), .A3(n_892), .B(n_860), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_862), .B(n_871), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_862), .B(n_907), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_859), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_876), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_908), .B(n_862), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_907), .B(n_854), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_924), .B(n_907), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_916), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_916), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_922), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_921), .Y(n_966) );
INVx1_ASAP7_75t_SL g967 ( .A(n_933), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_921), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_946), .B(n_903), .Y(n_969) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_935), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_953), .B(n_854), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_925), .Y(n_972) );
INVx3_ASAP7_75t_L g973 ( .A(n_932), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_925), .Y(n_974) );
INVx1_ASAP7_75t_SL g975 ( .A(n_933), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_953), .B(n_882), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_922), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_927), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_931), .B(n_887), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_931), .B(n_856), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_927), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_946), .B(n_902), .Y(n_982) );
NAND2x1_ASAP7_75t_L g983 ( .A(n_932), .B(n_902), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_936), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_930), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_937), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_930), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_954), .B(n_882), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_952), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_944), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_940), .B(n_904), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_940), .B(n_904), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_937), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_936), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_944), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_951), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_947), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_951), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_991), .B(n_956), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_969), .Y(n_1000) );
AOI222xp33_ASAP7_75t_SL g1001 ( .A1(n_967), .A2(n_911), .B1(n_934), .B2(n_912), .C1(n_929), .C2(n_932), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_975), .B(n_950), .Y(n_1002) );
AOI21xp33_ASAP7_75t_SL g1003 ( .A1(n_989), .A2(n_955), .B(n_943), .Y(n_1003) );
INVxp67_ASAP7_75t_L g1004 ( .A(n_970), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_963), .Y(n_1005) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_984), .B(n_939), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_994), .B(n_918), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_983), .A2(n_942), .B1(n_910), .B2(n_919), .Y(n_1008) );
INVx2_ASAP7_75t_L g1009 ( .A(n_965), .Y(n_1009) );
OAI21xp33_ASAP7_75t_L g1010 ( .A1(n_979), .A2(n_962), .B(n_991), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_992), .B(n_928), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_983), .A2(n_955), .B(n_910), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_973), .A2(n_910), .B1(n_982), .B2(n_960), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_982), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_992), .B(n_956), .Y(n_1015) );
A2O1A1Ixp33_ASAP7_75t_L g1016 ( .A1(n_973), .A2(n_910), .B(n_934), .C(n_897), .Y(n_1016) );
AOI21xp33_ASAP7_75t_L g1017 ( .A1(n_973), .A2(n_914), .B(n_948), .Y(n_1017) );
OAI31xp33_ASAP7_75t_L g1018 ( .A1(n_976), .A2(n_923), .A3(n_920), .B(n_957), .Y(n_1018) );
OAI221xp5_ASAP7_75t_L g1019 ( .A1(n_980), .A2(n_938), .B1(n_914), .B2(n_917), .C(n_915), .Y(n_1019) );
AOI211xp5_ASAP7_75t_SL g1020 ( .A1(n_1008), .A2(n_923), .B(n_920), .C(n_913), .Y(n_1020) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_1002), .Y(n_1021) );
NAND2x1_ASAP7_75t_L g1022 ( .A(n_1012), .B(n_965), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1005), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_1009), .Y(n_1024) );
XNOR2x1_ASAP7_75t_L g1025 ( .A(n_1014), .B(n_988), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1000), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1007), .Y(n_1027) );
NAND2xp5_ASAP7_75t_SL g1028 ( .A(n_1008), .B(n_998), .Y(n_1028) );
AOI322xp5_ASAP7_75t_L g1029 ( .A1(n_1021), .A2(n_1006), .A3(n_1011), .B1(n_1010), .B2(n_999), .C1(n_1015), .C2(n_1004), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_1027), .B(n_1006), .Y(n_1030) );
AOI32xp33_ASAP7_75t_L g1031 ( .A1(n_1020), .A2(n_1013), .A3(n_1001), .B1(n_1003), .B2(n_971), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1023), .Y(n_1032) );
AOI21xp33_ASAP7_75t_L g1033 ( .A1(n_1022), .A2(n_1018), .B(n_1019), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1025), .B(n_1017), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_1028), .A2(n_945), .B1(n_1016), .B2(n_941), .Y(n_1035) );
NOR5xp2_ASAP7_75t_L g1036 ( .A(n_1026), .B(n_997), .C(n_990), .D(n_995), .E(n_977), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1032), .Y(n_1037) );
OAI321xp33_ASAP7_75t_L g1038 ( .A1(n_1031), .A2(n_961), .A3(n_1024), .B1(n_915), .B2(n_981), .C(n_964), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1029), .B(n_1024), .Y(n_1039) );
NOR2x1_ASAP7_75t_L g1040 ( .A(n_1035), .B(n_990), .Y(n_1040) );
AOI322xp5_ASAP7_75t_L g1041 ( .A1(n_1034), .A2(n_926), .A3(n_968), .B1(n_985), .B2(n_978), .C1(n_966), .C2(n_987), .Y(n_1041) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_1033), .B(n_978), .C(n_968), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_1037), .B(n_1030), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_1039), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_1038), .B(n_1042), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_1040), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1041), .B(n_981), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_1044), .A2(n_974), .B1(n_972), .B2(n_997), .Y(n_1048) );
NOR3xp33_ASAP7_75t_L g1049 ( .A(n_1045), .B(n_972), .C(n_974), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1043), .Y(n_1050) );
NAND4xp75_ASAP7_75t_L g1051 ( .A(n_1050), .B(n_1047), .C(n_1046), .D(n_1036), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1048), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_1051), .A2(n_1049), .B1(n_890), .B2(n_996), .Y(n_1053) );
OAI22x1_ASAP7_75t_L g1054 ( .A1(n_1052), .A2(n_998), .B1(n_996), .B2(n_993), .Y(n_1054) );
AOI22x1_ASAP7_75t_L g1055 ( .A1(n_1054), .A2(n_986), .B1(n_958), .B2(n_949), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1053), .Y(n_1056) );
OAI22x1_ASAP7_75t_L g1057 ( .A1(n_1056), .A2(n_958), .B1(n_949), .B2(n_947), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1057), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_1058), .A2(n_1055), .B1(n_890), .B2(n_959), .Y(n_1059) );
endmodule