module fake_jpeg_20097_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_36),
.B1(n_26),
.B2(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_23),
.B1(n_27),
.B2(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_17),
.B1(n_19),
.B2(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_53),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_43),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_64),
.B1(n_36),
.B2(n_43),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_39),
.B1(n_19),
.B2(n_21),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_20),
.B1(n_27),
.B2(n_14),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_13),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_16),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_36),
.B1(n_20),
.B2(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_25),
.B1(n_16),
.B2(n_53),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_48),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_63),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_47),
.B1(n_48),
.B2(n_45),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_71),
.B1(n_25),
.B2(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR4xp25_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_92),
.C(n_75),
.D(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_66),
.C(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.C(n_83),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_103),
.B1(n_80),
.B2(n_93),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_77),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_88),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_79),
.B(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_52),
.C(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

AO221x1_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_52),
.B1(n_101),
.B2(n_51),
.C(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_93),
.B1(n_85),
.B2(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_84),
.B1(n_51),
.B2(n_40),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_106),
.C(n_112),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_105),
.B(n_111),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_124),
.B(n_52),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.C(n_118),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_113),
.B1(n_117),
.B2(n_116),
.Y(n_123)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_127),
.B(n_121),
.Y(n_130)
);

AOI31xp67_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_9),
.A3(n_10),
.B(n_5),
.Y(n_126)
);

AOI31xp67_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_128),
.A3(n_6),
.B(n_3),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_8),
.B(n_12),
.C(n_6),
.D(n_7),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_123),
.A3(n_121),
.B1(n_124),
.B2(n_59),
.C1(n_60),
.C2(n_12),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.C(n_46),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_46),
.C(n_2),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_132),
.B(n_2),
.Y(n_135)
);


endmodule