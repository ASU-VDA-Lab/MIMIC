module real_jpeg_23652_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_0),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_2),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_2),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_84),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_2),
.B(n_52),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_2),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_84),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_3),
.B(n_52),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_3),
.B(n_49),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_3),
.B(n_40),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_3),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_3),
.B(n_109),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_7),
.B(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_84),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_7),
.B(n_40),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_7),
.B(n_29),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_7),
.B(n_25),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_7),
.B(n_109),
.Y(n_304)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_40),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_9),
.B(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_9),
.B(n_84),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_25),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_103),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_10),
.B(n_84),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_10),
.B(n_52),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_11),
.B(n_49),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_11),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_11),
.B(n_84),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_12),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_84),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_12),
.B(n_52),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_12),
.B(n_49),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_12),
.B(n_40),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_12),
.B(n_29),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_15),
.B(n_243),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_15),
.B(n_52),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_16),
.B(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_16),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_16),
.B(n_52),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_16),
.B(n_84),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_16),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_29),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_16),
.B(n_25),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_16),
.B(n_109),
.Y(n_287)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_17),
.Y(n_192)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_17),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_54),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_118),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_63),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.CI(n_32),
.CON(n_23),
.SN(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_26),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_26),
.B(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.C(n_41),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_40),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_43),
.B(n_54),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.C(n_51),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_45),
.B(n_48),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_58),
.C(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_46),
.A2(n_51),
.B1(n_59),
.B2(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_48),
.B(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_51),
.B(n_79),
.C(n_82),
.Y(n_116)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_111),
.C(n_117),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_75),
.A2(n_76),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_95),
.C(n_97),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_77),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.C(n_91),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_78),
.B(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_100),
.C(n_105),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_82),
.A2(n_86),
.B1(n_100),
.B2(n_101),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_83),
.B(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_87),
.B(n_91),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_88),
.B(n_89),
.CI(n_90),
.CON(n_330),
.SN(n_330)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_91),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.CI(n_94),
.CON(n_91),
.SN(n_91)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_367),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_95),
.Y(n_367)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.C(n_110),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_99),
.B(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_100),
.A2(n_101),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_100),
.B(n_308),
.C(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_105),
.B(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_340),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_110),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_110),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_110),
.B(n_336),
.C(n_339),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_111),
.B(n_117),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_112),
.A2(n_113),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_115),
.B(n_116),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_368),
.C(n_369),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_356),
.C(n_357),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_344),
.C(n_345),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_320),
.C(n_321),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_289),
.C(n_290),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_254),
.C(n_255),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_222),
.C(n_223),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_197),
.C(n_198),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_158),
.C(n_169),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_137),
.C(n_142),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_132),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_151),
.C(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_157),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_168),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_193),
.C(n_194),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.C(n_183),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_188),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_211),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_212),
.C(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_205),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_207),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.CI(n_210),
.CON(n_207),
.SN(n_207)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_238),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_227),
.C(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_234),
.C(n_237),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_229),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.CI(n_232),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_246),
.C(n_252),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_246),
.B1(n_252),
.B2(n_253),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_241),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_244),
.B(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_244),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_245),
.B(n_279),
.C(n_280),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_275),
.B2(n_288),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_276),
.C(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_260),
.C(n_268),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_268),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_264),
.C(n_267),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_316),
.C(n_317),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.CI(n_287),
.CON(n_281),
.SN(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_318),
.B2(n_319),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_310),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_310),
.C(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_301),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_302),
.C(n_303),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_297),
.C(n_299),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_309),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.C(n_343),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_343),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_330),
.Y(n_374)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_331),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_342),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_339),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_355),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_349),
.C(n_355),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_352),
.C(n_353),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_360),
.C(n_365),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_364),
.B2(n_365),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);


endmodule