module fake_ibex_755_n_3181 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3181);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3181;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_1782;
wire n_963;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_2723;
wire n_1616;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_822;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1599;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_3070;
wire n_2711;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_634;
wire n_991;
wire n_1349;
wire n_1223;
wire n_1331;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1860;
wire n_1491;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1839;
wire n_1617;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_1622;
wire n_897;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_3102;
wire n_2872;
wire n_2790;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_980;
wire n_849;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_1379;
wire n_759;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_635;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2303;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2961;
wire n_2996;
wire n_2704;
wire n_2770;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_436),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_146),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_222),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_297),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_466),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_232),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_508),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_175),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_8),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_31),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_297),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_600),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_77),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_249),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_570),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_535),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_226),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_270),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_346),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_279),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_203),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_281),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_91),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_543),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_413),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_376),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_597),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_348),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_52),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_88),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_152),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_407),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_72),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_229),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_334),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_463),
.Y(n_670)
);

BUFx8_ASAP7_75t_SL g671 ( 
.A(n_540),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_14),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_605),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_357),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_551),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_591),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_344),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_56),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_414),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_448),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_273),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_20),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_318),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_448),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_0),
.Y(n_685)
);

BUFx2_ASAP7_75t_R g686 ( 
.A(n_174),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_596),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_193),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_373),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_246),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_616),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_98),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_345),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_245),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_330),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_253),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_465),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_111),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_173),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_633),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_488),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_151),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_145),
.Y(n_703)
);

BUFx8_ASAP7_75t_SL g704 ( 
.A(n_52),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_341),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_117),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_432),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_366),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_168),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_304),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_100),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_617),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_569),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_25),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_112),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_129),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_25),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_240),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_517),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_202),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_135),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_58),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_53),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_375),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_629),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_265),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_100),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_579),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_598),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_275),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_58),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_236),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_91),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_441),
.Y(n_735)
);

BUFx2_ASAP7_75t_SL g736 ( 
.A(n_450),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_138),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_334),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_168),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_343),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_180),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_478),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_263),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_250),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_376),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_264),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_391),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_108),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_309),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_328),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_61),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_114),
.Y(n_752)
);

INVxp33_ASAP7_75t_R g753 ( 
.A(n_95),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_13),
.Y(n_754)
);

BUFx8_ASAP7_75t_SL g755 ( 
.A(n_187),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_14),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_343),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_556),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_239),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_240),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_565),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_531),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_521),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_614),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_125),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_95),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_357),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_373),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_470),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_253),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_64),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_190),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_541),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_50),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_138),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_564),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_571),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_289),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_555),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_536),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_479),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_537),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_593),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_403),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_458),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_532),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_411),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_207),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_20),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_504),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_552),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_74),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_503),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_375),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_532),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_476),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_0),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_322),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_50),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_493),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_324),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_27),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_492),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_458),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_442),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_134),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_405),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_320),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_426),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_257),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_142),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_498),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_90),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_242),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_484),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_355),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_490),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_175),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_567),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_189),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_254),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_285),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_248),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_576),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_302),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_54),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_160),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_182),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_603),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_624),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_444),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_324),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_189),
.Y(n_833)
);

CKINVDCx14_ASAP7_75t_R g834 ( 
.A(n_549),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_520),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_68),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_243),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_302),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_408),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_255),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_426),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_526),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_286),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_319),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_583),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_585),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_92),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_608),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_421),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_517),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_613),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_145),
.Y(n_852)
);

BUFx5_ASAP7_75t_L g853 ( 
.A(n_15),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_358),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_500),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_440),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_498),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_1),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_1),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_184),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_560),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_94),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_285),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_30),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_73),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_619),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_114),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_179),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_533),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_54),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_9),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_374),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_40),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_559),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_580),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_98),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_67),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_171),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_172),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_219),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_252),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_421),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_148),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_420),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_178),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_404),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_383),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_590),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_611),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_123),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_428),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_459),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_267),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_500),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_496),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_508),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_466),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_339),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_117),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_310),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_320),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_394),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_126),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_162),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_526),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_37),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_312),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_398),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_439),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_122),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_76),
.Y(n_911)
);

CKINVDCx16_ASAP7_75t_R g912 ( 
.A(n_402),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_2),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_23),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_475),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_400),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_602),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_630),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_23),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_363),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_86),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_340),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_7),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_293),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_519),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_247),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_522),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_209),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_60),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_103),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_42),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_38),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_273),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_365),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_65),
.Y(n_935)
);

BUFx2_ASAP7_75t_SL g936 ( 
.A(n_103),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_509),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_41),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_490),
.Y(n_939)
);

BUFx10_ASAP7_75t_L g940 ( 
.A(n_574),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_325),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_355),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_33),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_210),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_546),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_170),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_311),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_28),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_242),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_32),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_153),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_537),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_394),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_326),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_214),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_44),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_26),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_184),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_464),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_314),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_16),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_577),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_519),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_197),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_88),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_57),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_444),
.Y(n_967)
);

BUFx10_ASAP7_75t_L g968 ( 
.A(n_19),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_587),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_13),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_154),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_190),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_22),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_393),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_288),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_516),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_366),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_514),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_256),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_148),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_68),
.Y(n_981)
);

BUFx2_ASAP7_75t_R g982 ( 
.A(n_612),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_509),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_329),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_222),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_83),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_499),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_563),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_258),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_278),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_575),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_43),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_4),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_211),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_572),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_56),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_384),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_281),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_206),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_471),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_35),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_131),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_248),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_329),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_483),
.Y(n_1005)
);

CKINVDCx16_ASAP7_75t_R g1006 ( 
.A(n_251),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_327),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_365),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_221),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_16),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_335),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_172),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_232),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_419),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_44),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_695),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_912),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_695),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_713),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_695),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_1006),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_645),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_740),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_691),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_982),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_834),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_752),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_635),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_641),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_643),
.Y(n_1030)
);

CKINVDCx16_ASAP7_75t_R g1031 ( 
.A(n_731),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_752),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_671),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_704),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_646),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_825),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_755),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_648),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_648),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_740),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_898),
.B(n_2),
.Y(n_1041)
);

INVxp33_ASAP7_75t_SL g1042 ( 
.A(n_634),
.Y(n_1042)
);

INVxp33_ASAP7_75t_SL g1043 ( 
.A(n_634),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_820),
.B(n_4),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_986),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_661),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_673),
.B(n_3),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_661),
.Y(n_1048)
);

INVxp33_ASAP7_75t_SL g1049 ( 
.A(n_637),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_986),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1003),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_647),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_700),
.B(n_3),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_660),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1003),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_676),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_719),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_719),
.Y(n_1058)
);

NOR2xp67_ASAP7_75t_L g1059 ( 
.A(n_787),
.B(n_5),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_728),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_676),
.Y(n_1061)
);

CKINVDCx14_ASAP7_75t_R g1062 ( 
.A(n_940),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_655),
.A2(n_554),
.B(n_553),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_687),
.Y(n_1064)
);

INVxp33_ASAP7_75t_SL g1065 ( 
.A(n_637),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_728),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_763),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_740),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_687),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_962),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_740),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_763),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_962),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_638),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_665),
.Y(n_1075)
);

INVxp33_ASAP7_75t_SL g1076 ( 
.A(n_638),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_903),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_678),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_988),
.Y(n_1079)
);

INVxp67_ASAP7_75t_SL g1080 ( 
.A(n_989),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_731),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_731),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_706),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_707),
.Y(n_1084)
);

CKINVDCx16_ASAP7_75t_R g1085 ( 
.A(n_742),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_751),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_989),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_701),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_701),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_705),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_988),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_642),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_705),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_708),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_708),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_734),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_734),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_642),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_748),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_785),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_649),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_748),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_756),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_792),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_756),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_766),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_766),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_718),
.B(n_730),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_742),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_774),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_740),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_649),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_774),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_794),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_651),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_651),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_652),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_782),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_803),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_740),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_758),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_807),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_816),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_653),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_790),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_790),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_809),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_809),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_653),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_740),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_811),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_811),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_892),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_654),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_892),
.B(n_6),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_654),
.Y(n_1136)
);

CKINVDCx16_ASAP7_75t_R g1137 ( 
.A(n_742),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_835),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_909),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_909),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_656),
.B(n_1010),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_928),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_928),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_842),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_996),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_656),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_1121),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1023),
.B(n_1040),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1040),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1027),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1068),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1032),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1063),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1068),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1036),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1066),
.B(n_930),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1062),
.B(n_930),
.Y(n_1157)
);

AND2x6_ASAP7_75t_L g1158 ( 
.A(n_1016),
.B(n_758),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1071),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1121),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1042),
.A2(n_658),
.B1(n_659),
.B2(n_657),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_L g1163 ( 
.A(n_1038),
.B(n_740),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1042),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1050),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1136),
.B(n_930),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1051),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1018),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1063),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1055),
.B(n_1022),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1071),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1043),
.A2(n_658),
.B1(n_659),
.B2(n_657),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_1132),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1020),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1057),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1111),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1058),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1120),
.Y(n_1178)
);

AND3x2_ASAP7_75t_L g1179 ( 
.A(n_1074),
.B(n_686),
.C(n_753),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1060),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1067),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1120),
.Y(n_1182)
);

INVxp33_ASAP7_75t_L g1183 ( 
.A(n_1112),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1072),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1080),
.B(n_1141),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1130),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1130),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1093),
.B(n_996),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1132),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1043),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1077),
.Y(n_1191)
);

BUFx8_ASAP7_75t_L g1192 ( 
.A(n_1049),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1132),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1087),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1107),
.B(n_955),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1118),
.B(n_955),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1081),
.B(n_655),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1128),
.B(n_663),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1088),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1089),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1090),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1094),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1095),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1096),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1097),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1041),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_1031),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1108),
.B(n_675),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1053),
.A2(n_888),
.B(n_675),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1102),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1103),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1115),
.B(n_663),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1105),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1106),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1049),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1065),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1110),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1113),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1125),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1126),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1127),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1131),
.Y(n_1223)
);

AND2x2_ASAP7_75t_SL g1224 ( 
.A(n_1082),
.B(n_1002),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1039),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1133),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1139),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_1065),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1140),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1142),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1143),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1145),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1044),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1085),
.B(n_968),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1109),
.B(n_968),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1047),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1046),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1076),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1048),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1135),
.B(n_1002),
.Y(n_1240)
);

XNOR2xp5_ASAP7_75t_L g1241 ( 
.A(n_1017),
.B(n_858),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1056),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1137),
.B(n_955),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1061),
.B(n_888),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1076),
.B(n_664),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1064),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1069),
.B(n_669),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1059),
.B(n_636),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1070),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1073),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1079),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1091),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1092),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1098),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1101),
.A2(n_819),
.B(n_783),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1116),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1124),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1129),
.B(n_824),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1134),
.Y(n_1260)
);

BUFx8_ASAP7_75t_L g1261 ( 
.A(n_1026),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1024),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1026),
.B(n_968),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1019),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1017),
.B(n_640),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1021),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1033),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1021),
.B(n_669),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1034),
.B(n_940),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1037),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1028),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1025),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1028),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1029),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1029),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1030),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1030),
.B(n_650),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1035),
.B(n_681),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1035),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1052),
.B(n_667),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1052),
.Y(n_1282)
);

AND2x2_ASAP7_75t_SL g1283 ( 
.A(n_1054),
.B(n_639),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1075),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1075),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1078),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1078),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1083),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1083),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1084),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1084),
.B(n_668),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1144),
.B(n_940),
.Y(n_1292)
);

INVxp33_ASAP7_75t_SL g1293 ( 
.A(n_1086),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1086),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1100),
.B(n_681),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1100),
.B(n_682),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1104),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1104),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1114),
.B(n_682),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1114),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1144),
.B(n_991),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1119),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1119),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1122),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1122),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1123),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1123),
.A2(n_881),
.B1(n_895),
.B2(n_879),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1138),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1138),
.B(n_991),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1027),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1063),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1063),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1022),
.B(n_829),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1023),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_L g1315 ( 
.A(n_1141),
.B(n_830),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1027),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1136),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1027),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1023),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1023),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1027),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1027),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1066),
.B(n_991),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1027),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1023),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1136),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1023),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1027),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1066),
.B(n_683),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1023),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1023),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1063),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1027),
.B(n_670),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1023),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1066),
.B(n_684),
.Y(n_1335)
);

XOR2xp5_ASAP7_75t_L g1336 ( 
.A(n_1028),
.B(n_932),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1023),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1063),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1023),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1023),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1044),
.B(n_736),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1066),
.B(n_853),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1136),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1063),
.A2(n_861),
.B(n_845),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1136),
.Y(n_1345)
);

CKINVDCx8_ASAP7_75t_R g1346 ( 
.A(n_1025),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1023),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1023),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1027),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1023),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1063),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1190),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1326),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1311),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1326),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1173),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1207),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1311),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1311),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1343),
.B(n_711),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1173),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1173),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1224),
.A2(n_693),
.B1(n_694),
.B2(n_688),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1193),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1162),
.B(n_693),
.C(n_688),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1185),
.B(n_918),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1343),
.B(n_694),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1233),
.A2(n_867),
.B1(n_853),
.B2(n_674),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1193),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1345),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1193),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1201),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1312),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1345),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1207),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.B(n_699),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1201),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1233),
.B(n_712),
.Y(n_1378)
);

BUFx8_ASAP7_75t_SL g1379 ( 
.A(n_1272),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1295),
.B(n_699),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1168),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1312),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1236),
.B(n_969),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1161),
.Y(n_1384)
);

AND2x2_ASAP7_75t_SL g1385 ( 
.A(n_1283),
.B(n_639),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1236),
.B(n_995),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1210),
.A2(n_867),
.B1(n_853),
.B2(n_672),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1168),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1332),
.B(n_875),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1341),
.B(n_677),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1161),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1332),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1201),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1332),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1338),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1201),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1150),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1198),
.B(n_726),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1206),
.B(n_729),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1338),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1218),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1192),
.Y(n_1402)
);

INVxp33_ASAP7_75t_L g1403 ( 
.A(n_1216),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1153),
.B(n_761),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1170),
.B(n_764),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1153),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1218),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1153),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1153),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1153),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1192),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1210),
.A2(n_1255),
.B1(n_1229),
.B2(n_1200),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1169),
.B(n_776),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1169),
.Y(n_1414)
);

AND2x2_ASAP7_75t_SL g1415 ( 
.A(n_1283),
.B(n_639),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1183),
.B(n_711),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1207),
.B(n_680),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1152),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1155),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1207),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1169),
.B(n_777),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1351),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1218),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1207),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1157),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1217),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1157),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1351),
.B(n_779),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1183),
.B(n_814),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1351),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1159),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1165),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1253),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1351),
.B(n_791),
.Y(n_1434)
);

NAND2xp33_ASAP7_75t_SL g1435 ( 
.A(n_1164),
.B(n_702),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1351),
.B(n_846),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1158),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1147),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1167),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1310),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_R g1441 ( 
.A(n_1252),
.B(n_702),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1170),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1344),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1341),
.A2(n_709),
.B1(n_813),
.B2(n_703),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1316),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1218),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1170),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1147),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1333),
.B(n_848),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1228),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1149),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1195),
.B(n_851),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_L g1453 ( 
.A(n_1158),
.B(n_853),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1318),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1180),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1182),
.B(n_866),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1182),
.B(n_874),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1228),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1219),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1182),
.B(n_889),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1151),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1210),
.A2(n_867),
.B1(n_853),
.B2(n_685),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1333),
.B(n_917),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1238),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1234),
.B(n_931),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1341),
.B(n_689),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1151),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1333),
.B(n_690),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1245),
.B(n_709),
.C(n_703),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1225),
.B(n_813),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1321),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1154),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1228),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1341),
.B(n_936),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1234),
.B(n_814),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1180),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1219),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1255),
.A2(n_867),
.B1(n_853),
.B2(n_692),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1322),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1253),
.B(n_696),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1324),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1147),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1219),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1225),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1328),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1160),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1195),
.B(n_853),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1262),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1244),
.B(n_698),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1182),
.B(n_853),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1219),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1172),
.B(n_927),
.C(n_823),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1244),
.B(n_710),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1249),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1235),
.B(n_937),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_L g1496 ( 
.A(n_1158),
.B(n_867),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1158),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1171),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1262),
.B(n_714),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1315),
.B(n_717),
.Y(n_1500)
);

OR2x2_ASAP7_75t_SL g1501 ( 
.A(n_1287),
.B(n_951),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1158),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1226),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1186),
.B(n_867),
.Y(n_1504)
);

OR2x2_ASAP7_75t_SL g1505 ( 
.A(n_1287),
.B(n_953),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1171),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1226),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1296),
.B(n_927),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1258),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_L g1510 ( 
.A(n_1271),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1158),
.Y(n_1511)
);

BUFx2_ASAP7_75t_SL g1512 ( 
.A(n_1243),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1349),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1255),
.A2(n_867),
.B1(n_723),
.B2(n_727),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1342),
.B(n_721),
.Y(n_1515)
);

AND3x2_ASAP7_75t_L g1516 ( 
.A(n_1279),
.B(n_1013),
.C(n_1014),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1229),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1243),
.B(n_934),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1261),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1258),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1186),
.B(n_867),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1196),
.B(n_1342),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1229),
.A2(n_735),
.B1(n_738),
.B2(n_733),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1186),
.B(n_639),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1209),
.Y(n_1525)
);

INVx4_ASAP7_75t_L g1526 ( 
.A(n_1260),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1226),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_SL g1528 ( 
.A(n_1252),
.B(n_929),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1260),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1176),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1211),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1176),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1221),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1260),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1174),
.A2(n_1188),
.B1(n_1313),
.B2(n_1202),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1178),
.Y(n_1536)
);

BUFx8_ASAP7_75t_SL g1537 ( 
.A(n_1272),
.Y(n_1537)
);

NAND2xp33_ASAP7_75t_L g1538 ( 
.A(n_1249),
.B(n_639),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_L g1539 ( 
.A(n_1249),
.B(n_720),
.Y(n_1539)
);

OAI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1293),
.A2(n_934),
.B1(n_937),
.B2(n_931),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1222),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1178),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1187),
.B(n_720),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1187),
.B(n_720),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1223),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1227),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1314),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1314),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1254),
.B(n_743),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1319),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1232),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1199),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1199),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1187),
.B(n_1319),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1257),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1156),
.B(n_946),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1249),
.B(n_720),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1188),
.B(n_939),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1320),
.Y(n_1559)
);

NOR2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1275),
.B(n_939),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1202),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1261),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1271),
.B(n_750),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1325),
.B(n_720),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1156),
.B(n_941),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1325),
.Y(n_1566)
);

AND2x6_ASAP7_75t_L g1567 ( 
.A(n_1249),
.B(n_854),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1327),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1327),
.B(n_854),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1299),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1254),
.B(n_771),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1197),
.B(n_775),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1203),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1330),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1203),
.Y(n_1575)
);

BUFx10_ASAP7_75t_L g1576 ( 
.A(n_1271),
.Y(n_1576)
);

AO22x2_ASAP7_75t_L g1577 ( 
.A1(n_1248),
.A2(n_784),
.B1(n_786),
.B2(n_778),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1204),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1204),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1205),
.Y(n_1580)
);

XNOR2xp5_ASAP7_75t_L g1581 ( 
.A(n_1336),
.B(n_998),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1330),
.B(n_854),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1205),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1197),
.B(n_793),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1212),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1214),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1214),
.Y(n_1587)
);

AND2x6_ASAP7_75t_L g1588 ( 
.A(n_1237),
.B(n_854),
.Y(n_1588)
);

INVx5_ASAP7_75t_L g1589 ( 
.A(n_1215),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1331),
.Y(n_1590)
);

AND2x6_ASAP7_75t_L g1591 ( 
.A(n_1237),
.B(n_854),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1331),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1313),
.A2(n_796),
.B1(n_798),
.B2(n_795),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1334),
.B(n_880),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1215),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1189),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1166),
.B(n_943),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1336),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1269),
.Y(n_1599)
);

INVxp33_ASAP7_75t_L g1600 ( 
.A(n_1166),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1334),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1220),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1220),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1337),
.B(n_880),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1213),
.B(n_942),
.C(n_941),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1323),
.B(n_942),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1323),
.Y(n_1607)
);

BUFx10_ASAP7_75t_L g1608 ( 
.A(n_1271),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1337),
.Y(n_1609)
);

AND2x6_ASAP7_75t_L g1610 ( 
.A(n_1239),
.B(n_880),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1576),
.Y(n_1611)
);

AND2x4_ASAP7_75t_SL g1612 ( 
.A(n_1484),
.B(n_1264),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1535),
.B(n_1224),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1397),
.Y(n_1615)
);

AO221x1_ASAP7_75t_L g1616 ( 
.A1(n_1353),
.A2(n_1307),
.B1(n_1285),
.B2(n_1302),
.C(n_1305),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1484),
.B(n_1433),
.Y(n_1617)
);

BUFx5_ASAP7_75t_L g1618 ( 
.A(n_1567),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1596),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1418),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_R g1621 ( 
.A(n_1402),
.B(n_1261),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1359),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1535),
.B(n_1329),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1522),
.B(n_1239),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1442),
.B(n_1246),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1470),
.B(n_1260),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1419),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_R g1628 ( 
.A(n_1473),
.B(n_1346),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1359),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1528),
.B(n_1247),
.C(n_1264),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1455),
.B(n_1250),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1424),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1596),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1431),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1455),
.B(n_1250),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1432),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1439),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1600),
.B(n_1256),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1355),
.B(n_1241),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1440),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1476),
.B(n_1242),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1607),
.A2(n_1266),
.B1(n_1259),
.B2(n_1251),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1596),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1259),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1572),
.A2(n_1208),
.B(n_1163),
.C(n_1230),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1476),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1558),
.B(n_1248),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1390),
.B(n_1571),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1390),
.B(n_1248),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1502),
.B(n_1242),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1385),
.A2(n_1175),
.B1(n_1181),
.B2(n_1177),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1571),
.B(n_1184),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1385),
.A2(n_1415),
.B1(n_1515),
.B2(n_1383),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1445),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1417),
.B(n_1242),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1442),
.B(n_1263),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1454),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1370),
.B(n_1292),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1447),
.B(n_1292),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1412),
.B(n_1339),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1571),
.B(n_1447),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1426),
.Y(n_1663)
);

AND2x6_ASAP7_75t_SL g1664 ( 
.A(n_1598),
.B(n_1274),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1356),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1488),
.B(n_1301),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1465),
.A2(n_1266),
.B1(n_1263),
.B2(n_1309),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1480),
.A2(n_1231),
.B1(n_1230),
.B2(n_945),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1471),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1361),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1479),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1415),
.A2(n_1194),
.B1(n_1191),
.B2(n_1231),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1362),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1466),
.B(n_1265),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1475),
.A2(n_1266),
.B1(n_1309),
.B2(n_1301),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1379),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1481),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1474),
.B(n_1466),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1364),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1485),
.Y(n_1680)
);

INVx8_ASAP7_75t_L g1681 ( 
.A(n_1474),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1452),
.B(n_1380),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1416),
.B(n_1278),
.Y(n_1683)
);

INVx8_ASAP7_75t_L g1684 ( 
.A(n_1474),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1508),
.B(n_1270),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1367),
.B(n_1241),
.Y(n_1686)
);

BUFx8_ASAP7_75t_L g1687 ( 
.A(n_1520),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1417),
.B(n_1268),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1606),
.B(n_1163),
.Y(n_1689)
);

BUFx8_ASAP7_75t_L g1690 ( 
.A(n_1495),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1374),
.B(n_1275),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1513),
.B(n_1549),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1589),
.B(n_1278),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1549),
.B(n_1240),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1515),
.A2(n_1189),
.B1(n_1240),
.B2(n_1278),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1429),
.B(n_1240),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1589),
.B(n_1281),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1515),
.B(n_1281),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1480),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1512),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1556),
.B(n_1267),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1499),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1499),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1489),
.B(n_1281),
.Y(n_1704)
);

BUFx2_ASAP7_75t_R g1705 ( 
.A(n_1379),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1360),
.B(n_1291),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1369),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1589),
.B(n_1291),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1565),
.B(n_1267),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1425),
.B(n_1291),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1489),
.B(n_1493),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1493),
.B(n_943),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1359),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1371),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1441),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1383),
.A2(n_806),
.B1(n_808),
.B2(n_805),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1525),
.B(n_945),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1531),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1597),
.B(n_1276),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1533),
.B(n_947),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1541),
.Y(n_1721)
);

BUFx8_ASAP7_75t_L g1722 ( 
.A(n_1518),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1589),
.B(n_1285),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1359),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1424),
.B(n_1285),
.Y(n_1725)
);

AO221x1_ASAP7_75t_L g1726 ( 
.A1(n_1577),
.A2(n_1285),
.B1(n_1302),
.B2(n_1305),
.C(n_1287),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1437),
.B(n_1497),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1403),
.B(n_1273),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1545),
.B(n_1546),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1551),
.B(n_947),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1469),
.B(n_1276),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1552),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1468),
.B(n_949),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1468),
.B(n_949),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1403),
.A2(n_1290),
.B1(n_1294),
.B2(n_1289),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1487),
.A2(n_1290),
.B1(n_1294),
.B2(n_1289),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1561),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1437),
.B(n_1287),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1509),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1437),
.B(n_1302),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1500),
.B(n_950),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1500),
.B(n_950),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1386),
.B(n_1572),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1365),
.B(n_1605),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1497),
.B(n_1302),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1386),
.B(n_952),
.Y(n_1746)
);

NOR3xp33_ASAP7_75t_L g1747 ( 
.A(n_1540),
.B(n_1280),
.C(n_1277),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1584),
.B(n_952),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1449),
.B(n_1297),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1575),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1576),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1575),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1392),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1384),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1584),
.B(n_958),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1463),
.B(n_1298),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1497),
.B(n_1305),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1463),
.B(n_1298),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1553),
.A2(n_1340),
.B(n_1348),
.C(n_1347),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1580),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1378),
.B(n_1405),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1517),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1599),
.A2(n_961),
.B1(n_964),
.B2(n_958),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1563),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1580),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_L g1766 ( 
.A(n_1519),
.B(n_1300),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1411),
.B(n_1346),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1570),
.B(n_1303),
.Y(n_1768)
);

OAI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1363),
.A2(n_1306),
.B1(n_1308),
.B2(n_1304),
.C(n_1303),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1444),
.B(n_961),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1602),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1523),
.B(n_964),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1577),
.A2(n_818),
.B1(n_821),
.B2(n_810),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1352),
.A2(n_966),
.B1(n_967),
.B2(n_965),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1464),
.A2(n_966),
.B1(n_967),
.B2(n_965),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1523),
.B(n_971),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1555),
.B(n_1304),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1427),
.B(n_1492),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1602),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1441),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1497),
.B(n_1340),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1563),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1514),
.A2(n_1578),
.B1(n_1579),
.B2(n_1573),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1376),
.B(n_1306),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1384),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_SL g1786 ( 
.A(n_1563),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1608),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1514),
.A2(n_1308),
.B1(n_973),
.B2(n_974),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1581),
.B(n_1282),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1560),
.B(n_1305),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1583),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1537),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1608),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1511),
.B(n_972),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1511),
.B(n_972),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1435),
.B(n_1286),
.C(n_1284),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1451),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1585),
.A2(n_974),
.B1(n_975),
.B2(n_973),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1586),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1391),
.B(n_975),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1391),
.B(n_977),
.Y(n_1801)
);

INVxp33_ASAP7_75t_L g1802 ( 
.A(n_1537),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1357),
.B(n_977),
.Y(n_1803)
);

AND2x4_ASAP7_75t_SL g1804 ( 
.A(n_1526),
.B(n_1288),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1438),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1375),
.B(n_980),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1587),
.Y(n_1807)
);

AND2x2_ASAP7_75t_SL g1808 ( 
.A(n_1510),
.B(n_880),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1595),
.A2(n_983),
.B1(n_984),
.B2(n_981),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1562),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1398),
.B(n_981),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1593),
.A2(n_985),
.B1(n_987),
.B2(n_984),
.C(n_983),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1399),
.A2(n_987),
.B1(n_990),
.B2(n_985),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1438),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1603),
.B(n_990),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1399),
.B(n_992),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1526),
.B(n_992),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1368),
.A2(n_828),
.B1(n_831),
.B2(n_826),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1420),
.B(n_993),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1593),
.B(n_1368),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1461),
.B(n_993),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1516),
.B(n_1179),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1450),
.B(n_998),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1458),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1467),
.B(n_1000),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1472),
.B(n_1000),
.Y(n_1826)
);

NAND2xp33_ASAP7_75t_L g1827 ( 
.A(n_1567),
.B(n_1348),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1510),
.B(n_1001),
.Y(n_1828)
);

NAND2xp33_ASAP7_75t_L g1829 ( 
.A(n_1567),
.B(n_1350),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1472),
.B(n_1001),
.Y(n_1830)
);

A2O1A1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1381),
.A2(n_1350),
.B(n_1148),
.C(n_833),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1478),
.B(n_1010),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1529),
.B(n_662),
.C(n_644),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1388),
.Y(n_1834)
);

INVx8_ASAP7_75t_L g1835 ( 
.A(n_1567),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1387),
.A2(n_837),
.B(n_839),
.C(n_832),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1529),
.B(n_1011),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1478),
.A2(n_1012),
.B1(n_1011),
.B2(n_715),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1534),
.A2(n_1012),
.B1(n_843),
.B2(n_850),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1501),
.B(n_666),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1534),
.B(n_840),
.Y(n_1841)
);

A2O1A1Ixp33_ASAP7_75t_L g1842 ( 
.A1(n_1387),
.A2(n_860),
.B(n_868),
.C(n_859),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1392),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1486),
.B(n_679),
.Y(n_1844)
);

INVx8_ASAP7_75t_L g1845 ( 
.A(n_1567),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1494),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1498),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1498),
.B(n_697),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1462),
.A2(n_870),
.B1(n_882),
.B2(n_869),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1506),
.B(n_716),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_L g1851 ( 
.A(n_1453),
.B(n_724),
.C(n_722),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1530),
.B(n_725),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1532),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1536),
.B(n_1542),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1536),
.B(n_732),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1448),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1547),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1547),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1448),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1548),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1548),
.B(n_737),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1550),
.B(n_739),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1559),
.A2(n_884),
.B1(n_894),
.B2(n_893),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_L g1864 ( 
.A1(n_1389),
.A2(n_901),
.B(n_914),
.C(n_908),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1566),
.A2(n_933),
.B1(n_935),
.B2(n_916),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1496),
.A2(n_744),
.B1(n_745),
.B2(n_741),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1482),
.B(n_938),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1456),
.Y(n_1868)
);

OAI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1568),
.A2(n_788),
.B1(n_801),
.B2(n_767),
.C(n_746),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1574),
.A2(n_948),
.B1(n_954),
.B2(n_944),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1590),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_SL g1872 ( 
.A(n_1610),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1482),
.B(n_1404),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1592),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1592),
.Y(n_1875)
);

AND2x6_ASAP7_75t_SL g1876 ( 
.A(n_1505),
.B(n_957),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1456),
.A2(n_1460),
.B1(n_1457),
.B2(n_1404),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1601),
.B(n_747),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1457),
.B(n_959),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1601),
.B(n_749),
.Y(n_1880)
);

OR2x2_ASAP7_75t_SL g1881 ( 
.A(n_1443),
.B(n_960),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1609),
.B(n_754),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1609),
.B(n_757),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1460),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1413),
.A2(n_760),
.B1(n_762),
.B2(n_759),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1588),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1490),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1446),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1421),
.B(n_765),
.Y(n_1889)
);

NOR3xp33_ASAP7_75t_L g1890 ( 
.A(n_1428),
.B(n_913),
.C(n_910),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1490),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1446),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1874),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1661),
.A2(n_1408),
.B(n_1406),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1682),
.B(n_768),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1685),
.B(n_1434),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1615),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1622),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1685),
.B(n_1436),
.Y(n_1899)
);

O2A1O1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1743),
.A2(n_976),
.B(n_924),
.C(n_970),
.Y(n_1900)
);

OR2x6_ASAP7_75t_L g1901 ( 
.A(n_1681),
.B(n_1409),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1622),
.A2(n_1430),
.B(n_1422),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1888),
.A2(n_1358),
.B(n_1354),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1786),
.Y(n_1904)
);

A2O1A1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1689),
.A2(n_1624),
.B(n_1682),
.C(n_1646),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1624),
.B(n_769),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1620),
.Y(n_1907)
);

O2A1O1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1704),
.A2(n_979),
.B(n_994),
.C(n_978),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1668),
.B(n_770),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1629),
.A2(n_1382),
.B(n_1373),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1627),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1874),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1668),
.B(n_772),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1635),
.B(n_773),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1675),
.B(n_1554),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1713),
.Y(n_1916)
);

AOI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1626),
.A2(n_1400),
.B(n_1395),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1692),
.B(n_780),
.Y(n_1918)
);

INVxp67_ASAP7_75t_L g1919 ( 
.A(n_1786),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1613),
.B(n_781),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1663),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1713),
.A2(n_1394),
.B(n_1392),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1724),
.A2(n_1394),
.B(n_1409),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1724),
.B(n_1394),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1761),
.A2(n_999),
.B(n_1004),
.C(n_997),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1724),
.A2(n_1394),
.B(n_1409),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1724),
.A2(n_1410),
.B(n_1409),
.Y(n_1927)
);

AOI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1832),
.A2(n_1521),
.B(n_1504),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_SL g1929 ( 
.A(n_1705),
.B(n_1588),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1859),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1634),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1753),
.A2(n_1414),
.B(n_1410),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1753),
.A2(n_1414),
.B(n_1410),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1654),
.A2(n_1377),
.B1(n_1393),
.B2(n_1372),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1820),
.A2(n_905),
.B1(n_956),
.B2(n_880),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1663),
.B(n_789),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1623),
.B(n_797),
.Y(n_1937)
);

AO21x1_ASAP7_75t_L g1938 ( 
.A1(n_1689),
.A2(n_1569),
.B(n_1564),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1621),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1666),
.B(n_799),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1649),
.B(n_800),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1687),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1637),
.Y(n_1943)
);

OAI321xp33_ASAP7_75t_L g1944 ( 
.A1(n_1773),
.A2(n_1005),
.A3(n_1008),
.B1(n_1015),
.B2(n_1009),
.C(n_1007),
.Y(n_1944)
);

AO21x2_ASAP7_75t_L g1945 ( 
.A1(n_1726),
.A2(n_1543),
.B(n_1524),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1683),
.B(n_802),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1638),
.B(n_804),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1641),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1700),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1706),
.B(n_812),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1655),
.B(n_1658),
.Y(n_1951)
);

NOR3xp33_ASAP7_75t_L g1952 ( 
.A(n_1630),
.B(n_817),
.C(n_815),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1672),
.A2(n_1396),
.B1(n_1401),
.B2(n_1372),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1843),
.A2(n_1594),
.B(n_1582),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1669),
.B(n_822),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_SL g1956 ( 
.A(n_1676),
.B(n_1588),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1671),
.B(n_827),
.Y(n_1957)
);

NAND2x1_ASAP7_75t_L g1958 ( 
.A(n_1847),
.B(n_1396),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1677),
.B(n_836),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1680),
.B(n_838),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1646),
.A2(n_1864),
.B(n_1711),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1718),
.B(n_841),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1843),
.A2(n_1604),
.B(n_1543),
.Y(n_1963)
);

NOR2x1p5_ASAP7_75t_SL g1964 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1721),
.B(n_844),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1699),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1729),
.Y(n_1967)
);

CKINVDCx10_ASAP7_75t_R g1968 ( 
.A(n_1628),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1700),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1843),
.A2(n_1544),
.B(n_1524),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1611),
.B(n_1401),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1867),
.Y(n_1972)
);

AOI33xp33_ASAP7_75t_L g1973 ( 
.A1(n_1695),
.A2(n_1716),
.A3(n_1784),
.B1(n_1773),
.B2(n_1870),
.B3(n_1863),
.Y(n_1973)
);

O2A1O1Ixp5_ASAP7_75t_L g1974 ( 
.A1(n_1864),
.A2(n_1544),
.B(n_1423),
.C(n_1477),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1672),
.A2(n_1652),
.B1(n_1662),
.B2(n_1764),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1824),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1701),
.B(n_847),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1709),
.B(n_849),
.Y(n_1978)
);

AOI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1642),
.A2(n_1459),
.B(n_1446),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1810),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1709),
.B(n_852),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1835),
.Y(n_1982)
);

BUFx4f_ASAP7_75t_L g1983 ( 
.A(n_1681),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1703),
.B(n_855),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1719),
.B(n_856),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1835),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1860),
.A2(n_1423),
.B(n_1407),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1719),
.B(n_857),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1859),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1694),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1875),
.A2(n_1507),
.B(n_1483),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1702),
.B(n_923),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1749),
.B(n_862),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1702),
.B(n_926),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1892),
.A2(n_1527),
.B(n_1459),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1691),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1841),
.Y(n_1997)
);

O2A1O1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1869),
.A2(n_1539),
.B(n_1557),
.C(n_1538),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1667),
.B(n_863),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1797),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1782),
.B(n_864),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1756),
.B(n_865),
.Y(n_2002)
);

CKINVDCx10_ASAP7_75t_R g2003 ( 
.A(n_1628),
.Y(n_2003)
);

AOI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1651),
.A2(n_1491),
.B(n_1459),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1808),
.B(n_871),
.Y(n_2005)
);

NOR2xp67_ASAP7_75t_L g2006 ( 
.A(n_1792),
.B(n_1640),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1835),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1841),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1844),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1758),
.B(n_1645),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1759),
.A2(n_1610),
.B(n_1591),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1845),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1751),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1758),
.B(n_872),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1645),
.B(n_873),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1653),
.A2(n_1503),
.B1(n_877),
.B2(n_878),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1648),
.B(n_876),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1690),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1848),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1845),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1698),
.B(n_883),
.Y(n_2021)
);

AO21x1_ASAP7_75t_L g2022 ( 
.A1(n_1873),
.A2(n_1610),
.B(n_1591),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1850),
.B(n_885),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1659),
.A2(n_887),
.B1(n_890),
.B2(n_886),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1853),
.A2(n_896),
.B(n_891),
.Y(n_2025)
);

A2O1A1Ixp33_ASAP7_75t_L g2026 ( 
.A1(n_1731),
.A2(n_956),
.B(n_963),
.C(n_905),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1748),
.B(n_897),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1881),
.A2(n_900),
.B1(n_902),
.B2(n_899),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1696),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1831),
.A2(n_1610),
.B(n_1591),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1808),
.B(n_904),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1755),
.B(n_906),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1857),
.A2(n_911),
.B(n_907),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1858),
.A2(n_919),
.B(n_915),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1674),
.B(n_920),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1871),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1887),
.A2(n_1891),
.B(n_1619),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1614),
.A2(n_922),
.B(n_921),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1633),
.A2(n_925),
.B(n_905),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1845),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1791),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1805),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1644),
.A2(n_956),
.B(n_905),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1631),
.A2(n_1636),
.B(n_1821),
.Y(n_2044)
);

NOR2x1p5_ASAP7_75t_L g2045 ( 
.A(n_1822),
.B(n_905),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1612),
.B(n_1768),
.Y(n_2046)
);

INVx5_ASAP7_75t_L g2047 ( 
.A(n_1681),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1678),
.B(n_1739),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1854),
.Y(n_2049)
);

INVxp67_ASAP7_75t_L g2050 ( 
.A(n_1817),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1799),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1768),
.B(n_963),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1674),
.B(n_7),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1747),
.A2(n_963),
.B1(n_11),
.B2(n_8),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1678),
.B(n_10),
.Y(n_2055)
);

A2O1A1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_1744),
.A2(n_1657),
.B(n_1639),
.C(n_1836),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1650),
.B(n_10),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1809),
.B(n_11),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1825),
.A2(n_558),
.B(n_557),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1809),
.B(n_12),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1826),
.A2(n_562),
.B(n_561),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_L g2062 ( 
.A(n_1747),
.B(n_1796),
.C(n_1769),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1830),
.A2(n_568),
.B(n_566),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1777),
.B(n_15),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1807),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1715),
.B(n_17),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1690),
.Y(n_2067)
);

AND2x6_ASAP7_75t_L g2068 ( 
.A(n_1846),
.B(n_573),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1823),
.B(n_1839),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1766),
.B(n_17),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1621),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1852),
.A2(n_581),
.B(n_578),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1842),
.A2(n_586),
.B(n_582),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_1790),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1722),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1625),
.Y(n_2076)
);

O2A1O1Ixp33_ASAP7_75t_L g2077 ( 
.A1(n_1736),
.A2(n_21),
.B(n_18),
.C(n_19),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1855),
.A2(n_589),
.B(n_588),
.Y(n_2078)
);

O2A1O1Ixp33_ASAP7_75t_L g2079 ( 
.A1(n_1735),
.A2(n_24),
.B(n_21),
.C(n_22),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1722),
.B(n_24),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1783),
.A2(n_1643),
.B1(n_1746),
.B2(n_1849),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1778),
.B(n_26),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1618),
.B(n_592),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1710),
.Y(n_2084)
);

AOI21xp5_ASAP7_75t_L g2085 ( 
.A1(n_1861),
.A2(n_595),
.B(n_594),
.Y(n_2085)
);

OAI321xp33_ASAP7_75t_L g2086 ( 
.A1(n_1840),
.A2(n_29),
.A3(n_32),
.B1(n_27),
.B2(n_28),
.C(n_31),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1778),
.B(n_29),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1862),
.A2(n_1882),
.B(n_1880),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1625),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1763),
.B(n_1774),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1715),
.B(n_33),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1883),
.A2(n_601),
.B(n_599),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1772),
.B(n_34),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1776),
.B(n_34),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1657),
.B(n_35),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1780),
.B(n_36),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1873),
.A2(n_1811),
.B(n_1815),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1780),
.B(n_36),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1717),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1712),
.B(n_37),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1833),
.B(n_38),
.Y(n_2101)
);

XNOR2xp5_ASAP7_75t_L g2102 ( 
.A(n_1802),
.B(n_39),
.Y(n_2102)
);

NOR2x1_ASAP7_75t_L g2103 ( 
.A(n_1617),
.B(n_39),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_1762),
.A2(n_607),
.B(n_606),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1775),
.B(n_40),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1660),
.B(n_41),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1790),
.B(n_43),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1664),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1632),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1886),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1688),
.B(n_45),
.Y(n_2111)
);

O2A1O1Ixp33_ASAP7_75t_L g2112 ( 
.A1(n_1693),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2112)
);

AND2x2_ASAP7_75t_SL g2113 ( 
.A(n_1827),
.B(n_47),
.Y(n_2113)
);

BUFx4f_ASAP7_75t_L g2114 ( 
.A(n_1684),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1816),
.B(n_1697),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1710),
.B(n_48),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1834),
.A2(n_610),
.B(n_609),
.Y(n_2117)
);

O2A1O1Ixp33_ASAP7_75t_L g2118 ( 
.A1(n_1708),
.A2(n_51),
.B(n_48),
.C(n_49),
.Y(n_2118)
);

BUFx12f_ASAP7_75t_L g2119 ( 
.A(n_1876),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1833),
.B(n_49),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1787),
.B(n_55),
.Y(n_2121)
);

CKINVDCx20_ASAP7_75t_R g2122 ( 
.A(n_1684),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1660),
.B(n_55),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1720),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1741),
.B(n_59),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1793),
.B(n_61),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_1684),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1730),
.A2(n_618),
.B(n_615),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1889),
.A2(n_621),
.B(n_620),
.Y(n_2129)
);

INVx1_ASAP7_75t_SL g2130 ( 
.A(n_1804),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1618),
.B(n_622),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1879),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1742),
.B(n_62),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1665),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1849),
.A2(n_1818),
.B1(n_1734),
.B2(n_1733),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1770),
.B(n_63),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1670),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1813),
.B(n_63),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1673),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_1686),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1798),
.B(n_64),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_1800),
.B(n_65),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1781),
.A2(n_625),
.B(n_623),
.Y(n_2143)
);

O2A1O1Ixp5_ASAP7_75t_SL g2144 ( 
.A1(n_1723),
.A2(n_627),
.B(n_628),
.C(n_626),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1812),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1837),
.B(n_1890),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1781),
.A2(n_631),
.B(n_632),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1679),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1837),
.B(n_70),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1818),
.A2(n_74),
.B1(n_71),
.B2(n_73),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1890),
.B(n_1863),
.Y(n_2151)
);

AOI222xp33_ASAP7_75t_L g2152 ( 
.A1(n_1728),
.A2(n_77),
.B1(n_79),
.B2(n_75),
.C1(n_76),
.C2(n_78),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1870),
.A2(n_79),
.B1(n_75),
.B2(n_78),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_1707),
.A2(n_80),
.B(n_81),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1788),
.B(n_80),
.Y(n_2155)
);

BUFx4f_ASAP7_75t_L g2156 ( 
.A(n_1789),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_1877),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1805),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1838),
.B(n_82),
.Y(n_2159)
);

AOI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_1765),
.A2(n_84),
.B(n_85),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1771),
.A2(n_84),
.B(n_85),
.Y(n_2161)
);

AOI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_1779),
.A2(n_86),
.B(n_87),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_1656),
.A2(n_89),
.B(n_90),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1801),
.B(n_89),
.Y(n_2164)
);

O2A1O1Ixp5_ASAP7_75t_L g2165 ( 
.A1(n_1725),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2165)
);

NAND2xp33_ASAP7_75t_SL g2166 ( 
.A(n_1872),
.B(n_93),
.Y(n_2166)
);

OAI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_1714),
.A2(n_96),
.B(n_97),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1803),
.B(n_96),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1767),
.B(n_97),
.Y(n_2169)
);

OAI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1851),
.A2(n_99),
.B(n_101),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1616),
.B(n_102),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_1814),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1732),
.A2(n_102),
.B(n_104),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1865),
.B(n_104),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1884),
.B(n_105),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1868),
.B(n_106),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1737),
.A2(n_1752),
.B(n_1750),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1885),
.B(n_107),
.Y(n_2178)
);

OAI321xp33_ASAP7_75t_L g2179 ( 
.A1(n_1866),
.A2(n_109),
.A3(n_112),
.B1(n_107),
.B2(n_108),
.C(n_110),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1814),
.Y(n_2180)
);

AND2x2_ASAP7_75t_SL g2181 ( 
.A(n_1829),
.B(n_109),
.Y(n_2181)
);

A2O1A1Ixp33_ASAP7_75t_L g2182 ( 
.A1(n_1760),
.A2(n_115),
.B(n_110),
.C(n_113),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_1806),
.B(n_113),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1647),
.A2(n_115),
.B(n_116),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1727),
.A2(n_116),
.B(n_118),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1819),
.B(n_118),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1878),
.Y(n_2187)
);

AOI21x1_ASAP7_75t_L g2188 ( 
.A1(n_1738),
.A2(n_119),
.B(n_120),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_1828),
.B(n_119),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1856),
.B(n_120),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_1740),
.B(n_121),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1856),
.B(n_121),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1745),
.B(n_122),
.Y(n_2193)
);

O2A1O1Ixp33_ASAP7_75t_L g2194 ( 
.A1(n_1757),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1794),
.A2(n_124),
.B(n_126),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_1795),
.A2(n_127),
.B(n_128),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1754),
.Y(n_2197)
);

O2A1O1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_1785),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_1785),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_1618),
.A2(n_130),
.B(n_132),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1618),
.B(n_133),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1618),
.B(n_133),
.Y(n_2202)
);

NOR2xp67_ASAP7_75t_L g2203 ( 
.A(n_1872),
.B(n_134),
.Y(n_2203)
);

O2A1O1Ixp5_ASAP7_75t_L g2204 ( 
.A1(n_1661),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2204)
);

AOI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1661),
.A2(n_136),
.B(n_137),
.Y(n_2205)
);

AOI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_1661),
.A2(n_139),
.B(n_140),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_1663),
.B(n_139),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_1661),
.A2(n_140),
.B(n_141),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1668),
.B(n_141),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_1786),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1668),
.A2(n_146),
.B1(n_143),
.B2(n_144),
.Y(n_2211)
);

O2A1O1Ixp5_ASAP7_75t_L g2212 ( 
.A1(n_1661),
.A2(n_150),
.B(n_147),
.C(n_149),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1967),
.B(n_150),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2047),
.B(n_152),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_1968),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_2140),
.B(n_2090),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2046),
.B(n_155),
.Y(n_2217)
);

AO21x1_ASAP7_75t_L g2218 ( 
.A1(n_2200),
.A2(n_156),
.B(n_157),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2088),
.A2(n_156),
.B(n_157),
.Y(n_2219)
);

AOI21x1_ASAP7_75t_L g2220 ( 
.A1(n_1924),
.A2(n_158),
.B(n_159),
.Y(n_2220)
);

O2A1O1Ixp33_ASAP7_75t_L g2221 ( 
.A1(n_2146),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2221)
);

AND3x1_ASAP7_75t_SL g2222 ( 
.A(n_2045),
.B(n_2003),
.C(n_2119),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_1898),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_2047),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_1905),
.A2(n_164),
.B(n_165),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_R g2226 ( 
.A(n_2122),
.B(n_164),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1898),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_2156),
.B(n_1996),
.Y(n_2228)
);

CKINVDCx12_ASAP7_75t_R g2229 ( 
.A(n_1901),
.Y(n_2229)
);

O2A1O1Ixp33_ASAP7_75t_L g2230 ( 
.A1(n_2101),
.A2(n_169),
.B(n_166),
.C(n_167),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1973),
.B(n_167),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1921),
.B(n_169),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1948),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2010),
.B(n_170),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_1921),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_1894),
.A2(n_171),
.B(n_173),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1897),
.Y(n_2237)
);

NOR2xp67_ASAP7_75t_SL g2238 ( 
.A(n_2018),
.B(n_174),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_1983),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2097),
.A2(n_176),
.B(n_177),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2029),
.B(n_176),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2113),
.B(n_177),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1893),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2009),
.B(n_2019),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_2156),
.B(n_178),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1999),
.B(n_2050),
.Y(n_2246)
);

OR2x6_ASAP7_75t_L g2247 ( 
.A(n_2075),
.B(n_179),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2151),
.B(n_180),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2135),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2099),
.B(n_181),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2124),
.B(n_1990),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_2067),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2012),
.B(n_185),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1907),
.B(n_1911),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1912),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2062),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_1939),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1931),
.B(n_191),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1999),
.B(n_192),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1943),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_1940),
.B(n_194),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2113),
.B(n_195),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1950),
.B(n_196),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2062),
.B(n_196),
.C(n_197),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2181),
.B(n_198),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2049),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2050),
.B(n_199),
.Y(n_2267)
);

AOI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2069),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_1895),
.B(n_200),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_1902),
.A2(n_201),
.B(n_203),
.Y(n_2270)
);

O2A1O1Ixp33_ASAP7_75t_L g2271 ( 
.A1(n_2120),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2053),
.B(n_208),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2053),
.B(n_208),
.Y(n_2273)
);

OR2x6_ASAP7_75t_L g2274 ( 
.A(n_1942),
.B(n_209),
.Y(n_2274)
);

BUFx8_ASAP7_75t_SL g2275 ( 
.A(n_2071),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2181),
.B(n_210),
.Y(n_2276)
);

NAND3xp33_ASAP7_75t_SL g2277 ( 
.A(n_2152),
.B(n_211),
.C(n_212),
.Y(n_2277)
);

AOI21x1_ASAP7_75t_L g2278 ( 
.A1(n_1979),
.A2(n_212),
.B(n_213),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_1949),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2041),
.Y(n_2280)
);

O2A1O1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_1900),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1936),
.B(n_216),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1951),
.B(n_217),
.Y(n_2283)
);

INVx4_ASAP7_75t_L g2284 ( 
.A(n_1983),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_2012),
.Y(n_2285)
);

INVx6_ASAP7_75t_L g2286 ( 
.A(n_1976),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_1896),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2012),
.B(n_223),
.Y(n_2288)
);

OAI22x1_ASAP7_75t_L g2289 ( 
.A1(n_2108),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1949),
.B(n_224),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2051),
.Y(n_2291)
);

OAI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_1899),
.A2(n_225),
.B(n_226),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1969),
.B(n_227),
.Y(n_2293)
);

A2O1A1Ixp33_ASAP7_75t_L g2294 ( 
.A1(n_1899),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2065),
.Y(n_2295)
);

O2A1O1Ixp5_ASAP7_75t_L g2296 ( 
.A1(n_1961),
.A2(n_231),
.B(n_228),
.C(n_230),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2081),
.A2(n_234),
.B1(n_231),
.B2(n_233),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1969),
.B(n_233),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2114),
.B(n_235),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2132),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2084),
.B(n_235),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2052),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2064),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2114),
.B(n_236),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2048),
.B(n_237),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2084),
.B(n_237),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1925),
.B(n_238),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2107),
.Y(n_2308)
);

O2A1O1Ixp33_ASAP7_75t_SL g2309 ( 
.A1(n_2056),
.A2(n_241),
.B(n_238),
.C(n_239),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2021),
.B(n_244),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_2048),
.B(n_244),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2134),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2137),
.Y(n_2313)
);

A2O1A1Ixp33_ASAP7_75t_L g2314 ( 
.A1(n_2125),
.A2(n_254),
.B(n_251),
.C(n_252),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2139),
.Y(n_2315)
);

O2A1O1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_1908),
.A2(n_2058),
.B(n_2209),
.C(n_1913),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1975),
.A2(n_1909),
.B1(n_2211),
.B2(n_2115),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_2012),
.Y(n_2318)
);

A2O1A1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2125),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_1910),
.A2(n_259),
.B(n_260),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2035),
.B(n_261),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_1944),
.B(n_262),
.Y(n_2322)
);

BUFx3_ASAP7_75t_L g2323 ( 
.A(n_1980),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1904),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2148),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2116),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2111),
.Y(n_2327)
);

NOR3xp33_ASAP7_75t_SL g2328 ( 
.A(n_2080),
.B(n_266),
.C(n_267),
.Y(n_2328)
);

BUFx12f_ASAP7_75t_L g2329 ( 
.A(n_1904),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_1915),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2070),
.B(n_268),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1915),
.A2(n_2133),
.B1(n_2136),
.B2(n_2060),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_1914),
.B(n_271),
.Y(n_2333)
);

AO32x1_ASAP7_75t_L g2334 ( 
.A1(n_2171),
.A2(n_274),
.A3(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_1901),
.Y(n_2335)
);

CKINVDCx16_ASAP7_75t_R g2336 ( 
.A(n_1929),
.Y(n_2336)
);

A2O1A1Ixp33_ASAP7_75t_SL g2337 ( 
.A1(n_2133),
.A2(n_277),
.B(n_274),
.C(n_276),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_2130),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_1966),
.B(n_276),
.Y(n_2339)
);

O2A1O1Ixp33_ASAP7_75t_L g2340 ( 
.A1(n_2141),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2340)
);

INVx5_ASAP7_75t_L g2341 ( 
.A(n_1901),
.Y(n_2341)
);

O2A1O1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_2175),
.A2(n_283),
.B(n_280),
.C(n_282),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2138),
.B(n_280),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_1919),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2136),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2105),
.B(n_284),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_1930),
.B(n_286),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1972),
.Y(n_2348)
);

CKINVDCx20_ASAP7_75t_R g2349 ( 
.A(n_1919),
.Y(n_2349)
);

O2A1O1Ixp5_ASAP7_75t_L g2350 ( 
.A1(n_1938),
.A2(n_290),
.B(n_287),
.C(n_289),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2095),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_2351)
);

NAND3xp33_ASAP7_75t_SL g2352 ( 
.A(n_2054),
.B(n_294),
.C(n_295),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_1982),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2210),
.B(n_296),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_1930),
.B(n_296),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_1966),
.B(n_298),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_1927),
.A2(n_298),
.B(n_299),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_2210),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2111),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2000),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_1937),
.A2(n_299),
.B(n_300),
.Y(n_2361)
);

AOI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_1932),
.A2(n_300),
.B(n_301),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_1982),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_1916),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2036),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_1982),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_SL g2367 ( 
.A1(n_2102),
.A2(n_2054),
.B1(n_2055),
.B2(n_2145),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2024),
.B(n_303),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2013),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2188),
.Y(n_2370)
);

O2A1O1Ixp33_ASAP7_75t_L g2371 ( 
.A1(n_2079),
.A2(n_306),
.B(n_303),
.C(n_305),
.Y(n_2371)
);

A2O1A1Ixp33_ASAP7_75t_L g2372 ( 
.A1(n_2077),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2372)
);

OAI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_1906),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_2373)
);

INVx5_ASAP7_75t_L g2374 ( 
.A(n_2068),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2150),
.A2(n_311),
.B1(n_308),
.B2(n_310),
.Y(n_2375)
);

INVxp67_ASAP7_75t_L g2376 ( 
.A(n_2207),
.Y(n_2376)
);

AOI21xp33_ASAP7_75t_L g2377 ( 
.A1(n_2100),
.A2(n_312),
.B(n_313),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1993),
.B(n_313),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_1982),
.Y(n_2379)
);

O2A1O1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_2002),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2149),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_1933),
.A2(n_318),
.B(n_319),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2189),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2076),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2158),
.B(n_321),
.Y(n_2385)
);

OAI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2155),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2203),
.B(n_323),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2055),
.Y(n_2388)
);

NOR3xp33_ASAP7_75t_SL g2389 ( 
.A(n_2086),
.B(n_325),
.C(n_326),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2014),
.B(n_327),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_1992),
.B(n_328),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_1974),
.A2(n_1920),
.B(n_2082),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2089),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_1994),
.B(n_330),
.Y(n_2394)
);

INVx2_ASAP7_75t_SL g2395 ( 
.A(n_2127),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2028),
.Y(n_2396)
);

OAI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_1974),
.A2(n_331),
.B(n_332),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_1997),
.Y(n_2398)
);

CKINVDCx11_ASAP7_75t_R g2399 ( 
.A(n_1986),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_1916),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1916),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2008),
.B(n_333),
.Y(n_2402)
);

A2O1A1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_2066),
.A2(n_2091),
.B(n_2098),
.C(n_2096),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_1923),
.A2(n_333),
.B(n_335),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_1977),
.B(n_336),
.Y(n_2405)
);

A2O1A1Ixp33_ASAP7_75t_L g2406 ( 
.A1(n_2066),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2191),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_1926),
.A2(n_340),
.B(n_341),
.Y(n_2408)
);

OR2x6_ASAP7_75t_L g2409 ( 
.A(n_1986),
.B(n_2007),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2174),
.Y(n_2410)
);

BUFx2_ASAP7_75t_L g2411 ( 
.A(n_1989),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_1922),
.A2(n_342),
.B(n_344),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2204),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_1916),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2023),
.B(n_346),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2093),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_2416)
);

AO32x1_ASAP7_75t_L g2417 ( 
.A1(n_2153),
.A2(n_347),
.A3(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_2417)
);

OAI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2087),
.A2(n_350),
.B(n_351),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2158),
.B(n_352),
.Y(n_2419)
);

O2A1O1Ixp33_ASAP7_75t_L g2420 ( 
.A1(n_2027),
.A2(n_353),
.B(n_354),
.C(n_356),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2094),
.A2(n_354),
.B1(n_356),
.B2(n_358),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_1986),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2176),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_1971),
.Y(n_2424)
);

A2O1A1Ixp33_ASAP7_75t_L g2425 ( 
.A1(n_2091),
.A2(n_359),
.B(n_360),
.C(n_361),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2074),
.B(n_359),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_SL g2427 ( 
.A(n_1956),
.B(n_360),
.Y(n_2427)
);

NAND3xp33_ASAP7_75t_L g2428 ( 
.A(n_2026),
.B(n_361),
.C(n_362),
.Y(n_2428)
);

A2O1A1Ixp33_ASAP7_75t_SL g2429 ( 
.A1(n_1935),
.A2(n_2170),
.B(n_2154),
.C(n_2167),
.Y(n_2429)
);

INVx4_ASAP7_75t_L g2430 ( 
.A(n_1986),
.Y(n_2430)
);

O2A1O1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2032),
.A2(n_362),
.B(n_363),
.C(n_364),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1978),
.B(n_364),
.Y(n_2432)
);

A2O1A1Ixp33_ASAP7_75t_L g2433 ( 
.A1(n_2096),
.A2(n_367),
.B(n_368),
.C(n_369),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_1989),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_1971),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2186),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_1984),
.B(n_370),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2007),
.B(n_370),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2057),
.A2(n_371),
.B1(n_372),
.B2(n_374),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1981),
.B(n_371),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_1917),
.A2(n_377),
.B(n_378),
.Y(n_2441)
);

O2A1O1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_1985),
.A2(n_378),
.B(n_379),
.C(n_380),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_1946),
.B(n_379),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2015),
.B(n_380),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2007),
.B(n_2020),
.Y(n_2445)
);

AOI222xp33_ASAP7_75t_L g2446 ( 
.A1(n_2006),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.C1(n_384),
.C2(n_385),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1988),
.B(n_381),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1918),
.B(n_382),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2192),
.Y(n_2449)
);

NAND3xp33_ASAP7_75t_SL g2450 ( 
.A(n_1952),
.B(n_385),
.C(n_386),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2017),
.B(n_1941),
.Y(n_2451)
);

A2O1A1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_2098),
.A2(n_386),
.B(n_387),
.C(n_388),
.Y(n_2452)
);

OAI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2159),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_2453)
);

AOI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2142),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1947),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2007),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_SL g2457 ( 
.A(n_2068),
.B(n_390),
.Y(n_2457)
);

O2A1O1Ixp5_ASAP7_75t_L g2458 ( 
.A1(n_2011),
.A2(n_392),
.B(n_393),
.C(n_395),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1955),
.B(n_396),
.Y(n_2459)
);

INVx6_ASAP7_75t_L g2460 ( 
.A(n_2158),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2001),
.B(n_397),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1957),
.Y(n_2462)
);

AOI22xp33_ASAP7_75t_L g2463 ( 
.A1(n_1952),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_2463)
);

AND2x6_ASAP7_75t_L g2464 ( 
.A(n_2020),
.B(n_2040),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1959),
.B(n_401),
.Y(n_2465)
);

O2A1O1Ixp33_ASAP7_75t_L g2466 ( 
.A1(n_2157),
.A2(n_2126),
.B(n_2121),
.C(n_2198),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2037),
.A2(n_402),
.B(n_403),
.Y(n_2467)
);

NAND3xp33_ASAP7_75t_L g2468 ( 
.A(n_2389),
.B(n_1935),
.C(n_2212),
.Y(n_2468)
);

BUFx2_ASAP7_75t_SL g2469 ( 
.A(n_2284),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2457),
.A2(n_2429),
.B(n_2392),
.Y(n_2470)
);

AOI221xp5_ASAP7_75t_SL g2471 ( 
.A1(n_2367),
.A2(n_2162),
.B1(n_2161),
.B2(n_2160),
.C(n_2182),
.Y(n_2471)
);

NAND2xp33_ASAP7_75t_SL g2472 ( 
.A(n_2226),
.B(n_2106),
.Y(n_2472)
);

OAI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2403),
.A2(n_2165),
.B(n_2205),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2235),
.Y(n_2474)
);

HB1xp67_ASAP7_75t_L g2475 ( 
.A(n_2279),
.Y(n_2475)
);

INVx2_ASAP7_75t_SL g2476 ( 
.A(n_2286),
.Y(n_2476)
);

OAI21x1_ASAP7_75t_L g2477 ( 
.A1(n_2370),
.A2(n_2004),
.B(n_1903),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2367),
.A2(n_2332),
.B1(n_2374),
.B2(n_2308),
.Y(n_2478)
);

OAI21x1_ASAP7_75t_L g2479 ( 
.A1(n_2413),
.A2(n_1995),
.B(n_2144),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2237),
.Y(n_2480)
);

OAI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2332),
.A2(n_2316),
.B(n_2317),
.Y(n_2481)
);

OA21x2_ASAP7_75t_L g2482 ( 
.A1(n_2397),
.A2(n_2073),
.B(n_2104),
.Y(n_2482)
);

BUFx10_ASAP7_75t_L g2483 ( 
.A(n_2247),
.Y(n_2483)
);

BUFx2_ASAP7_75t_L g2484 ( 
.A(n_2224),
.Y(n_2484)
);

AOI21x1_ASAP7_75t_L g2485 ( 
.A1(n_2278),
.A2(n_2131),
.B(n_2083),
.Y(n_2485)
);

AOI21x1_ASAP7_75t_L g2486 ( 
.A1(n_2242),
.A2(n_2201),
.B(n_2022),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2441),
.A2(n_1970),
.B(n_1963),
.Y(n_2487)
);

AO21x2_ASAP7_75t_L g2488 ( 
.A1(n_2225),
.A2(n_2218),
.B(n_2309),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2466),
.A2(n_2449),
.B(n_2410),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2251),
.B(n_2168),
.Y(n_2490)
);

CKINVDCx20_ASAP7_75t_R g2491 ( 
.A(n_2275),
.Y(n_2491)
);

OAI21x1_ASAP7_75t_L g2492 ( 
.A1(n_2220),
.A2(n_2043),
.B(n_1954),
.Y(n_2492)
);

O2A1O1Ixp33_ASAP7_75t_SL g2493 ( 
.A1(n_2262),
.A2(n_2031),
.B(n_2005),
.C(n_2173),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2280),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2260),
.Y(n_2495)
);

OA21x2_ASAP7_75t_L g2496 ( 
.A1(n_2458),
.A2(n_2184),
.B(n_2206),
.Y(n_2496)
);

INVx4_ASAP7_75t_L g2497 ( 
.A(n_2224),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2248),
.A2(n_2044),
.B(n_2072),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2427),
.B(n_2166),
.Y(n_2499)
);

O2A1O1Ixp33_ASAP7_75t_SL g2500 ( 
.A1(n_2265),
.A2(n_2276),
.B(n_2322),
.C(n_2294),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2423),
.A2(n_2085),
.B(n_2078),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2216),
.B(n_2168),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2295),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2396),
.B(n_2187),
.Y(n_2504)
);

AOI221xp5_ASAP7_75t_SL g2505 ( 
.A1(n_2281),
.A2(n_2112),
.B1(n_2118),
.B2(n_2163),
.C(n_2208),
.Y(n_2505)
);

BUFx2_ASAP7_75t_L g2506 ( 
.A(n_2369),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2347),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2246),
.B(n_2183),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2234),
.A2(n_2092),
.B(n_2061),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2337),
.A2(n_2063),
.B(n_2059),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_L g2511 ( 
.A(n_2285),
.B(n_2068),
.Y(n_2511)
);

OAI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2444),
.A2(n_2165),
.B(n_2183),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2446),
.B(n_2194),
.C(n_2193),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2261),
.B(n_1960),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2254),
.Y(n_2515)
);

A2O1A1Ixp33_ASAP7_75t_L g2516 ( 
.A1(n_2371),
.A2(n_2164),
.B(n_2193),
.C(n_1998),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2285),
.B(n_2068),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2455),
.B(n_1962),
.Y(n_2518)
);

OAI21x1_ASAP7_75t_L g2519 ( 
.A1(n_2350),
.A2(n_2129),
.B(n_2128),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2228),
.B(n_1965),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2388),
.B(n_2169),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2291),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2219),
.A2(n_1945),
.B(n_2030),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2239),
.Y(n_2524)
);

OAI21x1_ASAP7_75t_L g2525 ( 
.A1(n_2335),
.A2(n_2147),
.B(n_2143),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2462),
.B(n_2178),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2240),
.A2(n_2117),
.B(n_2177),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2244),
.B(n_2025),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_2323),
.Y(n_2529)
);

OAI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2345),
.A2(n_2123),
.B1(n_2103),
.B2(n_2172),
.Y(n_2530)
);

OAI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2345),
.A2(n_2249),
.B1(n_2247),
.B2(n_2375),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2321),
.A2(n_2196),
.B(n_2195),
.Y(n_2532)
);

CKINVDCx20_ASAP7_75t_R g2533 ( 
.A(n_2399),
.Y(n_2533)
);

AOI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_2272),
.A2(n_2273),
.B(n_2231),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_SL g2535 ( 
.A1(n_2247),
.A2(n_2068),
.B1(n_2202),
.B2(n_2172),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2259),
.B(n_2033),
.Y(n_2536)
);

OAI21x1_ASAP7_75t_L g2537 ( 
.A1(n_2335),
.A2(n_1928),
.B(n_1987),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2233),
.B(n_2199),
.Y(n_2538)
);

OAI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2296),
.A2(n_2372),
.B(n_2451),
.Y(n_2539)
);

OAI21x1_ASAP7_75t_L g2540 ( 
.A1(n_2302),
.A2(n_1991),
.B(n_2039),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2436),
.A2(n_1934),
.B(n_1953),
.Y(n_2541)
);

NOR2x1p5_ASAP7_75t_L g2542 ( 
.A(n_2284),
.B(n_2040),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2266),
.B(n_2034),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2312),
.Y(n_2544)
);

OA21x2_ASAP7_75t_L g2545 ( 
.A1(n_2236),
.A2(n_2185),
.B(n_2179),
.Y(n_2545)
);

AO21x1_ASAP7_75t_L g2546 ( 
.A1(n_2256),
.A2(n_2190),
.B(n_2016),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2223),
.A2(n_2197),
.B(n_1958),
.Y(n_2547)
);

O2A1O1Ixp33_ASAP7_75t_SL g2548 ( 
.A1(n_2314),
.A2(n_2199),
.B(n_2180),
.C(n_2042),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2318),
.Y(n_2549)
);

AO31x2_ASAP7_75t_L g2550 ( 
.A1(n_2467),
.A2(n_2038),
.A3(n_1964),
.B(n_2109),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2313),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2383),
.B(n_2042),
.Y(n_2552)
);

O2A1O1Ixp33_ASAP7_75t_SL g2553 ( 
.A1(n_2319),
.A2(n_2180),
.B(n_2158),
.C(n_2109),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2223),
.A2(n_2109),
.B(n_2110),
.Y(n_2554)
);

OAI21x1_ASAP7_75t_L g2555 ( 
.A1(n_2363),
.A2(n_2110),
.B(n_2109),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2407),
.B(n_404),
.Y(n_2556)
);

AOI221x1_ASAP7_75t_L g2557 ( 
.A1(n_2264),
.A2(n_2110),
.B1(n_406),
.B2(n_407),
.C(n_408),
.Y(n_2557)
);

BUFx12f_ASAP7_75t_L g2558 ( 
.A(n_2215),
.Y(n_2558)
);

AO21x1_ASAP7_75t_L g2559 ( 
.A1(n_2256),
.A2(n_405),
.B(n_409),
.Y(n_2559)
);

A2O1A1Ixp33_ASAP7_75t_L g2560 ( 
.A1(n_2292),
.A2(n_2110),
.B(n_410),
.C(n_411),
.Y(n_2560)
);

INVxp67_ASAP7_75t_L g2561 ( 
.A(n_2274),
.Y(n_2561)
);

NAND2x1_ASAP7_75t_L g2562 ( 
.A(n_2318),
.B(n_409),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2315),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2325),
.Y(n_2564)
);

AOI221xp5_ASAP7_75t_SL g2565 ( 
.A1(n_2373),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.C(n_414),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2223),
.A2(n_412),
.B(n_415),
.Y(n_2566)
);

BUFx3_ASAP7_75t_L g2567 ( 
.A(n_2252),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2341),
.B(n_415),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2347),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2243),
.Y(n_2570)
);

A2O1A1Ixp33_ASAP7_75t_L g2571 ( 
.A1(n_2249),
.A2(n_416),
.B(n_417),
.C(n_418),
.Y(n_2571)
);

HB1xp67_ASAP7_75t_L g2572 ( 
.A(n_2355),
.Y(n_2572)
);

OAI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2277),
.A2(n_416),
.B(n_417),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2255),
.Y(n_2574)
);

A2O1A1Ixp33_ASAP7_75t_L g2575 ( 
.A1(n_2361),
.A2(n_422),
.B(n_423),
.C(n_424),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2227),
.A2(n_422),
.B(n_423),
.Y(n_2576)
);

OAI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2310),
.A2(n_424),
.B(n_425),
.Y(n_2577)
);

A2O1A1Ixp33_ASAP7_75t_L g2578 ( 
.A1(n_2297),
.A2(n_427),
.B(n_428),
.C(n_429),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_2329),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2360),
.Y(n_2580)
);

AO31x2_ASAP7_75t_L g2581 ( 
.A1(n_2406),
.A2(n_2425),
.A3(n_2452),
.B(n_2433),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2327),
.B(n_2326),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2424),
.Y(n_2583)
);

AOI31xp67_ASAP7_75t_L g2584 ( 
.A1(n_2297),
.A2(n_430),
.A3(n_431),
.B(n_432),
.Y(n_2584)
);

CKINVDCx6p67_ASAP7_75t_R g2585 ( 
.A(n_2274),
.Y(n_2585)
);

OAI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2366),
.A2(n_431),
.B(n_433),
.Y(n_2586)
);

NAND2x1_ASAP7_75t_L g2587 ( 
.A(n_2460),
.B(n_434),
.Y(n_2587)
);

AO32x2_ASAP7_75t_L g2588 ( 
.A1(n_2330),
.A2(n_434),
.A3(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_2588)
);

OAI21x1_ASAP7_75t_L g2589 ( 
.A1(n_2379),
.A2(n_2362),
.B(n_2357),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2267),
.A2(n_438),
.B(n_439),
.Y(n_2590)
);

NAND3x1_ASAP7_75t_L g2591 ( 
.A(n_2245),
.B(n_442),
.C(n_443),
.Y(n_2591)
);

AO31x2_ASAP7_75t_L g2592 ( 
.A1(n_2270),
.A2(n_443),
.A3(n_445),
.B(n_446),
.Y(n_2592)
);

AOI31xp67_ASAP7_75t_L g2593 ( 
.A1(n_2385),
.A2(n_446),
.A3(n_447),
.B(n_449),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2359),
.B(n_447),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2303),
.B(n_2443),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2217),
.B(n_449),
.Y(n_2596)
);

CKINVDCx11_ASAP7_75t_R g2597 ( 
.A(n_2257),
.Y(n_2597)
);

OAI21x1_ASAP7_75t_L g2598 ( 
.A1(n_2382),
.A2(n_451),
.B(n_452),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2352),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_2599)
);

BUFx2_ASAP7_75t_SL g2600 ( 
.A(n_2214),
.Y(n_2600)
);

AOI21x1_ASAP7_75t_L g2601 ( 
.A1(n_2419),
.A2(n_454),
.B(n_455),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2364),
.A2(n_455),
.B(n_456),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2341),
.B(n_456),
.Y(n_2603)
);

O2A1O1Ixp33_ASAP7_75t_L g2604 ( 
.A1(n_2331),
.A2(n_457),
.B(n_459),
.C(n_460),
.Y(n_2604)
);

AOI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2400),
.A2(n_457),
.B(n_460),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2376),
.B(n_461),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2448),
.B(n_550),
.Y(n_2607)
);

INVxp67_ASAP7_75t_L g2608 ( 
.A(n_2274),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2349),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2324),
.Y(n_2610)
);

A2O1A1Ixp33_ASAP7_75t_L g2611 ( 
.A1(n_2420),
.A2(n_462),
.B(n_463),
.C(n_464),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_2336),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2343),
.B(n_549),
.Y(n_2613)
);

NAND3xp33_ASAP7_75t_L g2614 ( 
.A(n_2428),
.B(n_467),
.C(n_468),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2263),
.B(n_467),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2341),
.B(n_468),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2348),
.Y(n_2617)
);

OAI21x1_ASAP7_75t_L g2618 ( 
.A1(n_2404),
.A2(n_469),
.B(n_471),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2346),
.B(n_548),
.Y(n_2619)
);

NAND3xp33_ASAP7_75t_SL g2620 ( 
.A(n_2454),
.B(n_469),
.C(n_472),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2368),
.B(n_472),
.Y(n_2621)
);

AO21x2_ASAP7_75t_L g2622 ( 
.A1(n_2418),
.A2(n_548),
.B(n_474),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2300),
.B(n_473),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2401),
.A2(n_473),
.B(n_474),
.Y(n_2624)
);

OAI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_2378),
.A2(n_2390),
.B(n_2459),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_2344),
.Y(n_2626)
);

BUFx12f_ASAP7_75t_L g2627 ( 
.A(n_2358),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2375),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2338),
.B(n_477),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2232),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2414),
.A2(n_478),
.B(n_479),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2408),
.A2(n_480),
.B(n_481),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2412),
.A2(n_480),
.B(n_481),
.Y(n_2633)
);

AO31x2_ASAP7_75t_L g2634 ( 
.A1(n_2320),
.A2(n_482),
.A3(n_485),
.B(n_486),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2282),
.B(n_2213),
.Y(n_2635)
);

AOI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2414),
.A2(n_487),
.B(n_488),
.Y(n_2636)
);

NOR4xp25_ASAP7_75t_L g2637 ( 
.A(n_2221),
.B(n_487),
.C(n_489),
.D(n_491),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2435),
.B(n_489),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2405),
.A2(n_491),
.B(n_492),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2355),
.Y(n_2640)
);

A2O1A1Ixp33_ASAP7_75t_L g2641 ( 
.A1(n_2431),
.A2(n_493),
.B(n_494),
.C(n_495),
.Y(n_2641)
);

INVx4_ASAP7_75t_L g2642 ( 
.A(n_2497),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2480),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_SL g2644 ( 
.A1(n_2531),
.A2(n_2214),
.B1(n_2253),
.B2(n_2288),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2495),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_SL g2646 ( 
.A(n_2535),
.B(n_2253),
.Y(n_2646)
);

HB1xp67_ASAP7_75t_L g2647 ( 
.A(n_2474),
.Y(n_2647)
);

INVx6_ASAP7_75t_L g2648 ( 
.A(n_2497),
.Y(n_2648)
);

OAI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2585),
.A2(n_2289),
.B1(n_2307),
.B2(n_2450),
.Y(n_2649)
);

OAI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2616),
.A2(n_2293),
.B1(n_2290),
.B2(n_2387),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_2478),
.A2(n_2311),
.B1(n_2305),
.B2(n_2288),
.Y(n_2651)
);

BUFx8_ASAP7_75t_L g2652 ( 
.A(n_2558),
.Y(n_2652)
);

INVx6_ASAP7_75t_L g2653 ( 
.A(n_2529),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2503),
.Y(n_2654)
);

OAI22xp33_ASAP7_75t_R g2655 ( 
.A1(n_2579),
.A2(n_2356),
.B1(n_2339),
.B2(n_2461),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2544),
.Y(n_2656)
);

INVx6_ASAP7_75t_L g2657 ( 
.A(n_2567),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2508),
.A2(n_2437),
.B1(n_2377),
.B2(n_2386),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2474),
.B(n_2298),
.Y(n_2659)
);

CKINVDCx11_ASAP7_75t_R g2660 ( 
.A(n_2533),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2638),
.B(n_2365),
.Y(n_2661)
);

INVx6_ASAP7_75t_L g2662 ( 
.A(n_2483),
.Y(n_2662)
);

BUFx12f_ASAP7_75t_L g2663 ( 
.A(n_2597),
.Y(n_2663)
);

INVx1_ASAP7_75t_SL g2664 ( 
.A(n_2506),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2484),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2517),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2515),
.B(n_2398),
.Y(n_2667)
);

BUFx2_ASAP7_75t_L g2668 ( 
.A(n_2627),
.Y(n_2668)
);

OAI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2600),
.A2(n_2328),
.B1(n_2463),
.B2(n_2287),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2563),
.Y(n_2670)
);

OAI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2616),
.A2(n_2283),
.B1(n_2411),
.B2(n_2434),
.Y(n_2671)
);

BUFx4f_ASAP7_75t_SL g2672 ( 
.A(n_2491),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2513),
.A2(n_2620),
.B1(n_2481),
.B2(n_2472),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2513),
.A2(n_2380),
.B(n_2442),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_SL g2675 ( 
.A1(n_2483),
.A2(n_2438),
.B1(n_2381),
.B2(n_2351),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2564),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2511),
.Y(n_2677)
);

OAI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2628),
.A2(n_2439),
.B1(n_2304),
.B2(n_2299),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2551),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2617),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2630),
.B(n_2384),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2475),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2494),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2522),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2546),
.A2(n_2394),
.B1(n_2391),
.B2(n_2453),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2628),
.A2(n_2438),
.B1(n_2268),
.B2(n_2333),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2502),
.A2(n_2421),
.B1(n_2416),
.B2(n_2354),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_L g2688 ( 
.A(n_2517),
.Y(n_2688)
);

INVx1_ASAP7_75t_SL g2689 ( 
.A(n_2610),
.Y(n_2689)
);

CKINVDCx20_ASAP7_75t_R g2690 ( 
.A(n_2609),
.Y(n_2690)
);

OAI22xp33_ASAP7_75t_L g2691 ( 
.A1(n_2599),
.A2(n_2269),
.B1(n_2241),
.B2(n_2250),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2640),
.A2(n_2306),
.B1(n_2301),
.B2(n_2415),
.Y(n_2692)
);

BUFx4_ASAP7_75t_R g2693 ( 
.A(n_2469),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2559),
.A2(n_2426),
.B1(n_2440),
.B2(n_2447),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2573),
.A2(n_2432),
.B1(n_2238),
.B2(n_2465),
.Y(n_2695)
);

INVx6_ASAP7_75t_L g2696 ( 
.A(n_2542),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2580),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2586),
.Y(n_2698)
);

NAND2x1p5_ASAP7_75t_L g2699 ( 
.A(n_2603),
.B(n_2353),
.Y(n_2699)
);

INVxp67_ASAP7_75t_SL g2700 ( 
.A(n_2507),
.Y(n_2700)
);

INVx5_ASAP7_75t_L g2701 ( 
.A(n_2603),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2596),
.A2(n_2222),
.B1(n_2229),
.B2(n_2258),
.Y(n_2702)
);

INVx6_ASAP7_75t_L g2703 ( 
.A(n_2638),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2583),
.B(n_2393),
.Y(n_2704)
);

BUFx4f_ASAP7_75t_SL g2705 ( 
.A(n_2524),
.Y(n_2705)
);

BUFx2_ASAP7_75t_SL g2706 ( 
.A(n_2476),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_SL g2707 ( 
.A1(n_2569),
.A2(n_2464),
.B1(n_2353),
.B2(n_2422),
.Y(n_2707)
);

BUFx8_ASAP7_75t_SL g2708 ( 
.A(n_2612),
.Y(n_2708)
);

INVx6_ASAP7_75t_L g2709 ( 
.A(n_2538),
.Y(n_2709)
);

BUFx2_ASAP7_75t_L g2710 ( 
.A(n_2561),
.Y(n_2710)
);

BUFx12f_ASAP7_75t_L g2711 ( 
.A(n_2626),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_SL g2712 ( 
.A1(n_2572),
.A2(n_2464),
.B1(n_2430),
.B2(n_2422),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2520),
.A2(n_2402),
.B1(n_2395),
.B2(n_2464),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_SL g2714 ( 
.A1(n_2608),
.A2(n_2590),
.B1(n_2530),
.B2(n_2622),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_2536),
.A2(n_2464),
.B1(n_2445),
.B2(n_2430),
.Y(n_2715)
);

BUFx10_ASAP7_75t_L g2716 ( 
.A(n_2629),
.Y(n_2716)
);

OAI21xp5_ASAP7_75t_SL g2717 ( 
.A1(n_2599),
.A2(n_2342),
.B(n_2340),
.Y(n_2717)
);

INVxp67_ASAP7_75t_SL g2718 ( 
.A(n_2549),
.Y(n_2718)
);

INVx4_ASAP7_75t_L g2719 ( 
.A(n_2549),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2592),
.Y(n_2720)
);

INVxp67_ASAP7_75t_L g2721 ( 
.A(n_2606),
.Y(n_2721)
);

INVx6_ASAP7_75t_L g2722 ( 
.A(n_2514),
.Y(n_2722)
);

INVx4_ASAP7_75t_L g2723 ( 
.A(n_2622),
.Y(n_2723)
);

INVx6_ASAP7_75t_L g2724 ( 
.A(n_2570),
.Y(n_2724)
);

INVx6_ASAP7_75t_L g2725 ( 
.A(n_2574),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2592),
.Y(n_2726)
);

BUFx4f_ASAP7_75t_SL g2727 ( 
.A(n_2499),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2552),
.Y(n_2728)
);

OAI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2578),
.A2(n_2409),
.B1(n_2230),
.B2(n_2271),
.Y(n_2729)
);

OAI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2571),
.A2(n_2409),
.B1(n_2460),
.B2(n_2445),
.Y(n_2730)
);

OAI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2560),
.A2(n_2409),
.B1(n_2456),
.B2(n_2417),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2582),
.Y(n_2732)
);

INVx6_ASAP7_75t_L g2733 ( 
.A(n_2562),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2555),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2595),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2556),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2575),
.A2(n_2456),
.B1(n_2417),
.B2(n_2334),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2550),
.Y(n_2738)
);

BUFx8_ASAP7_75t_L g2739 ( 
.A(n_2588),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2623),
.Y(n_2740)
);

BUFx3_ASAP7_75t_L g2741 ( 
.A(n_2504),
.Y(n_2741)
);

INVx6_ASAP7_75t_L g2742 ( 
.A(n_2591),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2521),
.A2(n_2456),
.B1(n_2417),
.B2(n_2334),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2512),
.A2(n_2334),
.B1(n_495),
.B2(n_496),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2490),
.A2(n_494),
.B1(n_497),
.B2(n_499),
.Y(n_2745)
);

INVx2_ASAP7_75t_SL g2746 ( 
.A(n_2587),
.Y(n_2746)
);

CKINVDCx16_ASAP7_75t_R g2747 ( 
.A(n_2577),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2518),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2615),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2601),
.Y(n_2750)
);

BUFx10_ASAP7_75t_L g2751 ( 
.A(n_2568),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2635),
.B(n_501),
.Y(n_2752)
);

OAI22x1_ASAP7_75t_L g2753 ( 
.A1(n_2614),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2589),
.Y(n_2754)
);

CKINVDCx6p67_ASAP7_75t_R g2755 ( 
.A(n_2607),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2621),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2550),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2594),
.Y(n_2758)
);

AOI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_2489),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2526),
.B(n_507),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2613),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2634),
.Y(n_2762)
);

OAI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2468),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_2763)
);

AOI22xp33_ASAP7_75t_SL g2764 ( 
.A1(n_2468),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2471),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2625),
.A2(n_513),
.B1(n_515),
.B2(n_516),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2634),
.Y(n_2767)
);

INVx3_ASAP7_75t_SL g2768 ( 
.A(n_2545),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_SL g2769 ( 
.A1(n_2614),
.A2(n_518),
.B1(n_520),
.B2(n_521),
.Y(n_2769)
);

OAI22x1_ASAP7_75t_L g2770 ( 
.A1(n_2482),
.A2(n_518),
.B1(n_522),
.B2(n_523),
.Y(n_2770)
);

CKINVDCx11_ASAP7_75t_R g2771 ( 
.A(n_2593),
.Y(n_2771)
);

CKINVDCx8_ASAP7_75t_R g2772 ( 
.A(n_2545),
.Y(n_2772)
);

OAI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2557),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_2773)
);

BUFx12f_ASAP7_75t_L g2774 ( 
.A(n_2588),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2643),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2720),
.B(n_2473),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2643),
.Y(n_2777)
);

BUFx2_ASAP7_75t_SL g2778 ( 
.A(n_2642),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2645),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2645),
.Y(n_2780)
);

OAI21x1_ASAP7_75t_L g2781 ( 
.A1(n_2750),
.A2(n_2477),
.B(n_2479),
.Y(n_2781)
);

OA21x2_ASAP7_75t_L g2782 ( 
.A1(n_2738),
.A2(n_2523),
.B(n_2470),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2772),
.Y(n_2783)
);

BUFx12f_ASAP7_75t_L g2784 ( 
.A(n_2652),
.Y(n_2784)
);

HB1xp67_ASAP7_75t_L g2785 ( 
.A(n_2647),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2720),
.B(n_2726),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2732),
.B(n_2637),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2644),
.A2(n_2641),
.B1(n_2611),
.B2(n_2516),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2748),
.B(n_2619),
.Y(n_2789)
);

BUFx3_ASAP7_75t_L g2790 ( 
.A(n_2665),
.Y(n_2790)
);

OAI21x1_ASAP7_75t_L g2791 ( 
.A1(n_2750),
.A2(n_2485),
.B(n_2487),
.Y(n_2791)
);

OAI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2649),
.A2(n_2637),
.B(n_2534),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2754),
.Y(n_2793)
);

CKINVDCx20_ASAP7_75t_R g2794 ( 
.A(n_2660),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2682),
.B(n_2735),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2648),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2762),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2762),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2747),
.A2(n_2539),
.B1(n_2532),
.B2(n_2639),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2767),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2754),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2655),
.A2(n_2528),
.B1(n_2541),
.B2(n_2488),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2654),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2656),
.Y(n_2804)
);

OA21x2_ASAP7_75t_L g2805 ( 
.A1(n_2757),
.A2(n_2498),
.B(n_2537),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2774),
.A2(n_2675),
.B1(n_2739),
.B2(n_2673),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2679),
.B(n_2488),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2683),
.B(n_2565),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2670),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2676),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2678),
.A2(n_2669),
.B1(n_2691),
.B2(n_2686),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2680),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2652),
.Y(n_2813)
);

OR2x2_ASAP7_75t_L g2814 ( 
.A(n_2728),
.B(n_2700),
.Y(n_2814)
);

OAI21x1_ASAP7_75t_L g2815 ( 
.A1(n_2698),
.A2(n_2492),
.B(n_2525),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2739),
.A2(n_2636),
.B1(n_2566),
.B2(n_2576),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2665),
.Y(n_2817)
);

INVx3_ASAP7_75t_L g2818 ( 
.A(n_2754),
.Y(n_2818)
);

HB1xp67_ASAP7_75t_L g2819 ( 
.A(n_2724),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2734),
.Y(n_2820)
);

INVxp67_ASAP7_75t_L g2821 ( 
.A(n_2706),
.Y(n_2821)
);

AOI22xp33_ASAP7_75t_SL g2822 ( 
.A1(n_2703),
.A2(n_2482),
.B1(n_2632),
.B2(n_2598),
.Y(n_2822)
);

BUFx2_ASAP7_75t_L g2823 ( 
.A(n_2642),
.Y(n_2823)
);

BUFx3_ASAP7_75t_L g2824 ( 
.A(n_2648),
.Y(n_2824)
);

OAI21x1_ASAP7_75t_L g2825 ( 
.A1(n_2677),
.A2(n_2486),
.B(n_2519),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2697),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2742),
.A2(n_2471),
.B1(n_2505),
.B2(n_2500),
.Y(n_2827)
);

OR2x2_ASAP7_75t_L g2828 ( 
.A(n_2667),
.B(n_2581),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2734),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2684),
.B(n_2543),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2742),
.A2(n_2722),
.B1(n_2646),
.B2(n_2714),
.Y(n_2831)
);

AO21x2_ASAP7_75t_L g2832 ( 
.A1(n_2765),
.A2(n_2501),
.B(n_2527),
.Y(n_2832)
);

INVxp67_ASAP7_75t_SL g2833 ( 
.A(n_2718),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2768),
.B(n_2588),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2693),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2723),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2723),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2659),
.B(n_2496),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2677),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2724),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2681),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_L g2842 ( 
.A(n_2725),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2725),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2708),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2666),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2666),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2719),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2666),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2688),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2838),
.B(n_2688),
.Y(n_2850)
);

AOI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2811),
.A2(n_2651),
.B1(n_2650),
.B2(n_2721),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2779),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2838),
.B(n_2688),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2776),
.B(n_2710),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2779),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2821),
.B(n_2741),
.Y(n_2856)
);

A2O1A1Ixp33_ASAP7_75t_L g2857 ( 
.A1(n_2811),
.A2(n_2701),
.B(n_2717),
.C(n_2712),
.Y(n_2857)
);

INVx4_ASAP7_75t_L g2858 ( 
.A(n_2823),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2780),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2776),
.B(n_2740),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2792),
.A2(n_2764),
.B(n_2674),
.Y(n_2861)
);

OAI21x1_ASAP7_75t_L g2862 ( 
.A1(n_2791),
.A2(n_2731),
.B(n_2737),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2786),
.B(n_2722),
.Y(n_2863)
);

INVxp67_ASAP7_75t_L g2864 ( 
.A(n_2823),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2803),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2786),
.B(n_2743),
.Y(n_2866)
);

INVx4_ASAP7_75t_L g2867 ( 
.A(n_2847),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2827),
.A2(n_2671),
.B(n_2769),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2841),
.B(n_2736),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2834),
.B(n_2661),
.Y(n_2870)
);

AND2x4_ASAP7_75t_L g2871 ( 
.A(n_2783),
.B(n_2719),
.Y(n_2871)
);

OAI21x1_ASAP7_75t_SL g2872 ( 
.A1(n_2796),
.A2(n_2746),
.B(n_2702),
.Y(n_2872)
);

AO22x2_ASAP7_75t_L g2873 ( 
.A1(n_2775),
.A2(n_2777),
.B1(n_2828),
.B2(n_2795),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2780),
.Y(n_2874)
);

INVxp67_ASAP7_75t_SL g2875 ( 
.A(n_2847),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2775),
.B(n_2709),
.Y(n_2876)
);

OR2x6_ASAP7_75t_L g2877 ( 
.A(n_2778),
.B(n_2699),
.Y(n_2877)
);

OR2x2_ASAP7_75t_L g2878 ( 
.A(n_2795),
.B(n_2664),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2784),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2814),
.B(n_2689),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2777),
.B(n_2704),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2800),
.B(n_2803),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_SL g2883 ( 
.A(n_2835),
.Y(n_2883)
);

OAI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2827),
.A2(n_2763),
.B(n_2694),
.Y(n_2884)
);

NAND4xp25_ASAP7_75t_L g2885 ( 
.A(n_2831),
.B(n_2685),
.C(n_2658),
.D(n_2695),
.Y(n_2885)
);

AO21x1_ASAP7_75t_L g2886 ( 
.A1(n_2833),
.A2(n_2773),
.B(n_2730),
.Y(n_2886)
);

A2O1A1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2778),
.A2(n_2701),
.B(n_2707),
.C(n_2604),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2800),
.B(n_2771),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2804),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2800),
.B(n_2496),
.Y(n_2890)
);

OR2x2_ASAP7_75t_L g2891 ( 
.A(n_2814),
.B(n_2755),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2788),
.A2(n_2553),
.B(n_2548),
.Y(n_2892)
);

OR2x2_ASAP7_75t_L g2893 ( 
.A(n_2785),
.B(n_2752),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2784),
.B(n_2653),
.Y(n_2894)
);

OA21x2_ASAP7_75t_L g2895 ( 
.A1(n_2791),
.A2(n_2781),
.B(n_2815),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2804),
.Y(n_2896)
);

AO32x2_ASAP7_75t_L g2897 ( 
.A1(n_2796),
.A2(n_2692),
.A3(n_2745),
.B1(n_2729),
.B2(n_2584),
.Y(n_2897)
);

AOI21xp33_ASAP7_75t_L g2898 ( 
.A1(n_2787),
.A2(n_2753),
.B(n_2760),
.Y(n_2898)
);

OAI21x1_ASAP7_75t_L g2899 ( 
.A1(n_2781),
.A2(n_2510),
.B(n_2540),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2809),
.B(n_2744),
.Y(n_2900)
);

OAI22xp5_ASAP7_75t_SL g2901 ( 
.A1(n_2794),
.A2(n_2705),
.B1(n_2672),
.B2(n_2663),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2841),
.B(n_2749),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2809),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2882),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2882),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2873),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2875),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2860),
.B(n_2836),
.Y(n_2908)
);

INVxp67_ASAP7_75t_L g2909 ( 
.A(n_2873),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2860),
.B(n_2836),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2890),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2890),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2858),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2852),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2852),
.Y(n_2915)
);

OR2x2_ASAP7_75t_L g2916 ( 
.A(n_2878),
.B(n_2828),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2873),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2865),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2870),
.B(n_2836),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2889),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2855),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2896),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2858),
.Y(n_2923)
);

HB1xp67_ASAP7_75t_L g2924 ( 
.A(n_2858),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2903),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2855),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2850),
.B(n_2837),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2867),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2859),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2850),
.B(n_2782),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_2851),
.A2(n_2806),
.B1(n_2802),
.B2(n_2799),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2866),
.B(n_2810),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2859),
.Y(n_2933)
);

AOI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2885),
.A2(n_2727),
.B1(n_2789),
.B2(n_2716),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2874),
.Y(n_2935)
);

OR2x2_ASAP7_75t_L g2936 ( 
.A(n_2880),
.B(n_2807),
.Y(n_2936)
);

OR2x2_ASAP7_75t_L g2937 ( 
.A(n_2854),
.B(n_2807),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2853),
.B(n_2782),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2874),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2853),
.B(n_2820),
.Y(n_2940)
);

NOR2xp67_ASAP7_75t_L g2941 ( 
.A(n_2867),
.B(n_2701),
.Y(n_2941)
);

HB1xp67_ASAP7_75t_L g2942 ( 
.A(n_2867),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2866),
.B(n_2782),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2854),
.B(n_2782),
.Y(n_2944)
);

INVx3_ASAP7_75t_L g2945 ( 
.A(n_2913),
.Y(n_2945)
);

NAND3xp33_ASAP7_75t_L g2946 ( 
.A(n_2909),
.B(n_2857),
.C(n_2861),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2932),
.B(n_2881),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2931),
.B(n_2891),
.Y(n_2948)
);

OAI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2931),
.A2(n_2857),
.B(n_2887),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_SL g2950 ( 
.A1(n_2923),
.A2(n_2872),
.B1(n_2703),
.B2(n_2902),
.Y(n_2950)
);

OAI21xp5_ASAP7_75t_SL g2951 ( 
.A1(n_2923),
.A2(n_2887),
.B(n_2868),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2932),
.B(n_2881),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2911),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2936),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2936),
.Y(n_2955)
);

AOI221xp5_ASAP7_75t_L g2956 ( 
.A1(n_2909),
.A2(n_2898),
.B1(n_2884),
.B2(n_2886),
.C(n_2869),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2916),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2916),
.Y(n_2958)
);

BUFx2_ASAP7_75t_L g2959 ( 
.A(n_2924),
.Y(n_2959)
);

NAND3xp33_ASAP7_75t_L g2960 ( 
.A(n_2906),
.B(n_2892),
.C(n_2864),
.Y(n_2960)
);

NAND4xp25_ASAP7_75t_SL g2961 ( 
.A(n_2934),
.B(n_2883),
.C(n_2863),
.D(n_2690),
.Y(n_2961)
);

INVxp67_ASAP7_75t_SL g2962 ( 
.A(n_2924),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2937),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2937),
.Y(n_2964)
);

OAI321xp33_ASAP7_75t_L g2965 ( 
.A1(n_2906),
.A2(n_2877),
.A3(n_2888),
.B1(n_2901),
.B2(n_2856),
.C(n_2894),
.Y(n_2965)
);

HB1xp67_ASAP7_75t_L g2966 ( 
.A(n_2928),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2913),
.B(n_2862),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2943),
.B(n_2863),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2918),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2943),
.B(n_2876),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2913),
.A2(n_2877),
.B1(n_2824),
.B2(n_2819),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2927),
.B(n_2888),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2918),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2904),
.B(n_2893),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2920),
.Y(n_2975)
);

AND2x4_ASAP7_75t_L g2976 ( 
.A(n_2913),
.B(n_2862),
.Y(n_2976)
);

OR2x2_ASAP7_75t_L g2977 ( 
.A(n_2904),
.B(n_2876),
.Y(n_2977)
);

HB1xp67_ASAP7_75t_L g2978 ( 
.A(n_2928),
.Y(n_2978)
);

OAI221xp5_ASAP7_75t_L g2979 ( 
.A1(n_2917),
.A2(n_2879),
.B1(n_2877),
.B2(n_2816),
.C(n_2761),
.Y(n_2979)
);

BUFx2_ASAP7_75t_L g2980 ( 
.A(n_2942),
.Y(n_2980)
);

NOR2x1_ASAP7_75t_R g2981 ( 
.A(n_2940),
.B(n_2813),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2920),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2927),
.B(n_2871),
.Y(n_2983)
);

OAI221xp5_ASAP7_75t_L g2984 ( 
.A1(n_2917),
.A2(n_2877),
.B1(n_2713),
.B2(n_2822),
.C(n_2842),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2942),
.B(n_2871),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2922),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2972),
.B(n_2944),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2969),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2959),
.B(n_2944),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2980),
.B(n_2938),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2973),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2966),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2963),
.B(n_2938),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2975),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2982),
.Y(n_2995)
);

OAI21xp33_ASAP7_75t_SL g2996 ( 
.A1(n_2962),
.A2(n_2941),
.B(n_2907),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2957),
.B(n_2922),
.Y(n_2997)
);

HB1xp67_ASAP7_75t_L g2998 ( 
.A(n_2966),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2964),
.B(n_2930),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2958),
.B(n_2925),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2953),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2953),
.Y(n_3002)
);

AND2x4_ASAP7_75t_L g3003 ( 
.A(n_2967),
.B(n_2930),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2978),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2967),
.B(n_2930),
.Y(n_3005)
);

INVx1_ASAP7_75t_SL g3006 ( 
.A(n_2978),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2986),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2954),
.Y(n_3008)
);

INVx2_ASAP7_75t_SL g3009 ( 
.A(n_2985),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2955),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2997),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_3009),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2997),
.Y(n_3013)
);

INVx1_ASAP7_75t_SL g3014 ( 
.A(n_3006),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_3000),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_3009),
.B(n_2948),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2989),
.B(n_2967),
.Y(n_3017)
);

BUFx2_ASAP7_75t_SL g3018 ( 
.A(n_3006),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_3010),
.B(n_2962),
.Y(n_3019)
);

NAND2x1_ASAP7_75t_L g3020 ( 
.A(n_3003),
.B(n_2945),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_3001),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_3010),
.B(n_2947),
.Y(n_3022)
);

INVxp67_ASAP7_75t_SL g3023 ( 
.A(n_2992),
.Y(n_3023)
);

OR2x2_ASAP7_75t_L g3024 ( 
.A(n_3010),
.B(n_2952),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2989),
.B(n_2976),
.Y(n_3025)
);

OR2x2_ASAP7_75t_L g3026 ( 
.A(n_3008),
.B(n_2974),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_L g3027 ( 
.A(n_2996),
.B(n_2948),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_3000),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2990),
.B(n_2976),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_3008),
.B(n_2968),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2998),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_3001),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_3004),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2988),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2993),
.B(n_2956),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2988),
.Y(n_3036)
);

HB1xp67_ASAP7_75t_L g3037 ( 
.A(n_2991),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_3018),
.B(n_3012),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_3012),
.B(n_3003),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_3016),
.B(n_3003),
.Y(n_3040)
);

INVx3_ASAP7_75t_SL g3041 ( 
.A(n_3014),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_3037),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_3011),
.B(n_2991),
.Y(n_3043)
);

BUFx2_ASAP7_75t_L g3044 ( 
.A(n_3023),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_3031),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_3034),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_3036),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_3016),
.B(n_2946),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_3033),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_3017),
.B(n_3003),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_3027),
.B(n_2844),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_3026),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_3035),
.B(n_3027),
.Y(n_3053)
);

INVx2_ASAP7_75t_SL g3054 ( 
.A(n_3020),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3019),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_3013),
.A2(n_2949),
.B1(n_2984),
.B2(n_3005),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_3041),
.B(n_3022),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_SL g3058 ( 
.A1(n_3051),
.A2(n_2981),
.B(n_2668),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3044),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_3056),
.A2(n_2951),
.B1(n_2996),
.B2(n_2960),
.Y(n_3060)
);

AOI322xp5_ASAP7_75t_L g3061 ( 
.A1(n_3053),
.A2(n_3029),
.A3(n_3025),
.B1(n_3017),
.B2(n_3005),
.C1(n_3015),
.C2(n_3028),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_3041),
.B(n_3025),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_3041),
.B(n_3030),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_3038),
.A2(n_2979),
.B1(n_2961),
.B2(n_3029),
.Y(n_3064)
);

OAI222xp33_ASAP7_75t_L g3065 ( 
.A1(n_3048),
.A2(n_3054),
.B1(n_3045),
.B2(n_3039),
.C1(n_3040),
.C2(n_3052),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_3055),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_3049),
.B(n_3022),
.Y(n_3067)
);

HB1xp67_ASAP7_75t_L g3068 ( 
.A(n_3055),
.Y(n_3068)
);

OAI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_3065),
.A2(n_3049),
.B(n_3042),
.Y(n_3069)
);

OAI21xp33_ASAP7_75t_L g3070 ( 
.A1(n_3060),
.A2(n_3040),
.B(n_3054),
.Y(n_3070)
);

NAND4xp25_ASAP7_75t_L g3071 ( 
.A(n_3064),
.B(n_3050),
.C(n_2950),
.D(n_3047),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_3058),
.A2(n_2965),
.B(n_3046),
.Y(n_3072)
);

NOR2x1p5_ASAP7_75t_SL g3073 ( 
.A(n_3059),
.B(n_3046),
.Y(n_3073)
);

OAI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_3057),
.A2(n_3043),
.B1(n_3050),
.B2(n_3047),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_3068),
.Y(n_3075)
);

AOI322xp5_ASAP7_75t_L g3076 ( 
.A1(n_3062),
.A2(n_3005),
.A3(n_2990),
.B1(n_2999),
.B2(n_2993),
.C1(n_2950),
.C2(n_3032),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_3066),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_3063),
.Y(n_3078)
);

OR2x2_ASAP7_75t_L g3079 ( 
.A(n_3067),
.B(n_3024),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_3075),
.B(n_3061),
.Y(n_3080)
);

OAI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_3078),
.A2(n_3032),
.B(n_3021),
.Y(n_3081)
);

AOI221xp5_ASAP7_75t_L g3082 ( 
.A1(n_3074),
.A2(n_2976),
.B1(n_2907),
.B2(n_2971),
.C(n_3007),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3079),
.Y(n_3083)
);

AOI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_3070),
.A2(n_2657),
.B1(n_2711),
.B2(n_2985),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_3077),
.B(n_2994),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_3069),
.B(n_2994),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3073),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_3071),
.B(n_2995),
.Y(n_3088)
);

NAND3xp33_ASAP7_75t_L g3089 ( 
.A(n_3072),
.B(n_2766),
.C(n_2756),
.Y(n_3089)
);

XOR2x2_ASAP7_75t_L g3090 ( 
.A(n_3076),
.B(n_2985),
.Y(n_3090)
);

A2O1A1Ixp33_ASAP7_75t_SL g3091 ( 
.A1(n_3075),
.A2(n_2945),
.B(n_2759),
.C(n_3001),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_3075),
.B(n_2995),
.Y(n_3092)
);

AOI211x1_ASAP7_75t_L g3093 ( 
.A1(n_3087),
.A2(n_2999),
.B(n_2987),
.C(n_2970),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3083),
.Y(n_3094)
);

OA22x2_ASAP7_75t_L g3095 ( 
.A1(n_3080),
.A2(n_2987),
.B1(n_3002),
.B2(n_2770),
.Y(n_3095)
);

NOR3x1_ASAP7_75t_L g3096 ( 
.A(n_3089),
.B(n_2716),
.C(n_2618),
.Y(n_3096)
);

NOR3xp33_ASAP7_75t_L g3097 ( 
.A(n_3088),
.B(n_2605),
.C(n_2602),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_3084),
.B(n_2662),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3092),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3085),
.Y(n_3100)
);

NAND3xp33_ASAP7_75t_SL g3101 ( 
.A(n_3091),
.B(n_2631),
.C(n_2624),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3081),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_3086),
.B(n_2662),
.Y(n_3103)
);

NAND4xp25_ASAP7_75t_L g3104 ( 
.A(n_3082),
.B(n_2687),
.C(n_2824),
.D(n_2941),
.Y(n_3104)
);

HB1xp67_ASAP7_75t_L g3105 ( 
.A(n_3090),
.Y(n_3105)
);

OAI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_3095),
.A2(n_2696),
.B1(n_3002),
.B2(n_2733),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_3094),
.Y(n_3107)
);

INVxp67_ASAP7_75t_L g3108 ( 
.A(n_3102),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3105),
.B(n_2810),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_R g3110 ( 
.A(n_3098),
.B(n_525),
.Y(n_3110)
);

CKINVDCx16_ASAP7_75t_R g3111 ( 
.A(n_3099),
.Y(n_3111)
);

A2O1A1Ixp33_ASAP7_75t_L g3112 ( 
.A1(n_3103),
.A2(n_2758),
.B(n_2983),
.C(n_2633),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_3093),
.B(n_2812),
.Y(n_3113)
);

AND4x1_ASAP7_75t_L g3114 ( 
.A(n_3096),
.B(n_2715),
.C(n_528),
.D(n_529),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_L g3115 ( 
.A1(n_3101),
.A2(n_3100),
.B1(n_3104),
.B2(n_3097),
.Y(n_3115)
);

AOI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_3111),
.A2(n_2751),
.B1(n_2840),
.B2(n_2843),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_3108),
.A2(n_2940),
.B1(n_2900),
.B2(n_2977),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3107),
.Y(n_3118)
);

AOI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_3106),
.A2(n_2940),
.B1(n_2900),
.B2(n_2905),
.Y(n_3119)
);

AOI221x1_ASAP7_75t_SL g3120 ( 
.A1(n_3109),
.A2(n_3113),
.B1(n_3114),
.B2(n_3115),
.C(n_3112),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3107),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_3108),
.A2(n_2493),
.B(n_2509),
.Y(n_3122)
);

OAI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_3111),
.A2(n_2808),
.B1(n_2783),
.B2(n_2790),
.Y(n_3123)
);

OAI221xp5_ASAP7_75t_L g3124 ( 
.A1(n_3114),
.A2(n_2783),
.B1(n_2790),
.B2(n_2817),
.C(n_2830),
.Y(n_3124)
);

OAI211xp5_ASAP7_75t_L g3125 ( 
.A1(n_3110),
.A2(n_527),
.B(n_528),
.C(n_529),
.Y(n_3125)
);

OAI221xp5_ASAP7_75t_SL g3126 ( 
.A1(n_3114),
.A2(n_2790),
.B1(n_2817),
.B2(n_2908),
.C(n_2910),
.Y(n_3126)
);

OR2x2_ASAP7_75t_L g3127 ( 
.A(n_3118),
.B(n_527),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_3126),
.A2(n_2845),
.B1(n_2849),
.B2(n_2848),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_3121),
.B(n_530),
.Y(n_3129)
);

NOR2x1_ASAP7_75t_L g3130 ( 
.A(n_3125),
.B(n_530),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3116),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_3117),
.B(n_2910),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_3124),
.B(n_534),
.Y(n_3133)
);

NAND4xp75_ASAP7_75t_L g3134 ( 
.A(n_3122),
.B(n_535),
.C(n_536),
.D(n_538),
.Y(n_3134)
);

OR2x2_ASAP7_75t_L g3135 ( 
.A(n_3119),
.B(n_3123),
.Y(n_3135)
);

NAND2x1p5_ASAP7_75t_SL g3136 ( 
.A(n_3120),
.B(n_539),
.Y(n_3136)
);

CKINVDCx16_ASAP7_75t_R g3137 ( 
.A(n_3118),
.Y(n_3137)
);

O2A1O1Ixp33_ASAP7_75t_L g3138 ( 
.A1(n_3127),
.A2(n_3129),
.B(n_3133),
.C(n_3130),
.Y(n_3138)
);

CKINVDCx20_ASAP7_75t_R g3139 ( 
.A(n_3137),
.Y(n_3139)
);

OAI211xp5_ASAP7_75t_SL g3140 ( 
.A1(n_3131),
.A2(n_542),
.B(n_543),
.C(n_544),
.Y(n_3140)
);

XNOR2xp5_ASAP7_75t_L g3141 ( 
.A(n_3136),
.B(n_545),
.Y(n_3141)
);

NOR4xp75_ASAP7_75t_L g3142 ( 
.A(n_3134),
.B(n_547),
.C(n_2908),
.D(n_2919),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3135),
.Y(n_3143)
);

NAND3xp33_ASAP7_75t_SL g3144 ( 
.A(n_3132),
.B(n_2846),
.C(n_2839),
.Y(n_3144)
);

NOR3xp33_ASAP7_75t_L g3145 ( 
.A(n_3128),
.B(n_2554),
.C(n_2547),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3130),
.Y(n_3146)
);

INVx1_ASAP7_75t_SL g3147 ( 
.A(n_3131),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_3139),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_3143),
.B(n_2820),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_SL g3150 ( 
.A1(n_3141),
.A2(n_2911),
.B1(n_2912),
.B2(n_2939),
.Y(n_3150)
);

NAND3xp33_ASAP7_75t_SL g3151 ( 
.A(n_3147),
.B(n_2912),
.C(n_2911),
.Y(n_3151)
);

AND2x4_ASAP7_75t_L g3152 ( 
.A(n_3142),
.B(n_2820),
.Y(n_3152)
);

AOI211xp5_ASAP7_75t_L g3153 ( 
.A1(n_3140),
.A2(n_2926),
.B(n_2929),
.C(n_2912),
.Y(n_3153)
);

BUFx2_ASAP7_75t_L g3154 ( 
.A(n_3146),
.Y(n_3154)
);

AO22x2_ASAP7_75t_L g3155 ( 
.A1(n_3148),
.A2(n_3144),
.B1(n_3138),
.B2(n_3145),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3154),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3149),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3150),
.A2(n_2832),
.B1(n_2895),
.B2(n_2921),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_3152),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_3152),
.Y(n_3160)
);

AOI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_3151),
.A2(n_2832),
.B1(n_2895),
.B2(n_2921),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3153),
.Y(n_3162)
);

INVx1_ASAP7_75t_SL g3163 ( 
.A(n_3156),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_3160),
.B(n_2581),
.Y(n_3164)
);

OAI22xp5_ASAP7_75t_L g3165 ( 
.A1(n_3159),
.A2(n_2933),
.B1(n_2921),
.B2(n_2915),
.Y(n_3165)
);

AOI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_3157),
.A2(n_2935),
.B1(n_2933),
.B2(n_2915),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_3162),
.Y(n_3167)
);

OAI22x1_ASAP7_75t_L g3168 ( 
.A1(n_3158),
.A2(n_2933),
.B1(n_2915),
.B2(n_2914),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_3163),
.B(n_3155),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_3167),
.B(n_3161),
.Y(n_3170)
);

OAI22xp5_ASAP7_75t_SL g3171 ( 
.A1(n_3164),
.A2(n_2914),
.B1(n_2826),
.B2(n_2897),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3168),
.B(n_2581),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_3169),
.A2(n_3166),
.B1(n_3165),
.B2(n_2818),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_3170),
.A2(n_2801),
.B1(n_2818),
.B2(n_2793),
.Y(n_3174)
);

OA21x2_ASAP7_75t_L g3175 ( 
.A1(n_3172),
.A2(n_2899),
.B(n_2825),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3173),
.A2(n_3171),
.B1(n_2801),
.B2(n_2818),
.Y(n_3176)
);

OAI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_3176),
.A2(n_3174),
.B(n_3175),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3177),
.Y(n_3178)
);

OAI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_3177),
.A2(n_2793),
.B1(n_2801),
.B2(n_2829),
.Y(n_3179)
);

OAI221xp5_ASAP7_75t_R g3180 ( 
.A1(n_3178),
.A2(n_2897),
.B1(n_2826),
.B2(n_2805),
.C(n_2793),
.Y(n_3180)
);

AOI211xp5_ASAP7_75t_L g3181 ( 
.A1(n_3180),
.A2(n_3179),
.B(n_2798),
.C(n_2797),
.Y(n_3181)
);


endmodule