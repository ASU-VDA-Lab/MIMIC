module fake_netlist_1_12055_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_7), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_11), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AND3x1_ASAP7_75t_L g20 ( .A(n_18), .B(n_0), .C(n_1), .Y(n_20) );
AO22x2_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_17), .B1(n_16), .B2(n_1), .Y(n_21) );
AOI33xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .A3(n_20), .B1(n_15), .B2(n_14), .B3(n_13), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_2), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_25), .B(n_3), .C(n_8), .Y(n_26) );
INVx1_ASAP7_75t_SL g27 ( .A(n_26), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_28) );
endmodule