module fake_netlist_6_729_n_772 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_772);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_772;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_21),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_13),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_88),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_57),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_24),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_64),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_31),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_32),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_60),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_34),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_19),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_4),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_18),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_37),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_84),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_33),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_4),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_48),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_49),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_44),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_10),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_23),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_61),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_27),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_151),
.B(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_159),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_162),
.B(n_157),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_2),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_153),
.B(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_154),
.B(n_5),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_6),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_171),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_7),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_8),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_9),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_221),
.Y(n_254)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_207),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_201),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_204),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_216),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_10),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_208),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_R g266 ( 
.A(n_225),
.B(n_152),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_236),
.B(n_194),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_218),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_236),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_155),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_237),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_237),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_212),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_212),
.Y(n_289)
);

NOR2x1p5_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_244),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_231),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_258),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_224),
.C(n_223),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_213),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_241),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_244),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

BUFx6f_ASAP7_75t_SL g310 ( 
.A(n_253),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_267),
.B(n_156),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_260),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_239),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_213),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_276),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_224),
.C(n_223),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_245),
.C(n_233),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_239),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_279),
.B(n_245),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_274),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_262),
.B(n_282),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_266),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_158),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_255),
.B(n_160),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_239),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_243),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_213),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_259),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_161),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_251),
.B(n_164),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_243),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_243),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_252),
.B(n_166),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_195),
.C(n_175),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_254),
.B(n_243),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_256),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_273),
.B(n_246),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_248),
.B(n_173),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_246),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_267),
.B(n_180),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_247),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_181),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_246),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_210),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_317),
.B(n_186),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_298),
.A2(n_210),
.B1(n_188),
.B2(n_189),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_308),
.B(n_203),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_302),
.A2(n_200),
.B1(n_196),
.B2(n_192),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_335),
.B(n_203),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_221),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_11),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_312),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_17),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_20),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_307),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_347),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_315),
.B(n_347),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_356),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_311),
.A2(n_82),
.B1(n_144),
.B2(n_142),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

BUFx4f_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_318),
.B(n_12),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_301),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_352),
.A2(n_81),
.B1(n_141),
.B2(n_140),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_22),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_26),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_297),
.Y(n_399)
);

NOR2x2_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_14),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_309),
.Y(n_401)
);

BUFx4f_ASAP7_75t_L g402 ( 
.A(n_297),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_15),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_299),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_303),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_331),
.A2(n_86),
.B(n_28),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_326),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_328),
.B(n_29),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_330),
.A2(n_87),
.B(n_30),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_310),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_35),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_310),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_339),
.B(n_16),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_370),
.B(n_378),
.C(n_381),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_327),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_377),
.A2(n_357),
.B1(n_344),
.B2(n_337),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_343),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_403),
.B(n_357),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_306),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_345),
.B(n_350),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_345),
.B(n_350),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_336),
.Y(n_434)
);

OAI22x1_ASAP7_75t_L g435 ( 
.A1(n_374),
.A2(n_417),
.B1(n_414),
.B2(n_408),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_350),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_380),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_373),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_372),
.B(n_353),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_359),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_419),
.A2(n_353),
.B1(n_39),
.B2(n_40),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_353),
.B(n_41),
.C(n_42),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_387),
.B(n_38),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_387),
.B(n_45),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_46),
.B(n_47),
.C(n_50),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_415),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_54),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_386),
.B(n_55),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_56),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_400),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_375),
.A2(n_58),
.B(n_59),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_366),
.B(n_401),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_394),
.A2(n_62),
.B(n_63),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_376),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_398),
.A2(n_65),
.B(n_66),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_67),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_395),
.B(n_68),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_358),
.B(n_69),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_70),
.B(n_71),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

BUFx2_ASAP7_75t_SL g468 ( 
.A(n_405),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_421),
.A2(n_73),
.B(n_74),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_420),
.B(n_77),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_409),
.A2(n_79),
.B(n_83),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_358),
.B(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_406),
.B(n_89),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_410),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_363),
.A2(n_393),
.B1(n_383),
.B2(n_392),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_365),
.B(n_90),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

AO21x1_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_407),
.B(n_369),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_446),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_424),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_452),
.A2(n_399),
.B(n_418),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_474),
.A2(n_365),
.B(n_399),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_428),
.B(n_365),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_431),
.A2(n_91),
.B(n_94),
.Y(n_489)
);

AO21x2_ASAP7_75t_L g490 ( 
.A1(n_445),
.A2(n_96),
.B(n_97),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_426),
.B(n_149),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_432),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g494 ( 
.A(n_470),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

AOI22x1_ASAP7_75t_L g496 ( 
.A1(n_460),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_433),
.A2(n_105),
.B(n_107),
.Y(n_499)
);

OAI21x1_ASAP7_75t_SL g500 ( 
.A1(n_453),
.A2(n_108),
.B(n_109),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_423),
.B(n_422),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_454),
.A2(n_110),
.B(n_112),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_456),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_462),
.A2(n_139),
.B(n_116),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

NAND2x1p5_ASAP7_75t_L g511 ( 
.A(n_448),
.B(n_449),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_114),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_463),
.A2(n_117),
.B(n_118),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_434),
.A2(n_119),
.B(n_120),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_471),
.A2(n_436),
.B(n_478),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_121),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_461),
.A2(n_457),
.B(n_459),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_464),
.B(n_138),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_472),
.A2(n_123),
.B(n_124),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_466),
.A2(n_125),
.B(n_127),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_469),
.A2(n_129),
.B(n_132),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_476),
.B1(n_458),
.B2(n_472),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_467),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_521),
.A2(n_476),
.B1(n_442),
.B2(n_473),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_495),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_492),
.Y(n_529)
);

BUFx8_ASAP7_75t_SL g530 ( 
.A(n_494),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_491),
.B(n_475),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_494),
.Y(n_532)
);

OA21x2_ASAP7_75t_L g533 ( 
.A1(n_485),
.A2(n_451),
.B(n_450),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_483),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_427),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_497),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_492),
.Y(n_538)
);

BUFx8_ASAP7_75t_L g539 ( 
.A(n_522),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_491),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_492),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_516),
.A2(n_425),
.B1(n_522),
.B2(n_507),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_498),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_479),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_488),
.B(n_470),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_480),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_471),
.Y(n_549)
);

BUFx2_ASAP7_75t_R g550 ( 
.A(n_490),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_492),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_443),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_508),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_508),
.Y(n_559)
);

INVx8_ASAP7_75t_L g560 ( 
.A(n_495),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_489),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_510),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_485),
.A2(n_133),
.B(n_134),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_530),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_547),
.B(n_502),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_560),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_547),
.B(n_518),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_528),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_528),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_R g572 ( 
.A(n_536),
.B(n_488),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_525),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_532),
.B(n_507),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_524),
.B(n_511),
.Y(n_576)
);

AO31x2_ASAP7_75t_L g577 ( 
.A1(n_526),
.A2(n_481),
.A3(n_484),
.B(n_505),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_536),
.B(n_507),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_541),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_559),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_546),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_546),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_560),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_539),
.A2(n_519),
.B1(n_496),
.B2(n_509),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_559),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_531),
.B(n_511),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_548),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_518),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_527),
.B(n_504),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_541),
.B(n_560),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_548),
.B(n_487),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_543),
.A2(n_496),
.B1(n_509),
.B2(n_503),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_557),
.B(n_486),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_535),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g600 ( 
.A(n_555),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_527),
.B(n_504),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_544),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_SL g605 ( 
.A1(n_539),
.A2(n_511),
.B1(n_490),
.B2(n_512),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_539),
.A2(n_490),
.B1(n_512),
.B2(n_500),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_R g607 ( 
.A(n_532),
.B(n_495),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_545),
.B(n_487),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_564),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_554),
.B(n_505),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_553),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_579),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_584),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_573),
.B(n_556),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_569),
.B(n_563),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_590),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_591),
.B(n_550),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_515),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_599),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_599),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_578),
.B(n_552),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_609),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_612),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_612),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_610),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_589),
.B(n_515),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_583),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_596),
.B(n_533),
.C(n_565),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_589),
.B(n_515),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_594),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_585),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_610),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_565),
.Y(n_638)
);

OAI221xp5_ASAP7_75t_L g639 ( 
.A1(n_596),
.A2(n_512),
.B1(n_468),
.B2(n_549),
.C(n_533),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_578),
.B(n_565),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_562),
.Y(n_641)
);

NOR2x1_ASAP7_75t_SL g642 ( 
.A(n_576),
.B(n_542),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_588),
.B(n_562),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_598),
.B(n_562),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_597),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_567),
.B(n_561),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_604),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_628),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_628),
.B(n_582),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_627),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_627),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_631),
.B(n_577),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_631),
.B(n_623),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_625),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_629),
.B(n_577),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_634),
.B(n_577),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_616),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_645),
.B(n_567),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_644),
.B(n_608),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_635),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_622),
.B(n_587),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_645),
.B(n_605),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_623),
.B(n_605),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_625),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_634),
.B(n_606),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_608),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_622),
.B(n_587),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_637),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_640),
.B(n_594),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_621),
.B(n_600),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_620),
.B(n_606),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_621),
.B(n_592),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_637),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_651),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_652),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_654),
.B(n_647),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_655),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_619),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_672),
.B(n_641),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_654),
.B(n_647),
.Y(n_683)
);

NAND4xp25_ASAP7_75t_L g684 ( 
.A(n_663),
.B(n_620),
.C(n_624),
.D(n_619),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_667),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_666),
.B(n_640),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_665),
.B(n_641),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_671),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_672),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_649),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_676),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_650),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_672),
.B(n_642),
.Y(n_693)
);

NOR3xp33_ASAP7_75t_SL g694 ( 
.A(n_670),
.B(n_639),
.C(n_572),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_673),
.Y(n_695)
);

AOI32xp33_ASAP7_75t_L g696 ( 
.A1(n_686),
.A2(n_663),
.A3(n_670),
.B1(n_674),
.B2(n_668),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_686),
.B(n_668),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_674),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_679),
.B(n_672),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_693),
.B(n_669),
.Y(n_700)
);

OAI322xp33_ASAP7_75t_L g701 ( 
.A1(n_695),
.A2(n_660),
.A3(n_657),
.B1(n_656),
.B2(n_630),
.C1(n_662),
.C2(n_664),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_690),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_690),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_677),
.Y(n_704)
);

OAI33xp33_ASAP7_75t_L g705 ( 
.A1(n_681),
.A2(n_675),
.A3(n_643),
.B1(n_664),
.B2(n_662),
.B3(n_646),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_678),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_683),
.B(n_666),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_703),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_698),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_700),
.A2(n_694),
.B(n_684),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_702),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_705),
.A2(n_693),
.B1(n_694),
.B2(n_682),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_699),
.B(n_687),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_709),
.B(n_696),
.Y(n_714)
);

AOI211xp5_ASAP7_75t_L g715 ( 
.A1(n_710),
.A2(n_701),
.B(n_693),
.C(n_706),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_710),
.A2(n_712),
.B1(n_689),
.B2(n_682),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_708),
.A2(n_697),
.B1(n_689),
.B2(n_707),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_711),
.A2(n_701),
.B1(n_704),
.B2(n_691),
.C(n_688),
.Y(n_718)
);

OAI21xp33_ASAP7_75t_L g719 ( 
.A1(n_716),
.A2(n_689),
.B(n_659),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_715),
.A2(n_714),
.B1(n_718),
.B2(n_717),
.Y(n_720)
);

AND3x1_ASAP7_75t_L g721 ( 
.A(n_715),
.B(n_713),
.C(n_566),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_714),
.B(n_580),
.C(n_592),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_722),
.A2(n_685),
.B1(n_680),
.B2(n_682),
.Y(n_723)
);

AO22x2_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_633),
.B1(n_643),
.B2(n_614),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_SL g725 ( 
.A1(n_724),
.A2(n_720),
.B(n_719),
.C(n_530),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_723),
.A2(n_661),
.B1(n_653),
.B2(n_635),
.Y(n_726)
);

NAND5xp2_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_575),
.C(n_653),
.D(n_607),
.E(n_513),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_727),
.B(n_725),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_726),
.A2(n_635),
.B1(n_614),
.B2(n_594),
.Y(n_731)
);

NOR2x1_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_502),
.Y(n_732)
);

NOR2x1_ASAP7_75t_L g733 ( 
.A(n_727),
.B(n_593),
.Y(n_733)
);

AND3x4_ASAP7_75t_L g734 ( 
.A(n_725),
.B(n_626),
.C(n_601),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_580),
.C(n_513),
.Y(n_735)
);

XNOR2xp5_ASAP7_75t_L g736 ( 
.A(n_734),
.B(n_601),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_729),
.A2(n_635),
.B1(n_626),
.B2(n_638),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_732),
.Y(n_738)
);

XNOR2xp5_ASAP7_75t_L g739 ( 
.A(n_730),
.B(n_593),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_SL g740 ( 
.A1(n_731),
.A2(n_618),
.B(n_615),
.C(n_529),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_738),
.B(n_733),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_R g742 ( 
.A(n_739),
.B(n_555),
.Y(n_742)
);

OAI21xp33_ASAP7_75t_SL g743 ( 
.A1(n_737),
.A2(n_523),
.B(n_520),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_736),
.B(n_495),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_740),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_741),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

XNOR2xp5_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_735),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_742),
.Y(n_749)
);

AND4x1_ASAP7_75t_L g750 ( 
.A(n_743),
.B(n_136),
.C(n_137),
.D(n_555),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_741),
.A2(n_500),
.B1(n_581),
.B2(n_482),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_741),
.Y(n_752)
);

OA22x2_ASAP7_75t_L g753 ( 
.A1(n_741),
.A2(n_581),
.B1(n_615),
.B2(n_618),
.Y(n_753)
);

NOR2x1_ASAP7_75t_L g754 ( 
.A(n_752),
.B(n_495),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_746),
.A2(n_749),
.B1(n_748),
.B2(n_747),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_753),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_751),
.A2(n_568),
.B1(n_602),
.B2(n_586),
.Y(n_757)
);

OAI31xp33_ASAP7_75t_L g758 ( 
.A1(n_750),
.A2(n_549),
.A3(n_482),
.B(n_552),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_752),
.A2(n_568),
.B1(n_602),
.B2(n_586),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_752),
.A2(n_568),
.B1(n_602),
.B2(n_586),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_752),
.A2(n_635),
.B1(n_626),
.B2(n_636),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_642),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_754),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_758),
.A2(n_517),
.B(n_523),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_756),
.B(n_648),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_759),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_761),
.B1(n_760),
.B2(n_757),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_763),
.A2(n_542),
.B1(n_552),
.B2(n_538),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_767),
.B(n_762),
.C(n_765),
.Y(n_769)
);

AOI322xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_768),
.A3(n_764),
.B1(n_538),
.B2(n_529),
.C1(n_638),
.C2(n_632),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_770),
.B(n_538),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_514),
.B1(n_542),
.B2(n_499),
.Y(n_772)
);


endmodule