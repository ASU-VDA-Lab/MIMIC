module real_jpeg_16040_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_71, n_7, n_3, n_5, n_4, n_70, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_71;
input n_7;
input n_3;
input n_5;
input n_4;
input n_70;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_58;
wire n_52;
wire n_31;
wire n_49;
wire n_67;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_51;
wire n_45;
wire n_61;
wire n_47;
wire n_25;
wire n_42;
wire n_22;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_32;
wire n_30;

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_13),
.C(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_71),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_28),
.B(n_31),
.Y(n_27)
);

AOI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_50),
.B1(n_58),
.B2(n_61),
.C(n_68),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_20),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_34),
.B2(n_42),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_22),
.A2(n_34),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_24),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_33),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_66),
.Y(n_68)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_62),
.B(n_67),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_70),
.Y(n_29)
);


endmodule