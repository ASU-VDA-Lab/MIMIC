module fake_jpeg_27353_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_8),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_59),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_34),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_34),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_64),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_30),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_32),
.Y(n_92)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_19),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_77)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_67),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_16),
.C(n_27),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_40),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_89),
.B(n_96),
.Y(n_122)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_87),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_46),
.B1(n_56),
.B2(n_64),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_37),
.B1(n_18),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_99),
.B1(n_24),
.B2(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_42),
.A3(n_18),
.B1(n_32),
.B2(n_43),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_42),
.C(n_18),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_100),
.B1(n_103),
.B2(n_46),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_17),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_40),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

OR2x4_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_83),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_123),
.B1(n_81),
.B2(n_100),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_128),
.B1(n_131),
.B2(n_77),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_96),
.B(n_78),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_124),
.Y(n_133)
);

FAx1_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_79),
.CI(n_69),
.CON(n_120),
.SN(n_120)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_83),
.CI(n_87),
.CON(n_143),
.SN(n_143)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_56),
.B1(n_18),
.B2(n_28),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_39),
.C(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_89),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_135),
.B(n_142),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_143),
.B(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_71),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_81),
.B1(n_75),
.B2(n_74),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_155),
.B1(n_160),
.B2(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_90),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_58),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_94),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_73),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_152),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_73),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_76),
.B1(n_70),
.B2(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_70),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_13),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_76),
.B1(n_39),
.B2(n_16),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_51),
.B1(n_28),
.B2(n_27),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_29),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_51),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_122),
.C(n_115),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_189),
.C(n_170),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_120),
.C(n_126),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_174),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_120),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_118),
.B(n_120),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_177),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_132),
.B1(n_127),
.B2(n_111),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_190),
.B1(n_147),
.B2(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_112),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_188),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_132),
.B(n_112),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_107),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_131),
.C(n_107),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_133),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_156),
.Y(n_216)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_39),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_161),
.B(n_155),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_159),
.C(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_221),
.C(n_223),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_210),
.B1(n_196),
.B2(n_178),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_173),
.B(n_178),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_165),
.B1(n_181),
.B2(n_182),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_196),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_167),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_136),
.B1(n_143),
.B2(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_215),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_136),
.B(n_154),
.Y(n_213)
);

BUFx12f_ASAP7_75t_SL g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_168),
.B(n_142),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_191),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_39),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_194),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_218),
.B(n_207),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_242),
.B(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_165),
.B1(n_197),
.B2(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_234),
.B1(n_244),
.B2(n_245),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_197),
.B1(n_189),
.B2(n_190),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_176),
.C(n_195),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_246),
.C(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_215),
.B1(n_210),
.B2(n_220),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_201),
.Y(n_241)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_199),
.A2(n_173),
.B(n_166),
.C(n_151),
.Y(n_244)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_202),
.A2(n_191),
.B1(n_166),
.B2(n_29),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_39),
.C(n_58),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_231),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_252),
.B1(n_227),
.B2(n_232),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_200),
.B1(n_206),
.B2(n_224),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_222),
.C(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_214),
.C(n_221),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_200),
.C(n_211),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_217),
.B(n_203),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_244),
.B(n_10),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_201),
.C(n_29),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_244),
.C(n_2),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_242),
.B1(n_245),
.B2(n_232),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_9),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_7),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_9),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_270),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_276),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_237),
.B(n_229),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_256),
.B(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_242),
.B1(n_241),
.B2(n_231),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_241),
.B1(n_244),
.B2(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_249),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_282),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_265),
.B1(n_256),
.B2(n_266),
.C(n_251),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_277),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_261),
.C(n_264),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_287),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_282),
.B(n_278),
.Y(n_300)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_276),
.B1(n_271),
.B2(n_250),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_296),
.A2(n_300),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_12),
.C2(n_0),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_251),
.B1(n_279),
.B2(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_302),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_260),
.B1(n_259),
.B2(n_4),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_7),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_290),
.C(n_294),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_11),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_285),
.C(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_294),
.Y(n_309)
);

AOI31xp33_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_11),
.A3(n_14),
.B(n_13),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_312),
.B1(n_301),
.B2(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_299),
.Y(n_316)
);

AOI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_310),
.A3(n_307),
.B1(n_309),
.B2(n_304),
.C(n_302),
.Y(n_317)
);

OAI31xp33_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_307),
.A3(n_313),
.B(n_15),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_318),
.C2(n_311),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_5),
.Y(n_322)
);


endmodule