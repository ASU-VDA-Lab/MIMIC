module fake_jpeg_330_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx13_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_5),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_8),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_10),
.B(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_12),
.C(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_20),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_27),
.B(n_6),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_9),
.B1(n_6),
.B2(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_26),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_9),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_6),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_6),
.B(n_3),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_35),
.CI(n_3),
.CON(n_38),
.SN(n_38)
);

AOI311xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_2),
.A3(n_4),
.B(n_31),
.C(n_29),
.Y(n_39)
);


endmodule