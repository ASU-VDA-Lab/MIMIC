module fake_jpeg_1295_n_531 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_1),
.B(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_55),
.B(n_61),
.Y(n_121)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_70),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_18),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_71),
.A2(n_52),
.B1(n_17),
.B2(n_45),
.Y(n_148)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_79),
.B(n_103),
.Y(n_175)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_40),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_7),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_7),
.B(n_14),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_0),
.B(n_1),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_92),
.B(n_99),
.Y(n_159)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_22),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_109),
.Y(n_172)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_48),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_46),
.B1(n_36),
.B2(n_25),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_148),
.B1(n_52),
.B2(n_45),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_117),
.B(n_132),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_17),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_118),
.B(n_124),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_40),
.C(n_38),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_126),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_26),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_53),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_145),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_26),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_68),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_174),
.Y(n_186)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_57),
.B(n_31),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_126),
.A2(n_106),
.B1(n_100),
.B2(n_98),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_176),
.A2(n_183),
.B1(n_187),
.B2(n_220),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_84),
.B(n_101),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_178),
.A2(n_146),
.B(n_152),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_113),
.A2(n_60),
.B1(n_65),
.B2(n_94),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_184),
.B(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_54),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_212),
.Y(n_245)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_91),
.B1(n_89),
.B2(n_67),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_196),
.A2(n_214),
.B1(n_33),
.B2(n_146),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_150),
.A2(n_81),
.B1(n_21),
.B2(n_31),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_224),
.B1(n_226),
.B2(n_228),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_48),
.B1(n_47),
.B2(n_69),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_33),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_33),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_54),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_221),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_150),
.A2(n_70),
.B1(n_96),
.B2(n_28),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_121),
.B(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_114),
.B(n_58),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_225),
.Y(n_259)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_168),
.A2(n_21),
.B1(n_31),
.B2(n_49),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_119),
.B(n_75),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_22),
.B1(n_28),
.B2(n_47),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_153),
.A2(n_49),
.B(n_44),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_178),
.C(n_179),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g230 ( 
.A1(n_176),
.A2(n_97),
.B1(n_154),
.B2(n_151),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_240),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_238),
.B(n_208),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_166),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_249),
.A2(n_194),
.B1(n_207),
.B2(n_21),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_128),
.C(n_122),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_198),
.B(n_144),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_141),
.Y(n_255)
);

OAI22x1_ASAP7_75t_SL g258 ( 
.A1(n_187),
.A2(n_168),
.B1(n_115),
.B2(n_135),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_200),
.B1(n_197),
.B2(n_212),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_202),
.B(n_140),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_112),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_208),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_259),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_188),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_272),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_196),
.B1(n_204),
.B2(n_217),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_289),
.B1(n_296),
.B2(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_183),
.B1(n_182),
.B2(n_205),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_184),
.C(n_227),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_280),
.C(n_243),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_186),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_283),
.Y(n_325)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_185),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_234),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_206),
.C(n_203),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_209),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_240),
.B(n_216),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_286),
.Y(n_317)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_215),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_230),
.A2(n_210),
.B1(n_219),
.B2(n_189),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_233),
.B(n_262),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_237),
.A2(n_163),
.B1(n_211),
.B2(n_157),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_193),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_292),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_160),
.B1(n_201),
.B2(n_156),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_294),
.B1(n_199),
.B2(n_232),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_193),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_195),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_298),
.B(n_263),
.C(n_231),
.D(n_243),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_242),
.A2(n_200),
.B1(n_197),
.B2(n_163),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_233),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_195),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_228),
.B1(n_116),
.B2(n_190),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_305),
.C(n_313),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_230),
.B1(n_249),
.B2(n_252),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_304),
.A2(n_283),
.B1(n_287),
.B2(n_293),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_260),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_244),
.B(n_235),
.C(n_257),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_308),
.B(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_284),
.Y(n_343)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_232),
.B1(n_256),
.B2(n_253),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_288),
.B1(n_299),
.B2(n_286),
.Y(n_341)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_320),
.A2(n_327),
.B(n_329),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_324),
.B1(n_297),
.B2(n_292),
.Y(n_347)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_239),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_326),
.B(n_298),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_267),
.B(n_262),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_246),
.B(n_250),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_329),
.B(n_294),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_276),
.A2(n_246),
.B(n_250),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_341),
.B1(n_347),
.B2(n_323),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_313),
.B(n_273),
.CI(n_278),
.CON(n_331),
.SN(n_331)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_331),
.B(n_332),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_349),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_340),
.B(n_342),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_312),
.A2(n_272),
.B1(n_291),
.B2(n_296),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_345),
.B1(n_357),
.B2(n_304),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_289),
.B(n_275),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_343),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_302),
.A2(n_272),
.B1(n_288),
.B2(n_297),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_326),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_280),
.Y(n_351)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_321),
.A2(n_277),
.B(n_297),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_355),
.A2(n_308),
.B(n_318),
.Y(n_373)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_302),
.A2(n_272),
.B1(n_297),
.B2(n_277),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_273),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_309),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_305),
.C(n_301),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_364),
.C(n_365),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_369),
.B1(n_345),
.B2(n_357),
.Y(n_394)
);

OAI32xp33_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_318),
.A3(n_317),
.B1(n_325),
.B2(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_177),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_307),
.C(n_327),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_325),
.C(n_274),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_342),
.A2(n_316),
.B1(n_320),
.B2(n_328),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_370),
.B(n_384),
.Y(n_401)
);

AOI21xp33_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_49),
.B(n_44),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_385),
.B1(n_330),
.B2(n_347),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_332),
.B(n_311),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_377),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_322),
.C(n_300),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_382),
.C(n_386),
.Y(n_417)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_381),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_300),
.C(n_263),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_352),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_345),
.B1(n_339),
.B2(n_341),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_231),
.C(n_191),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_256),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_387),
.B(n_335),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_275),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_331),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_360),
.A2(n_334),
.B(n_355),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_397),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_333),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_395),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_402),
.B1(n_404),
.B2(n_406),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_331),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_396),
.A2(n_399),
.B1(n_410),
.B2(n_369),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_360),
.A2(n_340),
.B(n_330),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_409),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_385),
.A2(n_339),
.B1(n_353),
.B2(n_350),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_361),
.A2(n_356),
.B1(n_348),
.B2(n_336),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_374),
.A2(n_336),
.B1(n_335),
.B2(n_344),
.Y(n_404)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_344),
.B(n_223),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_253),
.B(n_191),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_408),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_366),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_373),
.A2(n_181),
.B1(n_180),
.B2(n_116),
.Y(n_410)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_412),
.Y(n_432)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_413),
.B(n_415),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_36),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_414),
.Y(n_436)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_28),
.B1(n_44),
.B2(n_36),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_416),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_394),
.A2(n_372),
.B1(n_377),
.B2(n_379),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_392),
.B1(n_404),
.B2(n_410),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_401),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_422),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_382),
.C(n_372),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_434),
.B1(n_130),
.B2(n_125),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_379),
.C(n_364),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_428),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_386),
.C(n_371),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_371),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_433),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_363),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_399),
.A2(n_380),
.B1(n_376),
.B2(n_368),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_407),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_15),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_411),
.B(n_376),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_437),
.B(n_415),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_380),
.C(n_152),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_428),
.C(n_423),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_398),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_419),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_414),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_453),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_408),
.B(n_412),
.C(n_390),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_452),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_406),
.B(n_397),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_451),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_448),
.A2(n_421),
.B1(n_436),
.B2(n_434),
.Y(n_465)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

INVx13_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_392),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_400),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_440),
.A2(n_389),
.B(n_403),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_457),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_441),
.B(n_418),
.C(n_423),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_424),
.A2(n_413),
.B1(n_389),
.B2(n_130),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_458),
.B(n_125),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_461),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_468),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_443),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_433),
.B1(n_419),
.B2(n_430),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_425),
.C(n_439),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_477),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_425),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_453),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_456),
.A2(n_130),
.B1(n_125),
.B2(n_111),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_476),
.B(n_478),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_457),
.A2(n_111),
.B1(n_46),
.B2(n_36),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_467),
.A2(n_449),
.B(n_459),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_484),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_483),
.B(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_444),
.C(n_446),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_470),
.B(n_462),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_458),
.Y(n_487)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_487),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

NOR2x1_ASAP7_75t_R g489 ( 
.A(n_468),
.B(n_452),
.Y(n_489)
);

AOI31xp67_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_11),
.A3(n_15),
.B(n_12),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_473),
.A2(n_452),
.B(n_455),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_490),
.A2(n_494),
.B(n_493),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_474),
.B(n_451),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_492),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_46),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_467),
.A2(n_464),
.B(n_475),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_480),
.A2(n_472),
.B(n_475),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_498),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_466),
.C(n_478),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_501),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_46),
.C(n_41),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_504),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_490),
.A2(n_39),
.B(n_10),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_482),
.A2(n_39),
.B1(n_41),
.B2(n_10),
.Y(n_505)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_489),
.A3(n_481),
.B1(n_39),
.B2(n_41),
.C1(n_16),
.C2(n_9),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_514),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_16),
.C(n_6),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_507),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_515),
.A2(n_505),
.B(n_501),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_496),
.B(n_6),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_516),
.B(n_1),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_517),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_513),
.C(n_500),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_SL g523 ( 
.A(n_519),
.B(n_521),
.C(n_522),
.Y(n_523)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g520 ( 
.A1(n_513),
.A2(n_499),
.B(n_498),
.C(n_506),
.D(n_503),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_511),
.A3(n_508),
.B1(n_515),
.B2(n_3),
.C1(n_1),
.C2(n_4),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_16),
.B(n_2),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_3),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_518),
.C(n_3),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_526),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_528),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_523),
.Y(n_531)
);


endmodule