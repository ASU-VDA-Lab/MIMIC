module fake_jpeg_19602_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_5),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_12),
.B1(n_9),
.B2(n_13),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_15),
.A2(n_18),
.B1(n_9),
.B2(n_4),
.Y(n_27)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_22),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_3),
.B1(n_4),
.B2(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_24),
.B1(n_15),
.B2(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.C(n_26),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_17),
.B1(n_22),
.B2(n_16),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_33),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_32),
.C(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_30),
.B(n_31),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_40),
.B1(n_37),
.B2(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.C(n_44),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_38),
.A3(n_28),
.B1(n_25),
.B2(n_10),
.C1(n_14),
.C2(n_16),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_10),
.B1(n_14),
.B2(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_4),
.Y(n_49)
);


endmodule