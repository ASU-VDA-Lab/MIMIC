module fake_jpeg_16836_n_396 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_43),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_7),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_7),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_6),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_40),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_79),
.B1(n_84),
.B2(n_90),
.Y(n_141)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_83),
.Y(n_122)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_30),
.B(n_31),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_31),
.C(n_2),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_32),
.B1(n_20),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_91),
.B1(n_4),
.B2(n_9),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_79)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_9),
.B1(n_12),
.B2(n_3),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_30),
.B1(n_36),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_15),
.B1(n_33),
.B2(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_96),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_37),
.B1(n_27),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_103),
.B1(n_31),
.B2(n_29),
.Y(n_142)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_35),
.B1(n_16),
.B2(n_25),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_105),
.Y(n_166)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_16),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_118),
.Y(n_137)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_44),
.B1(n_54),
.B2(n_57),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_123),
.A2(n_159),
.B1(n_161),
.B2(n_72),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_134),
.Y(n_181)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_133),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_48),
.B1(n_39),
.B2(n_30),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_170),
.B1(n_148),
.B2(n_135),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_25),
.B(n_42),
.C(n_30),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_144),
.Y(n_186)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_88),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_10),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_135),
.A2(n_148),
.B(n_2),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_73),
.A2(n_29),
.B1(n_14),
.B2(n_31),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_147),
.B1(n_163),
.B2(n_93),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_87),
.B(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_142),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_67),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_150),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_9),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_91),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_154),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_81),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_84),
.B(n_31),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_82),
.A2(n_113),
.A3(n_112),
.B1(n_77),
.B2(n_102),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_165),
.B(n_94),
.C(n_10),
.Y(n_184)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_5),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_104),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_160),
.B(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_76),
.B1(n_113),
.B2(n_82),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_115),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_71),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_5),
.B1(n_10),
.B2(n_3),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_4),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_167),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_115),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_172),
.A2(n_189),
.B1(n_204),
.B2(n_194),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_173),
.A2(n_216),
.B1(n_213),
.B2(n_198),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_76),
.B1(n_98),
.B2(n_96),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_213),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_184),
.B(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_83),
.B1(n_106),
.B2(n_78),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_192),
.B1(n_202),
.B2(n_120),
.Y(n_222)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_12),
.B1(n_94),
.B2(n_0),
.Y(n_189)
);

NAND2x1_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_0),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_191),
.B(n_205),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_0),
.B1(n_2),
.B2(n_141),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_126),
.A2(n_0),
.B1(n_2),
.B2(n_141),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_200),
.Y(n_235)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_134),
.A2(n_159),
.B1(n_147),
.B2(n_137),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_142),
.A2(n_128),
.B1(n_157),
.B2(n_132),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_128),
.A2(n_129),
.B1(n_161),
.B2(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_211),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_143),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_130),
.A2(n_122),
.A3(n_145),
.B1(n_124),
.B2(n_125),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_224),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_120),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_219),
.B(n_239),
.Y(n_281)
);

AOI22x1_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_167),
.B1(n_133),
.B2(n_127),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_220),
.A2(n_223),
.B(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_239),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_205),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_192),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_178),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_233),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_181),
.C(n_185),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_191),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_234),
.A2(n_243),
.B(n_244),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_182),
.A2(n_202),
.B1(n_175),
.B2(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_240),
.B1(n_242),
.B2(n_249),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_186),
.B1(n_201),
.B2(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_186),
.B1(n_210),
.B2(n_215),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_173),
.B(n_195),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_185),
.B(n_173),
.C(n_171),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_242),
.C(n_243),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_206),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_257),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_171),
.A2(n_176),
.B1(n_207),
.B2(n_197),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_176),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_177),
.A2(n_214),
.B1(n_198),
.B2(n_196),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_229),
.B1(n_221),
.B2(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_177),
.B(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_225),
.B1(n_227),
.B2(n_220),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_211),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_256),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_188),
.B(n_194),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_260),
.A2(n_285),
.B(n_231),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_264),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_273),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_267),
.B(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_253),
.A2(n_238),
.B1(n_223),
.B2(n_224),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_275),
.B1(n_279),
.B2(n_283),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_222),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_289),
.C(n_271),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_228),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_238),
.B1(n_223),
.B2(n_227),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_225),
.B(n_219),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_246),
.B(n_231),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_278),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_237),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_225),
.A2(n_234),
.B1(n_247),
.B2(n_244),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_244),
.B1(n_245),
.B2(n_240),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_226),
.A2(n_257),
.B1(n_248),
.B2(n_232),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_246),
.B1(n_292),
.B2(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_297),
.A2(n_299),
.B(n_307),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_309),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_294),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_279),
.B(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_289),
.C(n_274),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_314),
.C(n_317),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_288),
.B(n_260),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_320),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_267),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_319),
.B1(n_261),
.B2(n_287),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_269),
.C(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_265),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_275),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_259),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_321),
.C(n_317),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_290),
.B1(n_265),
.B2(n_282),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_261),
.C(n_264),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_322),
.A2(n_298),
.B(n_293),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_278),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_332),
.C(n_335),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_277),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_326),
.B(n_341),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_333),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_302),
.C(n_314),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_294),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_338),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_307),
.C(n_310),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_319),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_304),
.A2(n_320),
.B1(n_298),
.B2(n_296),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_339),
.A2(n_330),
.B1(n_342),
.B2(n_331),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_342),
.Y(n_351)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_343),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_323),
.B1(n_335),
.B2(n_304),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_346),
.A2(n_352),
.B(n_357),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_296),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_358),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_312),
.B(n_301),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_327),
.A2(n_312),
.B(n_301),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_306),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_338),
.A2(n_316),
.B1(n_313),
.B2(n_306),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_329),
.B1(n_322),
.B2(n_337),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_333),
.A2(n_324),
.B1(n_313),
.B2(n_332),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_324),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_374),
.C(n_364),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_325),
.C(n_334),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_366),
.C(n_353),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_361),
.C(n_353),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_352),
.A2(n_357),
.B(n_350),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_346),
.B1(n_351),
.B2(n_360),
.Y(n_378)
);

BUFx12_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_355),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_SL g372 ( 
.A(n_359),
.B(n_348),
.C(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_372),
.Y(n_375)
);

NAND4xp25_ASAP7_75t_SL g373 ( 
.A(n_349),
.B(n_354),
.C(n_347),
.D(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_373),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_351),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_379),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_367),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_381),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_366),
.C(n_365),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_382),
.A2(n_383),
.B(n_370),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_377),
.A2(n_370),
.B(n_373),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_375),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_386),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_388),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_365),
.B(n_371),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_389),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_390),
.C(n_362),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_392),
.A2(n_371),
.B1(n_376),
.B2(n_368),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_378),
.C(n_369),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_394),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_368),
.Y(n_396)
);


endmodule