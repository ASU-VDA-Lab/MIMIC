module fake_aes_3068_n_1257 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1257);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1257;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_659;
wire n_432;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g337 ( .A(n_22), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_189), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_155), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_208), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_68), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_316), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_291), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_1), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_32), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_82), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_179), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_256), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_221), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_232), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_76), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_65), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_41), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_89), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_240), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_115), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_233), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_103), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_125), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_37), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_215), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_44), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_315), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_214), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_55), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_267), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_234), .Y(n_370) );
INVxp33_ASAP7_75t_SL g371 ( .A(n_160), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_272), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_161), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_306), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_5), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_226), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_95), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_260), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_133), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_102), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_180), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_141), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_167), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_11), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_247), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_26), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_190), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_157), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_171), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_16), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_113), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_101), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_24), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_198), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_52), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_70), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_207), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_177), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_33), .Y(n_401) );
INVx4_ASAP7_75t_R g402 ( .A(n_328), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_187), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g404 ( .A(n_333), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_194), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_136), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_276), .Y(n_407) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_308), .Y(n_408) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_210), .B(n_143), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_102), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_209), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_47), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_206), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_223), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_72), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_106), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_312), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_117), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_195), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_87), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_288), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_222), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_134), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_139), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_36), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_81), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_191), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_34), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_193), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_305), .Y(n_430) );
BUFx5_ASAP7_75t_L g431 ( .A(n_21), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_218), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_331), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_97), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_15), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_24), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_20), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_74), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_294), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_81), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_61), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_32), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_280), .Y(n_443) );
INVxp33_ASAP7_75t_SL g444 ( .A(n_148), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_165), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_259), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_262), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_279), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_109), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_302), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_83), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_25), .Y(n_452) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_33), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_336), .Y(n_454) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_51), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_162), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_34), .B(n_170), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_268), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_287), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_152), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_254), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_127), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_19), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_270), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_241), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_146), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_185), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_192), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_211), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_58), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_137), .Y(n_471) );
BUFx8_ASAP7_75t_SL g472 ( .A(n_108), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_1), .Y(n_473) );
INVxp33_ASAP7_75t_SL g474 ( .A(n_55), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_115), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_20), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_238), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_175), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_35), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_27), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_301), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_164), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_153), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_176), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_237), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_126), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_297), .Y(n_487) );
CKINVDCx14_ASAP7_75t_R g488 ( .A(n_120), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_311), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_122), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_61), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_109), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_117), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_85), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_300), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_212), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_35), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_73), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_18), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_213), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_54), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_205), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_41), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_149), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_64), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_36), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_163), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_352), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_488), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_392), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_496), .B(n_0), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_392), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_403), .B(n_2), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_392), .B(n_3), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_403), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_417), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_431), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_450), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_403), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_403), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_426), .B(n_4), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_431), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_431), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_431), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_472), .Y(n_526) );
CKINVDCx8_ASAP7_75t_R g527 ( .A(n_339), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_472), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
INVx6_ASAP7_75t_L g530 ( .A(n_362), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_346), .B(n_4), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_446), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_413), .B(n_5), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_431), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_425), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_431), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_400), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_446), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_431), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_346), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_406), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_365), .B(n_6), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_489), .B(n_6), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_361), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_361), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_365), .Y(n_546) );
NOR2xp67_ASAP7_75t_L g547 ( .A(n_469), .B(n_7), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_446), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_523), .Y(n_549) );
NAND2xp33_ASAP7_75t_R g550 ( .A(n_526), .B(n_474), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_536), .Y(n_551) );
BUFx10_ASAP7_75t_L g552 ( .A(n_508), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_523), .B(n_342), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_531), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_536), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_515), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_536), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
INVx6_ASAP7_75t_L g559 ( .A(n_531), .Y(n_559) );
INVx5_ASAP7_75t_L g560 ( .A(n_530), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_517), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_535), .B(n_342), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_517), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_522), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_530), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_522), .Y(n_566) );
OR2x2_ASAP7_75t_SL g567 ( .A(n_533), .B(n_368), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_527), .B(n_339), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_524), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_525), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_531), .B(n_338), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_525), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_531), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_540), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_521), .B(n_404), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_521), .B(n_452), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_534), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_509), .A2(n_474), .B1(n_414), .B2(n_447), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_515), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_516), .B(n_371), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_530), .Y(n_584) );
INVx4_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_527), .B(n_357), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_518), .B(n_408), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_539), .Y(n_588) );
NOR2x1p5_ASAP7_75t_L g589 ( .A(n_528), .B(n_475), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_510), .B(n_357), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_512), .B(n_408), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_512), .B(n_396), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_577), .B(n_537), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_591), .B(n_543), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_576), .A2(n_533), .B1(n_509), .B2(n_511), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_575), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_576), .B(n_514), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_574), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_559), .A2(n_554), .B1(n_415), .B2(n_440), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_549), .B(n_547), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_574), .B(n_396), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_562), .B(n_540), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_589), .B(n_547), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_553), .B(n_577), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_572), .B(n_540), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_554), .B(n_504), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_554), .B(n_504), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_575), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_552), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_555), .B(n_539), .Y(n_612) );
INVx4_ASAP7_75t_L g613 ( .A(n_559), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_559), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_585), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_568), .B(n_444), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_567), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_590), .B(n_540), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_567), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_592), .B(n_444), .Y(n_620) );
AOI22xp5_ASAP7_75t_SL g621 ( .A1(n_579), .A2(n_541), .B1(n_415), .B2(n_440), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_586), .B(n_544), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_555), .B(n_341), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_557), .B(n_546), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_557), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
O2A1O1Ixp5_ASAP7_75t_L g627 ( .A1(n_566), .A2(n_513), .B(n_546), .C(n_366), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_551), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_552), .B(n_579), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_561), .A2(n_546), .B(n_349), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_589), .B(n_542), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_551), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_561), .A2(n_544), .B1(n_545), .B2(n_542), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_583), .A2(n_451), .B1(n_473), .B2(n_394), .Y(n_634) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_587), .B(n_477), .C(n_464), .Y(n_635) );
BUFx3_ASAP7_75t_L g636 ( .A(n_565), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_563), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_584), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_564), .B(n_343), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_550), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_564), .B(n_404), .Y(n_643) );
NOR3xp33_ASAP7_75t_SL g644 ( .A(n_569), .B(n_503), .C(n_475), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_570), .B(n_344), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_585), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_570), .B(n_545), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_585), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_560), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_571), .B(n_367), .Y(n_651) );
OR2x6_ASAP7_75t_L g652 ( .A(n_571), .B(n_368), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_560), .B(n_464), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_573), .B(n_348), .Y(n_654) );
INVx5_ASAP7_75t_L g655 ( .A(n_560), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_573), .B(n_350), .Y(n_656) );
OR2x6_ASAP7_75t_L g657 ( .A(n_578), .B(n_416), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_578), .A2(n_347), .B1(n_354), .B2(n_337), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_580), .B(n_369), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_556), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_580), .B(n_372), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_566), .B(n_351), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_588), .B(n_381), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_588), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_556), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_560), .B(n_405), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_560), .B(n_407), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_560), .B(n_490), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_556), .B(n_530), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_556), .Y(n_670) );
BUFx6f_ASAP7_75t_SL g671 ( .A(n_582), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_581), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_581), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_581), .B(n_503), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_581), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_581), .B(n_345), .Y(n_677) );
XOR2xp5_ASAP7_75t_L g678 ( .A(n_582), .B(n_477), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_605), .A2(n_428), .B(n_442), .C(n_412), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
AO22x1_ASAP7_75t_L g681 ( .A1(n_611), .A2(n_394), .B1(n_473), .B2(n_451), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_603), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_598), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_614), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_613), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_617), .A2(n_505), .B1(n_463), .B2(n_455), .C(n_453), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_603), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_621), .A2(n_505), .B1(n_481), .B2(n_483), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_626), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_626), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_645), .B(n_478), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_652), .Y(n_692) );
AO21x1_ASAP7_75t_L g693 ( .A1(n_654), .A2(n_360), .B(n_359), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_594), .A2(n_355), .B(n_358), .C(n_356), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_648), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_638), .A2(n_373), .B(n_364), .Y(n_696) );
OR2x6_ASAP7_75t_L g697 ( .A(n_653), .B(n_652), .Y(n_697) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_626), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_619), .A2(n_483), .B1(n_486), .B2(n_481), .Y(n_699) );
NOR2xp33_ASAP7_75t_SL g700 ( .A(n_653), .B(n_486), .Y(n_700) );
O2A1O1Ixp5_ASAP7_75t_L g701 ( .A1(n_627), .A2(n_370), .B(n_376), .C(n_340), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_631), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_640), .A2(n_375), .B(n_374), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_597), .A2(n_379), .B(n_382), .C(n_377), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_652), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_625), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_612), .A2(n_380), .B(n_378), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_657), .A2(n_507), .B1(n_388), .B2(n_393), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_619), .A2(n_507), .B1(n_395), .B2(n_397), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_657), .A2(n_398), .B1(n_410), .B2(n_386), .Y(n_710) );
NOR2xp33_ASAP7_75t_SL g711 ( .A(n_671), .B(n_409), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_657), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_594), .B(n_401), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_596), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_600), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_629), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_604), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_595), .B(n_434), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_604), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_642), .B(n_501), .Y(n_721) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_606), .A2(n_376), .B(n_370), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_602), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_612), .A2(n_384), .B(n_383), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_615), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_624), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_613), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_616), .B(n_418), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_600), .Y(n_729) );
OR2x6_ASAP7_75t_L g730 ( .A(n_607), .B(n_493), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_618), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_636), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_643), .B(n_385), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_608), .B(n_420), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_658), .A2(n_436), .B1(n_437), .B2(n_435), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_658), .A2(n_441), .B1(n_449), .B2(n_438), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_609), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_610), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_649), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_651), .A2(n_661), .B(n_659), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_620), .B(n_387), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_639), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_633), .A2(n_470), .B1(n_479), .B2(n_476), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_601), .B(n_480), .Y(n_744) );
INVx5_ASAP7_75t_L g745 ( .A(n_626), .Y(n_745) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_655), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_663), .A2(n_390), .B(n_389), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g748 ( .A1(n_654), .A2(n_491), .B(n_494), .C(n_492), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_628), .Y(n_749) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_655), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_620), .B(n_497), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_656), .A2(n_498), .B(n_506), .C(n_499), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_671), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_635), .B(n_493), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_656), .B(n_391), .Y(n_755) );
BUFx2_ASAP7_75t_L g756 ( .A(n_644), .Y(n_756) );
INVx3_ASAP7_75t_L g757 ( .A(n_647), .Y(n_757) );
OR2x6_ASAP7_75t_SL g758 ( .A(n_675), .B(n_402), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g759 ( .A1(n_622), .A2(n_457), .B(n_411), .C(n_421), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_664), .B(n_353), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_641), .B(n_419), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_633), .B(n_353), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_646), .B(n_422), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_623), .B(n_423), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_630), .B(n_353), .Y(n_765) );
CKINVDCx8_ASAP7_75t_R g766 ( .A(n_655), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_627), .A2(n_424), .B(n_429), .C(n_427), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_677), .B(n_430), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_632), .B(n_353), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_637), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_623), .B(n_363), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_662), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_655), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_662), .B(n_432), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_650), .B(n_666), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_L g776 ( .A1(n_669), .A2(n_443), .B(n_445), .C(n_433), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_667), .Y(n_777) );
BUFx2_ASAP7_75t_SL g778 ( .A(n_670), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_668), .B(n_448), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_672), .Y(n_780) );
INVx5_ASAP7_75t_L g781 ( .A(n_660), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_660), .B(n_454), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_660), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_L g784 ( .A1(n_673), .A2(n_458), .B(n_459), .C(n_456), .Y(n_784) );
INVx4_ASAP7_75t_L g785 ( .A(n_665), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_665), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_665), .B(n_460), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_676), .B(n_461), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_674), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g790 ( .A1(n_674), .A2(n_465), .B(n_466), .C(n_462), .Y(n_790) );
INVx2_ASAP7_75t_SL g791 ( .A(n_674), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_603), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_597), .B(n_363), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_603), .Y(n_794) );
AOI22x1_ASAP7_75t_L g795 ( .A1(n_638), .A2(n_519), .B1(n_529), .B2(n_520), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_598), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_678), .Y(n_797) );
INVx4_ASAP7_75t_L g798 ( .A(n_611), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_645), .A2(n_468), .B(n_467), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_598), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_594), .A2(n_482), .B(n_484), .C(n_471), .Y(n_801) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_626), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_678), .Y(n_803) );
A2O1A1Ixp33_ASAP7_75t_L g804 ( .A1(n_594), .A2(n_487), .B(n_495), .C(n_485), .Y(n_804) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_722), .A2(n_439), .B(n_399), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_793), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_706), .Y(n_807) );
INVx4_ASAP7_75t_L g808 ( .A(n_697), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_701), .A2(n_502), .B(n_500), .Y(n_809) );
AND2x4_ASAP7_75t_L g810 ( .A(n_682), .B(n_362), .Y(n_810) );
NAND2x1p5_ASAP7_75t_L g811 ( .A(n_692), .B(n_399), .Y(n_811) );
AO21x2_ASAP7_75t_L g812 ( .A1(n_740), .A2(n_439), .B(n_519), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_770), .Y(n_813) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_759), .B(n_520), .C(n_519), .Y(n_814) );
OAI21x1_ASAP7_75t_L g815 ( .A1(n_786), .A2(n_529), .B(n_520), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_789), .A2(n_532), .B(n_529), .Y(n_816) );
OR2x6_ASAP7_75t_L g817 ( .A(n_697), .B(n_532), .Y(n_817) );
AOI31xp67_ASAP7_75t_L g818 ( .A1(n_760), .A2(n_532), .A3(n_548), .B(n_538), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_687), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_792), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_749), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_775), .A2(n_582), .B(n_548), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_794), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_693), .A2(n_538), .A3(n_515), .B(n_9), .Y(n_824) );
OA21x2_ASAP7_75t_L g825 ( .A1(n_779), .A2(n_769), .B(n_762), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_782), .A2(n_787), .B(n_780), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_700), .A2(n_538), .B1(n_515), .B2(n_9), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_779), .A2(n_538), .B(n_123), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_737), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_765), .A2(n_124), .B(n_121), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_795), .A2(n_129), .B(n_128), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_771), .A2(n_131), .B(n_130), .Y(n_832) );
NOR2x1_ASAP7_75t_R g833 ( .A(n_797), .B(n_7), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_731), .Y(n_834) );
AO21x2_ASAP7_75t_L g835 ( .A1(n_767), .A2(n_582), .B(n_132), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_738), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_768), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_713), .B(n_8), .Y(n_838) );
BUFx8_ASAP7_75t_L g839 ( .A(n_773), .Y(n_839) );
AND2x4_ASAP7_75t_L g840 ( .A(n_692), .B(n_10), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_681), .Y(n_841) );
OAI21x1_ASAP7_75t_L g842 ( .A1(n_747), .A2(n_138), .B(n_135), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_783), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_691), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_691), .B(n_12), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_733), .A2(n_142), .B(n_140), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_768), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_708), .Y(n_848) );
NAND2x1p5_ASAP7_75t_L g849 ( .A(n_705), .B(n_13), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_724), .A2(n_145), .B(n_144), .Y(n_850) );
CKINVDCx14_ASAP7_75t_R g851 ( .A(n_708), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_689), .Y(n_852) );
INVx1_ASAP7_75t_SL g853 ( .A(n_803), .Y(n_853) );
AO21x2_ASAP7_75t_L g854 ( .A1(n_790), .A2(n_150), .B(n_147), .Y(n_854) );
OAI21x1_ASAP7_75t_L g855 ( .A1(n_799), .A2(n_154), .B(n_151), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_744), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_751), .B(n_16), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_695), .B(n_17), .Y(n_858) );
NAND2x1p5_ASAP7_75t_L g859 ( .A(n_753), .B(n_17), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_723), .A2(n_158), .B(n_156), .Y(n_860) );
INVxp67_ASAP7_75t_L g861 ( .A(n_700), .Y(n_861) );
OA21x2_ASAP7_75t_L g862 ( .A1(n_755), .A2(n_166), .B(n_159), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_791), .A2(n_169), .B(n_168), .Y(n_863) );
OAI21x1_ASAP7_75t_L g864 ( .A1(n_684), .A2(n_173), .B(n_172), .Y(n_864) );
OAI21x1_ASAP7_75t_L g865 ( .A1(n_715), .A2(n_178), .B(n_174), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_754), .B(n_18), .C(n_19), .Y(n_866) );
OA21x2_ASAP7_75t_L g867 ( .A1(n_755), .A2(n_182), .B(n_181), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_699), .B(n_23), .Y(n_868) );
OAI21x1_ASAP7_75t_L g869 ( .A1(n_707), .A2(n_184), .B(n_183), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_689), .Y(n_870) );
OAI21x1_ASAP7_75t_L g871 ( .A1(n_707), .A2(n_188), .B(n_186), .Y(n_871) );
INVx6_ASAP7_75t_L g872 ( .A(n_798), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_756), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_689), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_690), .Y(n_875) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_753), .B(n_30), .Y(n_876) );
INVxp67_ASAP7_75t_SL g877 ( .A(n_690), .Y(n_877) );
OR2x6_ASAP7_75t_L g878 ( .A(n_798), .B(n_712), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_777), .A2(n_197), .B(n_196), .Y(n_879) );
INVx3_ASAP7_75t_L g880 ( .A(n_766), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_717), .B(n_31), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_690), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_702), .B(n_37), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_746), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_734), .Y(n_885) );
INVx3_ASAP7_75t_L g886 ( .A(n_746), .Y(n_886) );
OA21x2_ASAP7_75t_L g887 ( .A1(n_776), .A2(n_200), .B(n_199), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_719), .B(n_38), .Y(n_888) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_746), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_698), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_726), .B(n_39), .Y(n_891) );
OAI21x1_ASAP7_75t_L g892 ( .A1(n_696), .A2(n_202), .B(n_201), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_732), .B(n_40), .Y(n_893) );
OAI21x1_ASAP7_75t_L g894 ( .A1(n_703), .A2(n_204), .B(n_203), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_698), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_750), .Y(n_896) );
OAI21x1_ASAP7_75t_L g897 ( .A1(n_772), .A2(n_217), .B(n_216), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_741), .A2(n_220), .B(n_219), .Y(n_898) );
CKINVDCx11_ASAP7_75t_R g899 ( .A(n_758), .Y(n_899) );
OAI21x1_ASAP7_75t_L g900 ( .A1(n_685), .A2(n_225), .B(n_224), .Y(n_900) );
OAI21x1_ASAP7_75t_L g901 ( .A1(n_685), .A2(n_228), .B(n_227), .Y(n_901) );
BUFx12f_ASAP7_75t_L g902 ( .A(n_718), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_698), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_743), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_729), .Y(n_905) );
OAI21x1_ASAP7_75t_L g906 ( .A1(n_788), .A2(n_230), .B(n_229), .Y(n_906) );
OAI21x1_ASAP7_75t_L g907 ( .A1(n_725), .A2(n_235), .B(n_231), .Y(n_907) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_739), .A2(n_239), .B(n_236), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_757), .A2(n_243), .B(n_242), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_710), .Y(n_910) );
OAI21x1_ASAP7_75t_L g911 ( .A1(n_757), .A2(n_245), .B(n_244), .Y(n_911) );
OAI21x1_ASAP7_75t_L g912 ( .A1(n_784), .A2(n_248), .B(n_246), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_709), .B(n_714), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_801), .A2(n_250), .B(n_249), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_694), .B(n_43), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_680), .A2(n_252), .B(n_251), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_704), .Y(n_917) );
OA21x2_ASAP7_75t_L g918 ( .A1(n_804), .A2(n_335), .B(n_332), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_743), .A2(n_736), .B1(n_735), .B2(n_728), .Y(n_919) );
AND2x4_ASAP7_75t_SL g920 ( .A(n_732), .B(n_45), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_735), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_716), .B(n_45), .Y(n_922) );
OAI21x1_ASAP7_75t_SL g923 ( .A1(n_785), .A2(n_46), .B(n_48), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_742), .A2(n_330), .B(n_329), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_736), .A2(n_46), .B1(n_48), .B2(n_49), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_802), .Y(n_926) );
INVx2_ASAP7_75t_SL g927 ( .A(n_720), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_683), .A2(n_327), .B(n_326), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_802), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_750), .Y(n_930) );
NOR3xp33_ASAP7_75t_SL g931 ( .A(n_748), .B(n_49), .C(n_50), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_730), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_763), .A2(n_53), .B1(n_54), .B2(n_56), .Y(n_933) );
OAI21x1_ASAP7_75t_L g934 ( .A1(n_742), .A2(n_325), .B(n_324), .Y(n_934) );
OAI21x1_ASAP7_75t_L g935 ( .A1(n_796), .A2(n_800), .B(n_774), .Y(n_935) );
OAI21x1_ASAP7_75t_L g936 ( .A1(n_781), .A2(n_323), .B(n_322), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_752), .A2(n_53), .A3(n_56), .B(n_57), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_763), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_802), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_764), .A2(n_321), .B(n_318), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_679), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_727), .Y(n_942) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_761), .A2(n_281), .B(n_314), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_848), .A2(n_711), .B1(n_745), .B2(n_721), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_851), .A2(n_711), .B1(n_745), .B2(n_778), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_823), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_820), .B(n_59), .Y(n_947) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_919), .A2(n_781), .B1(n_62), .B2(n_63), .C(n_64), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_919), .A2(n_60), .B1(n_62), .B2(n_63), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_891), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_820), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_891), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_837), .A2(n_69), .B1(n_71), .B2(n_72), .C(n_73), .Y(n_953) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_841), .A2(n_71), .B1(n_74), .B2(n_75), .Y(n_954) );
OAI222xp33_ASAP7_75t_L g955 ( .A1(n_861), .A2(n_75), .B1(n_77), .B2(n_78), .C1(n_79), .C2(n_80), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_821), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_841), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_921), .B(n_84), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_891), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_959) );
AO222x2_ASAP7_75t_L g960 ( .A1(n_833), .A2(n_88), .B1(n_89), .B2(n_90), .C1(n_91), .C2(n_92), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_843), .B(n_88), .Y(n_961) );
AOI222xp33_ASAP7_75t_L g962 ( .A1(n_899), .A2(n_90), .B1(n_91), .B2(n_92), .C1(n_93), .C2(n_94), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_843), .B(n_93), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_847), .A2(n_94), .B1(n_95), .B2(n_96), .C(n_97), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_861), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_834), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_819), .B(n_100), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_807), .Y(n_968) );
AOI21xp5_ASAP7_75t_L g969 ( .A1(n_812), .A2(n_273), .B(n_313), .Y(n_969) );
AO21x2_ASAP7_75t_L g970 ( .A1(n_828), .A2(n_274), .B(n_310), .Y(n_970) );
OR2x6_ASAP7_75t_L g971 ( .A(n_817), .B(n_104), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_917), .A2(n_883), .B1(n_941), .B2(n_868), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_813), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_883), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_885), .A2(n_107), .B1(n_108), .B2(n_110), .C(n_111), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_856), .B(n_107), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_838), .B(n_110), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_821), .Y(n_978) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_889), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_812), .A2(n_277), .B(n_309), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_883), .A2(n_112), .B1(n_114), .B2(n_116), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g982 ( .A1(n_822), .A2(n_278), .B(n_307), .Y(n_982) );
AO31x2_ASAP7_75t_L g983 ( .A1(n_844), .A2(n_118), .A3(n_119), .B(n_253), .Y(n_983) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_920), .A2(n_255), .B1(n_257), .B2(n_258), .Y(n_984) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_893), .Y(n_985) );
OAI211xp5_ASAP7_75t_L g986 ( .A1(n_904), .A2(n_261), .B(n_263), .C(n_264), .Y(n_986) );
OAI211xp5_ASAP7_75t_SL g987 ( .A1(n_931), .A2(n_317), .B(n_266), .C(n_269), .Y(n_987) );
INVx2_ASAP7_75t_SL g988 ( .A(n_839), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_805), .A2(n_806), .B(n_825), .Y(n_989) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_857), .A2(n_845), .B(n_888), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_920), .A2(n_265), .B1(n_271), .B2(n_275), .Y(n_991) );
INVx3_ASAP7_75t_L g992 ( .A(n_896), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_805), .A2(n_282), .B(n_283), .Y(n_993) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_827), .A2(n_853), .B1(n_915), .B2(n_922), .C(n_905), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_827), .A2(n_284), .B1(n_285), .B2(n_286), .C(n_289), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_829), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_840), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_893), .Y(n_998) );
AO21x2_ASAP7_75t_L g999 ( .A1(n_828), .A2(n_293), .B(n_295), .Y(n_999) );
AO21x2_ASAP7_75t_L g1000 ( .A1(n_809), .A2(n_296), .B(n_298), .Y(n_1000) );
A2O1A1Ixp33_ASAP7_75t_L g1001 ( .A1(n_866), .A2(n_299), .B(n_303), .C(n_304), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_829), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_817), .A2(n_811), .B1(n_840), .B2(n_881), .Y(n_1003) );
OAI21xp5_ASAP7_75t_L g1004 ( .A1(n_858), .A2(n_814), .B(n_935), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_836), .B(n_808), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_836), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_810), .B(n_904), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_810), .B(n_925), .Y(n_1008) );
AOI21xp5_ASAP7_75t_SL g1009 ( .A1(n_943), .A2(n_811), .B(n_849), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_899), .A2(n_810), .B1(n_932), .B2(n_902), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_902), .A2(n_942), .B1(n_938), .B2(n_933), .Y(n_1011) );
INVx3_ASAP7_75t_L g1012 ( .A(n_930), .Y(n_1012) );
OR2x6_ASAP7_75t_L g1013 ( .A(n_859), .B(n_876), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_933), .A2(n_938), .B1(n_925), .B2(n_927), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_872), .A2(n_878), .B1(n_880), .B2(n_873), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_880), .B(n_878), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_846), .A2(n_825), .B1(n_918), .B2(n_914), .C(n_860), .Y(n_1017) );
AO21x2_ASAP7_75t_L g1018 ( .A1(n_835), .A2(n_831), .B(n_934), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_937), .B(n_930), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_937), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g1021 ( .A1(n_914), .A2(n_918), .B1(n_867), .B2(n_862), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_884), .B(n_886), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_937), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_923), .A2(n_886), .B1(n_884), .B2(n_914), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_937), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_877), .A2(n_889), .B1(n_939), .B2(n_895), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_L g1027 ( .A1(n_912), .A2(n_842), .B(n_855), .C(n_894), .Y(n_1027) );
OAI211xp5_ASAP7_75t_SL g1028 ( .A1(n_898), .A2(n_863), .B(n_939), .C(n_852), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_824), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_862), .A2(n_867), .B(n_815), .Y(n_1030) );
NOR3xp33_ASAP7_75t_L g1031 ( .A(n_842), .B(n_892), .C(n_894), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_889), .B(n_882), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_852), .B(n_895), .Y(n_1033) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_862), .A2(n_815), .B(n_816), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_887), .A2(n_940), .B1(n_934), .B2(n_924), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_870), .B(n_903), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_870), .Y(n_1037) );
AOI33xp33_ASAP7_75t_L g1038 ( .A1(n_874), .A2(n_903), .A3(n_882), .B1(n_929), .B2(n_926), .B3(n_875), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_874), .B(n_929), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g1040 ( .A1(n_816), .A2(n_887), .B(n_926), .Y(n_1040) );
AND2x6_ASAP7_75t_L g1041 ( .A(n_875), .B(n_890), .Y(n_1041) );
A2O1A1Ixp33_ASAP7_75t_L g1042 ( .A1(n_855), .A2(n_892), .B(n_871), .C(n_869), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_900), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_887), .A2(n_940), .B1(n_826), .B2(n_854), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_890), .Y(n_1045) );
OAI21xp5_ASAP7_75t_L g1046 ( .A1(n_830), .A2(n_850), .B(n_906), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_854), .A2(n_830), .B1(n_850), .B2(n_832), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_901), .A2(n_911), .B1(n_909), .B2(n_818), .Y(n_1048) );
AOI21xp5_ASAP7_75t_L g1049 ( .A1(n_907), .A2(n_908), .B(n_865), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_936), .A2(n_879), .B1(n_897), .B2(n_864), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_916), .B(n_928), .Y(n_1051) );
AOI21xp33_ASAP7_75t_L g1052 ( .A1(n_913), .A2(n_861), .B(n_917), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_910), .B(n_919), .Y(n_1053) );
INVx3_ASAP7_75t_L g1054 ( .A(n_896), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_851), .B(n_717), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g1056 ( .A1(n_812), .A2(n_740), .B(n_822), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_820), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_848), .A2(n_851), .B1(n_678), .B2(n_700), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_919), .A2(n_688), .B1(n_599), .B2(n_634), .C(n_579), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_919), .A2(n_686), .B1(n_751), .B2(n_605), .C(n_719), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_910), .B(n_919), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_848), .A2(n_851), .B1(n_678), .B2(n_700), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1006), .Y(n_1063) );
INVx4_ASAP7_75t_L g1064 ( .A(n_971), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_996), .B(n_1002), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_956), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_978), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1053), .B(n_1061), .Y(n_1068) );
AND2x4_ASAP7_75t_SL g1069 ( .A(n_971), .B(n_1013), .Y(n_1069) );
AO21x2_ASAP7_75t_L g1070 ( .A1(n_1021), .A2(n_1030), .B(n_1031), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_985), .B(n_998), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1060), .B(n_1059), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_973), .B(n_968), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_998), .B(n_1057), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1057), .B(n_966), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1007), .B(n_1008), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_946), .B(n_951), .Y(n_1077) );
INVxp67_ASAP7_75t_SL g1078 ( .A(n_997), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1079 ( .A(n_1032), .B(n_979), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_971), .B(n_1020), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1023), .B(n_1025), .Y(n_1081) );
BUFx6f_ASAP7_75t_L g1082 ( .A(n_979), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1058), .B(n_1062), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1005), .B(n_1003), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_972), .B(n_958), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_947), .B(n_1055), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1029), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1038), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1036), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1019), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1033), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1045), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1013), .B(n_1039), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1014), .B(n_949), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1043), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_990), .B(n_1052), .Y(n_1096) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_1041), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_974), .B(n_981), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1037), .B(n_992), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_952), .B(n_983), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_970), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_970), .Y(n_1102) );
AO31x2_ASAP7_75t_L g1103 ( .A1(n_989), .A2(n_1027), .A3(n_1042), .B(n_1056), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_999), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1056), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1012), .B(n_1054), .Y(n_1106) );
NAND4xp25_ASAP7_75t_L g1107 ( .A(n_962), .B(n_1010), .C(n_1011), .D(n_960), .Y(n_1107) );
INVx3_ASAP7_75t_L g1108 ( .A(n_988), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1022), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1004), .Y(n_1110) );
AOI33xp33_ASAP7_75t_L g1111 ( .A1(n_961), .A2(n_963), .A3(n_967), .B1(n_977), .B2(n_954), .B3(n_957), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_950), .B(n_959), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1051), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1051), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1024), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1018), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1046), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_994), .B(n_948), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_984), .B(n_991), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_991), .B(n_1015), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1018), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_1016), .B(n_945), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1026), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_1031), .B(n_980), .Y(n_1124) );
INVx4_ASAP7_75t_R g1125 ( .A(n_1009), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1048), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_976), .B(n_944), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_965), .B(n_975), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_969), .B(n_993), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_953), .B(n_964), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1000), .B(n_1044), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1050), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1040), .Y(n_1133) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_1040), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1047), .B(n_1017), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1035), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1035), .B(n_995), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g1138 ( .A(n_1034), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1049), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_982), .B(n_1001), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1076), .B(n_986), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1076), .B(n_982), .Y(n_1142) );
OAI21xp33_ASAP7_75t_L g1143 ( .A1(n_1107), .A2(n_987), .B(n_955), .Y(n_1143) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_1069), .Y(n_1144) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_1084), .Y(n_1145) );
NAND2xp5_ASAP7_75t_SL g1146 ( .A(n_1064), .B(n_987), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1090), .B(n_1028), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1087), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_1120), .A2(n_1119), .B1(n_1072), .B2(n_1094), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1095), .Y(n_1150) );
INVx3_ASAP7_75t_L g1151 ( .A(n_1097), .Y(n_1151) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1113), .B(n_1114), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1068), .B(n_1081), .Y(n_1153) );
AOI33xp33_ASAP7_75t_L g1154 ( .A1(n_1096), .A2(n_1086), .A3(n_1077), .B1(n_1075), .B2(n_1069), .B3(n_1073), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1095), .Y(n_1155) );
AOI33xp33_ASAP7_75t_L g1156 ( .A1(n_1096), .A2(n_1086), .A3(n_1077), .B1(n_1075), .B2(n_1073), .B3(n_1112), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1083), .B(n_1084), .Y(n_1157) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_1099), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1065), .B(n_1136), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1065), .B(n_1136), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1089), .B(n_1063), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_1113), .B(n_1114), .Y(n_1162) );
OAI31xp33_ASAP7_75t_L g1163 ( .A1(n_1118), .A2(n_1130), .A3(n_1128), .B(n_1098), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1063), .B(n_1066), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1074), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1066), .B(n_1100), .Y(n_1166) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_1108), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1071), .B(n_1085), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1109), .B(n_1111), .Y(n_1169) );
OAI33xp33_ASAP7_75t_L g1170 ( .A1(n_1088), .A2(n_1115), .A3(n_1109), .B1(n_1122), .B2(n_1135), .B3(n_1105), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1091), .B(n_1093), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1100), .B(n_1115), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1091), .B(n_1093), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1067), .B(n_1092), .Y(n_1174) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_1088), .A2(n_1122), .A3(n_1135), .B1(n_1102), .B2(n_1127), .B3(n_1132), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1080), .B(n_1078), .Y(n_1176) );
INVxp67_ASAP7_75t_SL g1177 ( .A(n_1097), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1178 ( .A(n_1099), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1079), .B(n_1117), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1079), .B(n_1117), .Y(n_1180) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_1137), .A2(n_1110), .B1(n_1123), .B2(n_1138), .C(n_1132), .Y(n_1181) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_1167), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1153), .B(n_1106), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1164), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1172), .B(n_1133), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1157), .B(n_1103), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1145), .B(n_1133), .Y(n_1187) );
AOI221xp5_ASAP7_75t_L g1188 ( .A1(n_1163), .A2(n_1124), .B1(n_1139), .B2(n_1134), .C(n_1126), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1159), .B(n_1124), .Y(n_1189) );
NAND4xp25_ASAP7_75t_SL g1190 ( .A(n_1154), .B(n_1125), .C(n_1131), .D(n_1104), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1168), .B(n_1103), .Y(n_1191) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_1178), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1148), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1160), .B(n_1070), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1150), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1150), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1160), .B(n_1129), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1155), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1156), .B(n_1129), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1155), .Y(n_1200) );
AND2x4_ASAP7_75t_SL g1201 ( .A(n_1144), .B(n_1082), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1165), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1174), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1161), .B(n_1121), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1161), .B(n_1121), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1174), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1166), .B(n_1116), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1143), .A2(n_1140), .B1(n_1104), .B2(n_1101), .Y(n_1208) );
NAND4xp75_ASAP7_75t_L g1209 ( .A(n_1188), .B(n_1144), .C(n_1146), .D(n_1169), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1193), .Y(n_1210) );
AOI21xp5_ASAP7_75t_L g1211 ( .A1(n_1190), .A2(n_1175), .B(n_1170), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1195), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1185), .B(n_1147), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1184), .B(n_1149), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1197), .B(n_1179), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1196), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1197), .B(n_1180), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1198), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1185), .B(n_1147), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1200), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1203), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1204), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1186), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1189), .B(n_1162), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1205), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1205), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1194), .B(n_1162), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1191), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1194), .B(n_1152), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1213), .B(n_1202), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1213), .B(n_1183), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1232 ( .A1(n_1211), .A2(n_1199), .B(n_1182), .C(n_1208), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1219), .B(n_1206), .Y(n_1233) );
OAI21xp33_ASAP7_75t_L g1234 ( .A1(n_1222), .A2(n_1187), .B(n_1207), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_1214), .A2(n_1141), .B1(n_1142), .B2(n_1173), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1222), .B(n_1192), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1237 ( .A(n_1232), .B(n_1209), .C(n_1181), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1234), .B(n_1225), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1230), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1238), .B(n_1231), .Y(n_1240) );
OAI211xp5_ASAP7_75t_SL g1241 ( .A1(n_1237), .A2(n_1235), .B(n_1236), .C(n_1233), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g1242 ( .A(n_1239), .Y(n_1242) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_1241), .A2(n_1171), .B1(n_1226), .B2(n_1224), .Y(n_1243) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_1242), .A2(n_1223), .B1(n_1228), .B2(n_1221), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1243), .B(n_1240), .Y(n_1245) );
NOR4xp25_ASAP7_75t_L g1246 ( .A(n_1244), .B(n_1216), .C(n_1212), .D(n_1220), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1245), .Y(n_1247) );
NOR3xp33_ASAP7_75t_SL g1248 ( .A(n_1246), .B(n_1177), .C(n_1210), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1247), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_1248), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1249), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_1250), .A2(n_1229), .B1(n_1227), .B2(n_1158), .Y(n_1252) );
INVx3_ASAP7_75t_L g1253 ( .A(n_1251), .Y(n_1253) );
OAI22xp5_ASAP7_75t_SL g1254 ( .A1(n_1252), .A2(n_1151), .B1(n_1176), .B2(n_1158), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1253), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_1255), .A2(n_1254), .B1(n_1201), .B2(n_1218), .Y(n_1256) );
OAI21xp5_ASAP7_75t_L g1257 ( .A1(n_1256), .A2(n_1215), .B(n_1217), .Y(n_1257) );
endmodule