module real_aes_6604_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g258 ( .A(n_0), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_1), .A2(n_32), .B1(n_102), .B2(n_109), .Y(n_101) );
AOI211xp5_ASAP7_75t_L g151 ( .A1(n_2), .A2(n_152), .B(n_154), .C(n_161), .Y(n_151) );
AOI22xp33_ASAP7_75t_SL g113 ( .A1(n_3), .A2(n_73), .B1(n_114), .B2(n_118), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_4), .A2(n_31), .B1(n_214), .B2(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_5), .B(n_238), .Y(n_247) );
INVx1_ASAP7_75t_L g195 ( .A(n_6), .Y(n_195) );
AND2x6_ASAP7_75t_L g231 ( .A(n_6), .B(n_193), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_6), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_7), .Y(n_100) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_25), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g210 ( .A(n_9), .Y(n_210) );
INVx1_ASAP7_75t_L g251 ( .A(n_10), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_11), .B(n_218), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_12), .B(n_206), .Y(n_322) );
AO32x2_ASAP7_75t_L g264 ( .A1(n_13), .A2(n_205), .A3(n_230), .B1(n_238), .B2(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_14), .B(n_214), .Y(n_290) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_15), .A2(n_29), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_16), .B(n_206), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_17), .A2(n_41), .B1(n_214), .B2(n_267), .Y(n_268) );
AOI22xp33_ASAP7_75t_SL g306 ( .A1(n_18), .A2(n_60), .B1(n_214), .B2(n_218), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_19), .B(n_214), .Y(n_279) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_20), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_21), .B(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_22), .A2(n_81), .B1(n_82), .B2(n_165), .Y(n_80) );
INVx1_ASAP7_75t_L g165 ( .A(n_22), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_23), .B(n_233), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_24), .A2(n_76), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_24), .Y(n_171) );
INVx2_ASAP7_75t_L g216 ( .A(n_26), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_27), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_28), .B(n_233), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g186 ( .A1(n_29), .A2(n_45), .B1(n_55), .B2(n_187), .C(n_188), .Y(n_186) );
INVxp67_ASAP7_75t_L g189 ( .A(n_29), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g142 ( .A1(n_30), .A2(n_72), .B1(n_143), .B2(n_146), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_33), .A2(n_81), .B1(n_82), .B2(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_33), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_34), .B(n_159), .Y(n_158) );
AOI22xp33_ASAP7_75t_SL g122 ( .A1(n_35), .A2(n_62), .B1(n_123), .B2(n_130), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_36), .B(n_214), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_37), .A2(n_68), .B1(n_267), .B2(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g516 ( .A(n_37), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_38), .B(n_214), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_39), .B(n_214), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_40), .B(n_225), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g320 ( .A1(n_42), .A2(n_47), .B1(n_214), .B2(n_218), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_43), .B(n_214), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_44), .A2(n_176), .B1(n_177), .B2(n_182), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_44), .Y(n_182) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_45), .A2(n_64), .B1(n_90), .B2(n_94), .Y(n_97) );
INVxp67_ASAP7_75t_L g190 ( .A(n_45), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_46), .B(n_214), .Y(n_285) );
INVx1_ASAP7_75t_L g193 ( .A(n_48), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_49), .B(n_214), .Y(n_259) );
INVx1_ASAP7_75t_L g209 ( .A(n_50), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_51), .Y(n_187) );
AO32x2_ASAP7_75t_L g302 ( .A1(n_52), .A2(n_230), .A3(n_238), .B1(n_303), .B2(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g179 ( .A(n_53), .Y(n_179) );
INVx1_ASAP7_75t_L g276 ( .A(n_54), .Y(n_276) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_55), .A2(n_71), .B1(n_90), .B2(n_91), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_56), .B(n_218), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_57), .Y(n_155) );
AOI22xp33_ASAP7_75t_SL g134 ( .A1(n_58), .A2(n_70), .B1(n_135), .B2(n_137), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_59), .A2(n_169), .B1(n_172), .B2(n_173), .Y(n_168) );
INVx1_ASAP7_75t_L g172 ( .A(n_59), .Y(n_172) );
AOI22xp5_ASAP7_75t_SL g506 ( .A1(n_60), .A2(n_81), .B1(n_82), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_60), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_61), .A2(n_178), .B1(n_180), .B2(n_181), .Y(n_177) );
INVx1_ASAP7_75t_L g180 ( .A(n_61), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_61), .B(n_267), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_63), .B(n_218), .Y(n_280) );
INVx2_ASAP7_75t_L g207 ( .A(n_65), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_66), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_67), .B(n_218), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_69), .A2(n_77), .B1(n_218), .B2(n_219), .Y(n_319) );
INVx1_ASAP7_75t_L g90 ( .A(n_74), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_74), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_75), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g170 ( .A(n_76), .Y(n_170) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_183), .B1(n_196), .B2(n_500), .C(n_505), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_166), .Y(n_79) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND3x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_133), .C(n_151), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_112), .Y(n_83) );
OAI21xp5_ASAP7_75t_SL g84 ( .A1(n_85), .A2(n_100), .B(n_101), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x6_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x4_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_93), .Y(n_88) );
AND2x2_ASAP7_75t_L g108 ( .A(n_89), .B(n_97), .Y(n_108) );
INVx2_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx2_ASAP7_75t_L g107 ( .A(n_93), .Y(n_107) );
INVx1_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
OR2x2_ASAP7_75t_L g128 ( .A(n_93), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g132 ( .A(n_93), .B(n_129), .Y(n_132) );
AND2x4_ASAP7_75t_L g136 ( .A(n_95), .B(n_132), .Y(n_136) );
AND2x2_ASAP7_75t_L g153 ( .A(n_95), .B(n_141), .Y(n_153) );
AND2x6_ASAP7_75t_L g164 ( .A(n_95), .B(n_127), .Y(n_164) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g126 ( .A(n_96), .B(n_99), .Y(n_126) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g140 ( .A(n_97), .B(n_121), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_97), .B(n_99), .Y(n_150) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g106 ( .A(n_99), .Y(n_106) );
INVx1_ASAP7_75t_L g121 ( .A(n_99), .Y(n_121) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g111 ( .A(n_106), .Y(n_111) );
AND2x2_ASAP7_75t_L g141 ( .A(n_107), .B(n_129), .Y(n_141) );
AND2x4_ASAP7_75t_L g110 ( .A(n_108), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g115 ( .A(n_108), .B(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_122), .Y(n_112) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g160 ( .A(n_117), .B(n_150), .Y(n_160) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x6_ASAP7_75t_L g131 ( .A(n_126), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g145 ( .A(n_126), .B(n_141), .Y(n_145) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_132), .B(n_140), .Y(n_157) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_142), .Y(n_133) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g148 ( .A(n_141), .B(n_149), .Y(n_148) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
OAI21xp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .Y(n_154) );
BUFx2_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx11_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B1(n_174), .B2(n_175), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_169), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g181 ( .A(n_178), .Y(n_181) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_224), .B(n_227), .C(n_228), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
AND3x1_ASAP7_75t_SL g185 ( .A(n_186), .B(n_191), .C(n_194), .Y(n_185) );
INVxp67_ASAP7_75t_L g511 ( .A(n_186), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx1_ASAP7_75t_SL g512 ( .A(n_191), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_191), .A2(n_503), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g522 ( .A(n_191), .Y(n_522) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_192), .B(n_195), .Y(n_515) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_SL g521 ( .A(n_194), .B(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR3x1_ASAP7_75t_L g198 ( .A(n_199), .B(n_428), .C(n_477), .Y(n_198) );
NAND5xp2_ASAP7_75t_L g199 ( .A(n_200), .B(n_343), .C(n_371), .D(n_401), .E(n_415), .Y(n_199) );
AOI221xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_261), .B1(n_293), .B2(n_298), .C(n_309), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_234), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_202), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g323 ( .A(n_203), .Y(n_323) );
AND2x2_ASAP7_75t_L g331 ( .A(n_203), .B(n_237), .Y(n_331) );
AND2x2_ASAP7_75t_L g354 ( .A(n_203), .B(n_236), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_203), .B(n_248), .Y(n_369) );
OR2x2_ASAP7_75t_L g378 ( .A(n_203), .B(n_316), .Y(n_378) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_203), .Y(n_381) );
AND2x2_ASAP7_75t_L g489 ( .A(n_203), .B(n_316), .Y(n_489) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_211), .B(n_232), .Y(n_203) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_204), .A2(n_249), .B(n_260), .Y(n_248) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_206), .Y(n_238) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_207), .B(n_208), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_223), .B(n_230), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_217), .B(n_220), .Y(n_212) );
INVx3_ASAP7_75t_L g275 ( .A(n_214), .Y(n_275) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g267 ( .A(n_215), .Y(n_267) );
BUFx3_ASAP7_75t_L g305 ( .A(n_215), .Y(n_305) );
AND2x6_ASAP7_75t_L g503 ( .A(n_215), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g219 ( .A(n_216), .Y(n_219) );
INVx1_ASAP7_75t_L g226 ( .A(n_216), .Y(n_226) );
INVx2_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_220), .A2(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g246 ( .A(n_220), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_SL g274 ( .A1(n_220), .A2(n_275), .B(n_276), .C(n_277), .Y(n_274) );
INVx5_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OAI22xp5_ASAP7_75t_SL g303 ( .A1(n_221), .A2(n_229), .B1(n_304), .B2(n_306), .Y(n_303) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_222), .Y(n_229) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
INVx1_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
INVx1_ASAP7_75t_L g504 ( .A(n_222), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_224), .A2(n_246), .B(n_258), .C(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_228), .A2(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_229), .A2(n_246), .B1(n_266), .B2(n_268), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_229), .A2(n_246), .B1(n_319), .B2(n_320), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_230), .B(n_317), .C(n_318), .Y(n_342) );
AND2x2_ASAP7_75t_L g502 ( .A(n_230), .B(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_231), .A2(n_240), .B(n_243), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_231), .A2(n_250), .B(n_257), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_231), .A2(n_274), .B(n_278), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_231), .A2(n_284), .B(n_289), .Y(n_283) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_233), .A2(n_273), .B(n_281), .Y(n_272) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_233), .A2(n_283), .B(n_292), .Y(n_282) );
INVx2_ASAP7_75t_L g307 ( .A(n_233), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_234), .B(n_381), .Y(n_437) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OAI311xp33_ASAP7_75t_L g379 ( .A1(n_235), .A2(n_380), .A3(n_381), .B1(n_382), .C1(n_397), .Y(n_379) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
AND2x2_ASAP7_75t_L g340 ( .A(n_236), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g347 ( .A(n_236), .Y(n_347) );
AND2x2_ASAP7_75t_L g468 ( .A(n_236), .B(n_297), .Y(n_468) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_237), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g324 ( .A(n_237), .B(n_248), .Y(n_324) );
AND2x2_ASAP7_75t_L g376 ( .A(n_237), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g390 ( .A(n_237), .B(n_323), .Y(n_390) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_247), .Y(n_237) );
INVx4_ASAP7_75t_L g317 ( .A(n_238), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_246), .Y(n_243) );
INVx2_ASAP7_75t_L g297 ( .A(n_248), .Y(n_297) );
AND2x2_ASAP7_75t_L g339 ( .A(n_248), .B(n_323), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .C(n_254), .Y(n_250) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_255), .A2(n_279), .B(n_280), .Y(n_278) );
INVx4_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_269), .Y(n_261) );
OR2x2_ASAP7_75t_L g434 ( .A(n_262), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_262), .B(n_440), .Y(n_451) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_263), .B(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
AND2x2_ASAP7_75t_L g375 ( .A(n_264), .B(n_302), .Y(n_375) );
AND2x2_ASAP7_75t_L g386 ( .A(n_264), .B(n_282), .Y(n_386) );
AND2x2_ASAP7_75t_L g395 ( .A(n_264), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_269), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_269), .B(n_336), .Y(n_380) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g367 ( .A(n_270), .B(n_326), .Y(n_367) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_282), .Y(n_270) );
INVx2_ASAP7_75t_L g300 ( .A(n_271), .Y(n_300) );
AND2x2_ASAP7_75t_L g394 ( .A(n_271), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g312 ( .A(n_272), .Y(n_312) );
OR2x2_ASAP7_75t_L g411 ( .A(n_272), .B(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_272), .Y(n_474) );
AND2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_308), .Y(n_313) );
INVx1_ASAP7_75t_L g334 ( .A(n_282), .Y(n_334) );
AND2x2_ASAP7_75t_L g355 ( .A(n_282), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g396 ( .A(n_282), .Y(n_396) );
INVx1_ASAP7_75t_L g412 ( .A(n_282), .Y(n_412) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_282), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_295), .B(n_400), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_295), .A2(n_385), .B1(n_434), .B2(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OAI211xp5_ASAP7_75t_SL g477 ( .A1(n_296), .A2(n_478), .B(n_480), .C(n_498), .Y(n_477) );
INVx2_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g388 ( .A(n_297), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g399 ( .A(n_297), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_298), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g372 ( .A(n_299), .B(n_336), .Y(n_372) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g404 ( .A(n_300), .B(n_395), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_300), .B(n_337), .Y(n_423) );
AND2x4_ASAP7_75t_L g359 ( .A(n_301), .B(n_333), .Y(n_359) );
AND2x2_ASAP7_75t_L g497 ( .A(n_301), .B(n_473), .Y(n_497) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
INVx1_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
INVx1_ASAP7_75t_L g436 ( .A(n_302), .Y(n_436) );
OR2x2_ASAP7_75t_L g327 ( .A(n_308), .B(n_312), .Y(n_327) );
AND2x2_ASAP7_75t_L g336 ( .A(n_308), .B(n_337), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_308), .B(n_357), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B1(n_325), .B2(n_328), .C(n_332), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_311), .A2(n_333), .B(n_335), .C(n_338), .Y(n_332) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_312), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_312), .B(n_334), .Y(n_440) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_312), .Y(n_447) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g402 ( .A(n_313), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_324), .Y(n_314) );
INVx2_ASAP7_75t_L g393 ( .A(n_315), .Y(n_393) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_315), .A2(n_326), .B1(n_443), .B2(n_445), .C1(n_446), .C2(n_448), .Y(n_442) );
AND2x2_ASAP7_75t_L g499 ( .A(n_315), .B(n_468), .Y(n_499) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_323), .Y(n_315) );
INVx1_ASAP7_75t_L g389 ( .A(n_316), .Y(n_389) );
AO21x1_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g341 ( .A(n_322), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g427 ( .A(n_324), .B(n_361), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_325), .A2(n_439), .B(n_441), .Y(n_438) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_326), .B(n_333), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_326), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx3_ASAP7_75t_L g392 ( .A(n_330), .Y(n_392) );
OR2x2_ASAP7_75t_L g444 ( .A(n_330), .B(n_366), .Y(n_444) );
AND2x2_ASAP7_75t_L g360 ( .A(n_331), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g398 ( .A(n_331), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_331), .B(n_392), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_331), .B(n_388), .Y(n_414) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_400), .Y(n_418) );
INVxp67_ASAP7_75t_L g350 ( .A(n_333), .Y(n_350) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_335), .A2(n_408), .B1(n_413), .B2(n_414), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_335), .B(n_440), .Y(n_470) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g456 ( .A(n_336), .B(n_447), .Y(n_456) );
AND2x2_ASAP7_75t_L g485 ( .A(n_336), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g490 ( .A(n_336), .B(n_440), .Y(n_490) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
BUFx2_ASAP7_75t_L g409 ( .A(n_337), .Y(n_409) );
INVx1_ASAP7_75t_L g494 ( .A(n_338), .Y(n_494) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_339), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_341), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g362 ( .A(n_341), .Y(n_362) );
INVx3_ASAP7_75t_L g400 ( .A(n_341), .Y(n_400) );
OR2x2_ASAP7_75t_L g466 ( .A(n_341), .B(n_467), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B(n_351), .C(n_363), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_344), .A2(n_481), .B1(n_488), .B2(n_490), .C(n_491), .Y(n_480) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_352), .B(n_358), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_354), .B(n_392), .Y(n_406) );
AND2x2_ASAP7_75t_L g448 ( .A(n_354), .B(n_388), .Y(n_448) );
INVx1_ASAP7_75t_SL g461 ( .A(n_355), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_355), .B(n_409), .Y(n_464) );
INVx1_ASAP7_75t_L g482 ( .A(n_356), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_360), .A2(n_450), .B1(n_452), .B2(n_456), .C(n_457), .Y(n_449) );
AND2x2_ASAP7_75t_L g476 ( .A(n_361), .B(n_468), .Y(n_476) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g460 ( .A(n_362), .Y(n_460) );
AOI21xp33_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_367), .B(n_368), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g431 ( .A(n_366), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g417 ( .A(n_367), .Y(n_417) );
INVx1_ASAP7_75t_L g445 ( .A(n_368), .Y(n_445) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_376), .C(n_379), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_372), .A2(n_410), .A3(n_497), .B(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g472 ( .A(n_375), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g493 ( .A(n_375), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_377), .B(n_392), .Y(n_420) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g495 ( .A(n_378), .B(n_392), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_387), .B1(n_391), .B2(n_394), .Y(n_382) );
NAND2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_386), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g422 ( .A(n_386), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g425 ( .A(n_386), .B(n_409), .Y(n_425) );
AND2x2_ASAP7_75t_L g479 ( .A(n_386), .B(n_474), .Y(n_479) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OAI32xp33_ASAP7_75t_L g457 ( .A1(n_392), .A2(n_426), .A3(n_458), .B1(n_460), .B2(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_405), .C(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_403), .B(n_440), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_404), .A2(n_416), .B1(n_417), .B2(n_418), .C(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g416 ( .A(n_414), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_426), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND4xp25_ASAP7_75t_SL g481 ( .A(n_424), .B(n_482), .C(n_483), .D(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
NAND4xp25_ASAP7_75t_SL g428 ( .A(n_429), .B(n_442), .C(n_449), .D(n_462), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_437), .C(n_438), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g459 ( .A(n_435), .Y(n_459) );
INVx2_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
OR2x2_ASAP7_75t_L g492 ( .A(n_447), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_469), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g488 ( .A(n_468), .B(n_489), .Y(n_488) );
AOI21xp33_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_471), .B(n_475), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_491) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
OAI322xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_508), .A3(n_512), .B1(n_513), .B2(n_516), .C1(n_517), .C2(n_519), .Y(n_505) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
endmodule