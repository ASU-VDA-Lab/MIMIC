module fake_netlist_6_3990_n_1059 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1059);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1059;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_940;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_962;
wire n_824;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_939;
wire n_819;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_77),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_166),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_94),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_141),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_100),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_18),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_44),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_90),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_74),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_57),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_36),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_15),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_24),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_129),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

INVxp33_ASAP7_75t_R g233 ( 
.A(n_53),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_49),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_147),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_84),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_118),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_102),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_131),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_121),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_97),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_157),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_76),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_119),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_155),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_184),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_175),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_15),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_38),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_159),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_89),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_176),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_35),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_202),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_234),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_202),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_0),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_241),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_198),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_244),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_244),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_212),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_214),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_193),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_200),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_224),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_207),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_217),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_225),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_196),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_208),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_209),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_215),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_203),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_275),
.A2(n_195),
.B1(n_218),
.B2(n_238),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_212),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_213),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_201),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_213),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_273),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_307),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_303),
.B(n_201),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_298),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_276),
.A2(n_236),
.B1(n_261),
.B2(n_250),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_277),
.B(n_236),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_250),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_269),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_261),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_272),
.B(n_281),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_262),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_302),
.B(n_196),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_216),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_274),
.B(n_225),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_274),
.A2(n_243),
.B1(n_263),
.B2(n_260),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_305),
.B(n_309),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_266),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_196),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_365),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_342),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_296),
.B1(n_301),
.B2(n_289),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_356),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_369),
.B(n_361),
.Y(n_381)
);

NOR2x1p5_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_276),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_311),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_219),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_340),
.B(n_282),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_221),
.C(n_220),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_325),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_282),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_322),
.B(n_233),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_369),
.B(n_284),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_284),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_286),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_367),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_371),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_338),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_322),
.B(n_225),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_359),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_331),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

NOR2x1p5_ASAP7_75t_L g426 ( 
.A(n_319),
.B(n_286),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_334),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_331),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_353),
.B(n_287),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_319),
.B(n_287),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_367),
.B(n_223),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_328),
.B(n_264),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_328),
.B(n_226),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_328),
.B(n_259),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_389),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_399),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_438),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_354),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_330),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_406),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_406),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_389),
.B(n_370),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_417),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_324),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_379),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_338),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_329),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_329),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_422),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_379),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_324),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_342),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_371),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_413),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_335),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_435),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_392),
.B(n_410),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_395),
.B(n_342),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_438),
.B(n_347),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_395),
.B(n_330),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_R g496 ( 
.A(n_435),
.B(n_322),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_380),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_426),
.B(n_337),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_408),
.B(n_360),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_400),
.Y(n_502)
);

BUFx6f_ASAP7_75t_SL g503 ( 
.A(n_395),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_381),
.B(n_318),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_403),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_386),
.B(n_354),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_419),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_401),
.B(n_345),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_409),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_388),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_445),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_391),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_437),
.B(n_350),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_390),
.B(n_350),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_439),
.B(n_229),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_462),
.A2(n_442),
.B(n_441),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_475),
.B(n_424),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_492),
.A2(n_395),
.B1(n_387),
.B2(n_441),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_475),
.B(n_432),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_446),
.B(n_410),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_462),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_446),
.B(n_375),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_486),
.B(n_395),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_492),
.A2(n_442),
.B1(n_432),
.B2(n_397),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_519),
.B(n_421),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_477),
.B(n_443),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_423),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_486),
.B(n_394),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_448),
.B(n_429),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_477),
.A2(n_396),
.B(n_394),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_465),
.B(n_500),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_502),
.B(n_443),
.Y(n_544)
);

AND2x6_ASAP7_75t_SL g545 ( 
.A(n_471),
.B(n_345),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_504),
.A2(n_378),
.B(n_398),
.C(n_405),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_500),
.B(n_443),
.Y(n_548)
);

BUFx12f_ASAP7_75t_SL g549 ( 
.A(n_471),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_487),
.A2(n_351),
.B1(n_352),
.B2(n_239),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_459),
.B(n_443),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_452),
.B(n_429),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_506),
.B(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_470),
.Y(n_556)
);

AND2x6_ASAP7_75t_SL g557 ( 
.A(n_471),
.B(n_351),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_509),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_352),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_467),
.B(n_430),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_455),
.B(n_430),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_476),
.A2(n_407),
.B(n_414),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_488),
.B(n_407),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_494),
.B(n_431),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_378),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_494),
.B(n_348),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_457),
.B(n_378),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_458),
.B(n_398),
.Y(n_570)
);

AOI221xp5_ASAP7_75t_L g571 ( 
.A1(n_460),
.A2(n_230),
.B1(n_232),
.B2(n_258),
.C(n_242),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_450),
.B(n_358),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_512),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_464),
.A2(n_245),
.B1(n_252),
.B2(n_254),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_478),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_256),
.C(n_255),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_515),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_524),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_495),
.A2(n_416),
.B1(n_415),
.B2(n_414),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_565),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_529),
.B(n_461),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_549),
.B(n_496),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_530),
.B(n_540),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_529),
.B(n_460),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_531),
.A2(n_463),
.B1(n_466),
.B2(n_480),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_531),
.A2(n_495),
.B(n_482),
.C(n_485),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_533),
.A2(n_490),
.B(n_483),
.C(n_489),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_SL g593 ( 
.A(n_577),
.B(n_496),
.C(n_493),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_560),
.B(n_507),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_552),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_550),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_559),
.B(n_537),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_552),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_575),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_547),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_R g604 ( 
.A(n_577),
.B(n_503),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_557),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_536),
.B(n_453),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_559),
.B(n_537),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_551),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_558),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_576),
.A2(n_497),
.B1(n_491),
.B2(n_505),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_559),
.B(n_514),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_574),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_521),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_580),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_541),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_527),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_544),
.B(n_503),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_566),
.B(n_522),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_451),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_555),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_555),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_528),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_578),
.B(n_514),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_579),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_567),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_571),
.B(n_499),
.Y(n_629)
);

AO22x1_ASAP7_75t_L g630 ( 
.A1(n_561),
.A2(n_501),
.B1(n_499),
.B2(n_516),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_570),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_R g633 ( 
.A(n_538),
.B(n_447),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_499),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_588),
.A2(n_553),
.B1(n_539),
.B2(n_568),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_591),
.A2(n_562),
.B(n_542),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_584),
.B(n_571),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_627),
.A2(n_542),
.B(n_562),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_627),
.A2(n_525),
.B(n_581),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_583),
.Y(n_640)
);

AO31x2_ASAP7_75t_L g641 ( 
.A1(n_591),
.A2(n_525),
.A3(n_546),
.B(n_520),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_621),
.A2(n_548),
.B(n_535),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_606),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_623),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_619),
.B(n_518),
.Y(n_645)
);

AO31x2_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_415),
.A3(n_416),
.B(n_510),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_629),
.A2(n_589),
.B(n_593),
.C(n_620),
.Y(n_647)
);

AO31x2_ASAP7_75t_L g648 ( 
.A1(n_592),
.A2(n_498),
.A3(n_484),
.B(n_454),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_618),
.A2(n_449),
.B1(n_398),
.B2(n_391),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_583),
.Y(n_651)
);

AOI211x1_ASAP7_75t_L g652 ( 
.A1(n_594),
.A2(n_597),
.B(n_602),
.C(n_595),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_632),
.A2(n_385),
.B(n_341),
.Y(n_653)
);

OAI21xp33_ASAP7_75t_L g654 ( 
.A1(n_589),
.A2(n_362),
.B(n_358),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_601),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_610),
.A2(n_427),
.B(n_37),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_620),
.B(n_240),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_616),
.A2(n_427),
.A3(n_363),
.B(n_362),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_610),
.A2(n_427),
.B(n_40),
.Y(n_659)
);

OAI21x1_ASAP7_75t_SL g660 ( 
.A1(n_590),
.A2(n_41),
.B(n_34),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_596),
.A2(n_624),
.B(n_615),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_628),
.B(n_358),
.Y(n_662)
);

OAI21x1_ASAP7_75t_SL g663 ( 
.A1(n_590),
.A2(n_614),
.B(n_609),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_614),
.A2(n_427),
.B(n_43),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_630),
.A2(n_362),
.B(n_358),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_599),
.A2(n_45),
.B(n_42),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_617),
.A2(n_47),
.B(n_46),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_615),
.A2(n_363),
.B(n_362),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_626),
.A2(n_51),
.B(n_50),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_613),
.A2(n_582),
.A3(n_593),
.B(n_631),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_625),
.A2(n_611),
.B1(n_624),
.B2(n_607),
.Y(n_671)
);

AOI21x1_ASAP7_75t_L g672 ( 
.A1(n_625),
.A2(n_363),
.B(n_54),
.Y(n_672)
);

INVx6_ASAP7_75t_L g673 ( 
.A(n_582),
.Y(n_673)
);

OAI21x1_ASAP7_75t_SL g674 ( 
.A1(n_604),
.A2(n_56),
.B(n_52),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_59),
.B(n_58),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_601),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_611),
.A2(n_363),
.B1(n_240),
.B2(n_3),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_612),
.A2(n_240),
.B1(n_2),
.B2(n_3),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_598),
.A2(n_62),
.B(n_61),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_613),
.B(n_1),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_631),
.A2(n_623),
.B(n_622),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_63),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g683 ( 
.A(n_622),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_636),
.A2(n_631),
.B(n_623),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_640),
.B(n_603),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_647),
.A2(n_608),
.B1(n_634),
.B2(n_607),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_638),
.A2(n_631),
.B(n_633),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_661),
.A2(n_634),
.B(n_600),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_649),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_651),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_637),
.B(n_585),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_673),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_643),
.B(n_657),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_642),
.A2(n_604),
.B(n_605),
.Y(n_694)
);

O2A1O1Ixp5_ASAP7_75t_L g695 ( 
.A1(n_665),
.A2(n_633),
.B(n_619),
.C(n_585),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_635),
.A2(n_654),
.B(n_645),
.Y(n_696)
);

AOI221x1_ASAP7_75t_L g697 ( 
.A1(n_680),
.A2(n_623),
.B1(n_601),
.B2(n_587),
.C(n_7),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_655),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_652),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_673),
.Y(n_700)
);

AO32x2_ASAP7_75t_L g701 ( 
.A1(n_671),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_SL g702 ( 
.A1(n_677),
.A2(n_601),
.B(n_6),
.C(n_8),
.Y(n_702)
);

AOI221xp5_ASAP7_75t_L g703 ( 
.A1(n_678),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_644),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_662),
.B(n_64),
.Y(n_705)
);

INVx6_ASAP7_75t_L g706 ( 
.A(n_655),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_682),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_670),
.B(n_10),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_663),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_682),
.B(n_65),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_676),
.B(n_66),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_670),
.B(n_11),
.Y(n_712)
);

CKINVDCx6p67_ASAP7_75t_R g713 ( 
.A(n_644),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_683),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_714)
);

AO31x2_ASAP7_75t_L g715 ( 
.A1(n_668),
.A2(n_108),
.A3(n_189),
.B(n_188),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_681),
.A2(n_639),
.B(n_656),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_650),
.Y(n_717)
);

CKINVDCx8_ASAP7_75t_R g718 ( 
.A(n_644),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_670),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_672),
.B(n_67),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_641),
.B(n_12),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_674),
.B(n_13),
.C(n_14),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_659),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_653),
.A2(n_109),
.B(n_187),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_664),
.A2(n_107),
.B(n_186),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_675),
.A2(n_191),
.B(n_106),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_679),
.B(n_16),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_648),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_641),
.B(n_17),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_646),
.A2(n_110),
.A3(n_183),
.B(n_182),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_666),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_660),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_667),
.A2(n_185),
.B(n_111),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_641),
.B(n_22),
.Y(n_734)
);

AO31x2_ASAP7_75t_L g735 ( 
.A1(n_646),
.A2(n_648),
.A3(n_658),
.B(n_669),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_646),
.Y(n_736)
);

AOI221x1_ASAP7_75t_L g737 ( 
.A1(n_658),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_737)
);

OA21x2_ASAP7_75t_L g738 ( 
.A1(n_658),
.A2(n_114),
.B(n_181),
.Y(n_738)
);

AO31x2_ASAP7_75t_L g739 ( 
.A1(n_635),
.A2(n_112),
.A3(n_180),
.B(n_178),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_637),
.B(n_23),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_647),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_643),
.B(n_26),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_636),
.A2(n_177),
.B(n_105),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_638),
.A2(n_104),
.B(n_173),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_638),
.A2(n_103),
.B(n_172),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_688),
.B(n_69),
.Y(n_746)
);

INVx6_ASAP7_75t_L g747 ( 
.A(n_704),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_691),
.A2(n_703),
.B1(n_740),
.B2(n_694),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_690),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_722),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_686),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_717),
.A2(n_710),
.B1(n_693),
.B2(n_743),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_710),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_753)
);

CKINVDCx11_ASAP7_75t_R g754 ( 
.A(n_700),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_741),
.A2(n_32),
.B1(n_33),
.B2(n_70),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_707),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_689),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_713),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_718),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_759)
);

CKINVDCx11_ASAP7_75t_R g760 ( 
.A(n_698),
.Y(n_760)
);

INVxp33_ASAP7_75t_SL g761 ( 
.A(n_685),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_697),
.A2(n_75),
.B1(n_81),
.B2(n_82),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_706),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_692),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_684),
.Y(n_765)
);

BUFx8_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_706),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_714),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_742),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_709),
.A2(n_712),
.B1(n_727),
.B2(n_729),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_721),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_734),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_708),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_696),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_699),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_720),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_720),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_736),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

CKINVDCx8_ASAP7_75t_R g781 ( 
.A(n_738),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_719),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_695),
.Y(n_783)
);

NOR2x1_ASAP7_75t_L g784 ( 
.A(n_705),
.B(n_101),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_701),
.Y(n_785)
);

INVx6_ASAP7_75t_L g786 ( 
.A(n_687),
.Y(n_786)
);

CKINVDCx11_ASAP7_75t_R g787 ( 
.A(n_702),
.Y(n_787)
);

CKINVDCx14_ASAP7_75t_R g788 ( 
.A(n_701),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_726),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_733),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_701),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_716),
.Y(n_792)
);

BUFx4f_ASAP7_75t_SL g793 ( 
.A(n_730),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_730),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_739),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_735),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_735),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_739),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_737),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_779),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_774),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_797),
.A2(n_796),
.B(n_745),
.Y(n_802)
);

AO21x2_ASAP7_75t_L g803 ( 
.A1(n_794),
.A2(n_723),
.B(n_731),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_786),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_780),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_772),
.B(n_715),
.Y(n_806)
);

NOR2x1_ASAP7_75t_SL g807 ( 
.A(n_773),
.B(n_738),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_757),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_786),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_786),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_782),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_765),
.B(n_715),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_785),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_776),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_781),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_795),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_788),
.B(n_771),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_792),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_798),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_793),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_746),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_799),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_778),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_783),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_753),
.A2(n_732),
.B1(n_725),
.B2(n_744),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_755),
.A2(n_724),
.B(n_135),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_746),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_783),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_747),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_747),
.Y(n_831)
);

OAI21x1_ASAP7_75t_L g832 ( 
.A1(n_789),
.A2(n_133),
.B(n_136),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_752),
.B(n_138),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_769),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_790),
.A2(n_139),
.B(n_142),
.Y(n_836)
);

AO21x1_ASAP7_75t_L g837 ( 
.A1(n_762),
.A2(n_143),
.B(n_144),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_748),
.B(n_145),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_755),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_769),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_787),
.A2(n_146),
.B1(n_150),
.B2(n_153),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_784),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_764),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_775),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_764),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_807),
.A2(n_759),
.B(n_750),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_804),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_805),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_809),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_809),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_805),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_811),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_845),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_809),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_813),
.B(n_749),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_810),
.B(n_767),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_813),
.B(n_753),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_805),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_810),
.B(n_768),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_810),
.B(n_768),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_SL g862 ( 
.A1(n_823),
.A2(n_817),
.B1(n_839),
.B2(n_834),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_808),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_814),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_804),
.B(n_749),
.Y(n_866)
);

AO21x2_ASAP7_75t_L g867 ( 
.A1(n_807),
.A2(n_759),
.B(n_751),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_802),
.A2(n_777),
.B(n_767),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_822),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_821),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_845),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_811),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_804),
.Y(n_873)
);

OA21x2_ASAP7_75t_L g874 ( 
.A1(n_802),
.A2(n_827),
.B(n_816),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_864),
.B(n_822),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_856),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_861),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_861),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_864),
.B(n_817),
.Y(n_879)
);

AND2x4_ASAP7_75t_SL g880 ( 
.A(n_866),
.B(n_821),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_854),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_858),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_858),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_849),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_852),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_866),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_854),
.B(n_815),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_858),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_863),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_854),
.B(n_815),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_848),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_852),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_850),
.B(n_815),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_846),
.A2(n_837),
.B(n_827),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_848),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_851),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_866),
.B(n_818),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_851),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_850),
.B(n_804),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_862),
.B(n_825),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_881),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_877),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_881),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_894),
.A2(n_837),
.B1(n_846),
.B2(n_867),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_878),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_889),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_882),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_880),
.B(n_876),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_879),
.B(n_855),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_885),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_882),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_900),
.A2(n_872),
.B(n_869),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_892),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_875),
.B(n_855),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_880),
.B(n_876),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_888),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_887),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_902),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_910),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_907),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_SL g921 ( 
.A(n_904),
.B(n_862),
.C(n_818),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_907),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_905),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_914),
.B(n_855),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_906),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_910),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_886),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_908),
.B(n_886),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_909),
.B(n_754),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_926),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_929),
.A2(n_904),
.B1(n_823),
.B2(n_839),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_918),
.Y(n_932)
);

INVx3_ASAP7_75t_R g933 ( 
.A(n_920),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_927),
.B(n_928),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_928),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_919),
.B(n_915),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_929),
.B(n_915),
.Y(n_937)
);

AO221x2_ASAP7_75t_L g938 ( 
.A1(n_931),
.A2(n_921),
.B1(n_925),
.B2(n_923),
.C(n_903),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_931),
.A2(n_846),
.B1(n_857),
.B2(n_867),
.Y(n_939)
);

AO221x2_ASAP7_75t_L g940 ( 
.A1(n_930),
.A2(n_903),
.B1(n_901),
.B2(n_920),
.C(n_922),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_937),
.B(n_756),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_936),
.B(n_924),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_936),
.B(n_912),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_942),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_935),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_941),
.B(n_934),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_938),
.B(n_935),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_943),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_939),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_940),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_940),
.B(n_932),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_940),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_941),
.B(n_917),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_952),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_952),
.Y(n_955)
);

AOI211xp5_ASAP7_75t_L g956 ( 
.A1(n_949),
.A2(n_933),
.B(n_838),
.C(n_834),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_949),
.A2(n_846),
.B1(n_867),
.B2(n_844),
.Y(n_957)
);

OAI221xp5_ASAP7_75t_L g958 ( 
.A1(n_947),
.A2(n_838),
.B1(n_922),
.B2(n_800),
.C(n_901),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

AND2x2_ASAP7_75t_SL g960 ( 
.A(n_946),
.B(n_761),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_953),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_954),
.B(n_955),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_961),
.B(n_951),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_959),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_948),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_956),
.A2(n_950),
.B(n_945),
.Y(n_967)
);

OAI21xp33_ASAP7_75t_SL g968 ( 
.A1(n_957),
.A2(n_913),
.B(n_897),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_962),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_956),
.B1(n_913),
.B2(n_800),
.Y(n_970)
);

OAI221xp5_ASAP7_75t_L g971 ( 
.A1(n_967),
.A2(n_800),
.B1(n_841),
.B2(n_818),
.C(n_829),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_966),
.A2(n_912),
.B(n_770),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_968),
.A2(n_758),
.B(n_842),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_964),
.A2(n_820),
.B1(n_829),
.B2(n_825),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_969),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_970),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_971),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_972),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_973),
.B(n_965),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_969),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_969),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_977),
.Y(n_983)
);

AND3x4_ASAP7_75t_L g984 ( 
.A(n_979),
.B(n_760),
.C(n_856),
.Y(n_984)
);

NAND4xp25_ASAP7_75t_L g985 ( 
.A(n_980),
.B(n_820),
.C(n_842),
.D(n_857),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_975),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_981),
.B(n_766),
.Y(n_987)
);

NAND3xp33_ASAP7_75t_SL g988 ( 
.A(n_982),
.B(n_853),
.C(n_871),
.Y(n_988)
);

NOR3x1_ASAP7_75t_L g989 ( 
.A(n_978),
.B(n_763),
.C(n_833),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_976),
.B(n_766),
.Y(n_990)
);

AOI211xp5_ASAP7_75t_L g991 ( 
.A1(n_990),
.A2(n_976),
.B(n_826),
.C(n_833),
.Y(n_991)
);

NAND5xp2_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_860),
.C(n_859),
.D(n_857),
.E(n_844),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_987),
.B(n_843),
.C(n_836),
.Y(n_993)
);

OAI211xp5_ASAP7_75t_L g994 ( 
.A1(n_986),
.A2(n_871),
.B(n_853),
.C(n_843),
.Y(n_994)
);

NAND4xp25_ASAP7_75t_L g995 ( 
.A(n_989),
.B(n_860),
.C(n_859),
.D(n_821),
.Y(n_995)
);

OAI211xp5_ASAP7_75t_SL g996 ( 
.A1(n_984),
.A2(n_985),
.B(n_988),
.C(n_826),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_983),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_988),
.B(n_158),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_990),
.A2(n_916),
.B(n_911),
.C(n_832),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_997),
.A2(n_916),
.B(n_911),
.C(n_843),
.Y(n_1000)
);

OAI222xp33_ASAP7_75t_L g1001 ( 
.A1(n_996),
.A2(n_869),
.B1(n_843),
.B2(n_887),
.C1(n_890),
.C2(n_870),
.Y(n_1001)
);

OAI211xp5_ASAP7_75t_SL g1002 ( 
.A1(n_991),
.A2(n_830),
.B(n_831),
.C(n_835),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_998),
.B(n_993),
.C(n_994),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_995),
.B(n_884),
.C(n_835),
.Y(n_1004)
);

AOI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_992),
.A2(n_884),
.B(n_835),
.C(n_840),
.Y(n_1005)
);

NAND4xp25_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_860),
.C(n_859),
.D(n_821),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_997),
.A2(n_846),
.B(n_867),
.C(n_840),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_856),
.Y(n_1008)
);

AOI221x1_ASAP7_75t_L g1009 ( 
.A1(n_1002),
.A2(n_884),
.B1(n_856),
.B2(n_896),
.C(n_895),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_1004),
.Y(n_1010)
);

AOI221x1_ASAP7_75t_L g1011 ( 
.A1(n_1006),
.A2(n_884),
.B1(n_856),
.B2(n_896),
.C(n_895),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1000),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1005),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_SL g1014 ( 
.A1(n_1001),
.A2(n_831),
.B1(n_830),
.B2(n_840),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_1007),
.B(n_831),
.C(n_830),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_L g1016 ( 
.A(n_1003),
.B(n_884),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_SL g1017 ( 
.A(n_1003),
.B(n_890),
.C(n_824),
.Y(n_1017)
);

OR4x2_ASAP7_75t_L g1018 ( 
.A(n_1017),
.B(n_867),
.C(n_870),
.D(n_847),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1008),
.Y(n_1019)
);

AND3x2_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_824),
.C(n_828),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1013),
.B(n_893),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1016),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_1010),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_1011),
.B(n_870),
.C(n_893),
.Y(n_1025)
);

OR3x1_ASAP7_75t_L g1026 ( 
.A(n_1014),
.B(n_819),
.C(n_816),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_1009),
.B(n_898),
.C(n_891),
.Y(n_1027)
);

XNOR2xp5_ASAP7_75t_L g1028 ( 
.A(n_1008),
.B(n_160),
.Y(n_1028)
);

OR3x2_ASAP7_75t_L g1029 ( 
.A(n_1013),
.B(n_161),
.C(n_162),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_1010),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_899),
.B1(n_849),
.B2(n_870),
.Y(n_1031)
);

OAI211xp5_ASAP7_75t_SL g1032 ( 
.A1(n_1019),
.A2(n_164),
.B(n_165),
.C(n_167),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1029),
.A2(n_849),
.B1(n_898),
.B2(n_891),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_1028),
.Y(n_1034)
);

OA22x2_ASAP7_75t_L g1035 ( 
.A1(n_1020),
.A2(n_899),
.B1(n_883),
.B2(n_888),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_1030),
.B(n_168),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1024),
.A2(n_836),
.B(n_832),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1021),
.A2(n_849),
.B1(n_870),
.B2(n_847),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_1022),
.B(n_832),
.C(n_836),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1034),
.Y(n_1040)
);

INVxp33_ASAP7_75t_SL g1041 ( 
.A(n_1036),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1032),
.A2(n_1025),
.B1(n_1026),
.B2(n_1027),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1035),
.Y(n_1043)
);

AO22x2_ASAP7_75t_L g1044 ( 
.A1(n_1033),
.A2(n_1018),
.B1(n_883),
.B2(n_850),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1031),
.A2(n_849),
.B1(n_847),
.B2(n_873),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1038),
.A2(n_849),
.B1(n_847),
.B2(n_873),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1037),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1040),
.A2(n_1039),
.B1(n_849),
.B2(n_873),
.Y(n_1048)
);

NOR2xp67_ASAP7_75t_L g1049 ( 
.A(n_1042),
.B(n_171),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1043),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1044),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_1050),
.A2(n_1047),
.B1(n_1041),
.B2(n_1046),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1052),
.B(n_1051),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1053),
.A2(n_1049),
.B(n_1048),
.Y(n_1054)
);

OAI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1054),
.A2(n_1045),
.B1(n_849),
.B2(n_819),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1055),
.A2(n_174),
.B(n_812),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_1056),
.B(n_868),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_850),
.B1(n_874),
.B2(n_803),
.Y(n_1058)
);

AOI211xp5_ASAP7_75t_L g1059 ( 
.A1(n_1058),
.A2(n_806),
.B(n_812),
.C(n_865),
.Y(n_1059)
);


endmodule