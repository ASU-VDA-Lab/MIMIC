module fake_jpeg_15946_n_59 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_10),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_22),
.C(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_47),
.B1(n_12),
.B2(n_15),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_14),
.C(n_17),
.Y(n_43)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_8),
.B(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_52),
.B(n_51),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_53),
.B(n_54),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_41),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_43),
.C(n_44),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_45),
.Y(n_59)
);


endmodule