module fake_jpeg_9221_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_43),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_49),
.B1(n_59),
.B2(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_20),
.B1(n_30),
.B2(n_19),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_21),
.B1(n_24),
.B2(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_36),
.B1(n_39),
.B2(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_72),
.B1(n_47),
.B2(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_36),
.B1(n_43),
.B2(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_75),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_18),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_41),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_41),
.A3(n_42),
.B1(n_28),
.B2(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_87),
.B1(n_57),
.B2(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_28),
.B1(n_42),
.B2(n_41),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_46),
.C(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_101),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_58),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_62),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_106),
.B(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_72),
.B1(n_87),
.B2(n_54),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_65),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_73),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_32),
.B(n_44),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_83),
.B1(n_69),
.B2(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_117),
.B1(n_131),
.B2(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_69),
.B1(n_85),
.B2(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_122),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_122),
.A3(n_128),
.B1(n_116),
.B2(n_123),
.C1(n_124),
.C2(n_101),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_134),
.Y(n_136)
);

OAI22x1_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_82),
.B1(n_80),
.B2(n_23),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_68),
.B1(n_53),
.B2(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_44),
.B1(n_48),
.B2(n_73),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_82),
.C(n_2),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_63),
.B1(n_53),
.B2(n_68),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_76),
.B1(n_112),
.B2(n_78),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_143),
.B1(n_114),
.B2(n_117),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_92),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_140),
.C(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_125),
.C(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_145),
.B1(n_152),
.B2(n_153),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_96),
.B1(n_97),
.B2(n_89),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_76),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_101),
.C(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_89),
.B1(n_68),
.B2(n_53),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_104),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_105),
.B(n_106),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_131),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_90),
.B(n_102),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_150),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_161),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_159),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_103),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_178),
.C(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_102),
.B1(n_132),
.B2(n_78),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_153),
.B1(n_78),
.B2(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_104),
.C(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_99),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_158),
.B(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_176),
.B1(n_168),
.B2(n_16),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.C(n_191),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_143),
.B1(n_138),
.B2(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_189),
.B1(n_194),
.B2(n_195),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_138),
.B1(n_151),
.B2(n_136),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.C(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_179),
.B1(n_164),
.B2(n_160),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_42),
.C(n_27),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_167),
.C(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_179),
.B1(n_166),
.B2(n_160),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_206),
.B1(n_207),
.B2(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_177),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_203),
.B(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_212),
.C(n_3),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_1),
.Y(n_209)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_15),
.B(n_5),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_195),
.B(n_197),
.C(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_27),
.C(n_23),
.Y(n_212)
);

AO21x1_ASAP7_75t_SL g213 ( 
.A1(n_193),
.A2(n_187),
.B(n_28),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_196),
.B(n_2),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_211),
.C(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_4),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_3),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_4),
.B(n_6),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_224),
.C(n_217),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_210),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_4),
.C(n_6),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_202),
.B1(n_215),
.B2(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_7),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_233),
.C(n_216),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_233),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_204),
.B(n_8),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_227),
.B1(n_235),
.B2(n_214),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_234),
.C(n_205),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_7),
.B(n_8),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_9),
.C(n_10),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_249),
.C(n_13),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_251),
.B(n_10),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);


endmodule