module fake_jpeg_13370_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_25),
.Y(n_37)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_22),
.B1(n_14),
.B2(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_13),
.B1(n_10),
.B2(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_18),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_11),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_23),
.C(n_11),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_47),
.B1(n_39),
.B2(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_15),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_36),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_40),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_30),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_54),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_57),
.B(n_52),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_58),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_62),
.B(n_51),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_36),
.B(n_41),
.C(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_36),
.Y(n_67)
);


endmodule