module fake_jpeg_10915_n_236 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_37),
.B(n_54),
.Y(n_101)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_83),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_34),
.B1(n_15),
.B2(n_21),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_69),
.B(n_81),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_15),
.B(n_33),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_56),
.B1(n_52),
.B2(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_47),
.C(n_14),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_73),
.C(n_66),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_40),
.A2(n_34),
.B1(n_21),
.B2(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_33),
.B(n_31),
.C(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_102),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_103),
.B1(n_90),
.B2(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_39),
.B(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_38),
.B(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_25),
.B1(n_24),
.B2(n_6),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_73),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_95),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_121),
.Y(n_138)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_109),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_44),
.B1(n_5),
.B2(n_6),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_112),
.B1(n_116),
.B2(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_8),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_11),
.B1(n_12),
.B2(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_11),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_86),
.B1(n_76),
.B2(n_87),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_70),
.B1(n_109),
.B2(n_110),
.Y(n_155)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_73),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_66),
.B(n_82),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_80),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_70),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_92),
.C(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_153),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_155),
.B(n_142),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_131),
.C(n_118),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_134),
.B(n_120),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_78),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_127),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_121),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_162),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_126),
.B1(n_116),
.B2(n_122),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_176),
.B1(n_143),
.B2(n_142),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_158),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_173),
.C(n_178),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_131),
.B1(n_124),
.B2(n_114),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_132),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_114),
.B1(n_124),
.B2(n_155),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_146),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_157),
.B(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_194),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_140),
.B(n_144),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_174),
.B(n_175),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_186),
.B(n_188),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_192),
.B(n_191),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_146),
.C(n_138),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_141),
.C(n_139),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_172),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_199),
.B1(n_205),
.B2(n_195),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_181),
.C(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_212),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_208),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_180),
.C(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_181),
.C(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_190),
.C(n_178),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_197),
.B1(n_184),
.B2(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_215),
.B1(n_197),
.B2(n_210),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_213),
.B(n_200),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_189),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_224),
.B(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_211),
.B1(n_182),
.B2(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_228),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_182),
.A3(n_217),
.B1(n_186),
.B2(n_220),
.C1(n_176),
.C2(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_151),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_227),
.A2(n_177),
.B(n_148),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_157),
.B(n_148),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_230),
.B1(n_151),
.B2(n_152),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_233),
.B(n_152),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_139),
.Y(n_236)
);


endmodule