module fake_jpeg_15553_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g110 ( 
.A(n_39),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_25),
.A2(n_12),
.B1(n_6),
.B2(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_16),
.B1(n_21),
.B2(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_61),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_6),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_62),
.Y(n_120)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_66),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_36),
.B1(n_26),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_21),
.B1(n_18),
.B2(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_21),
.B1(n_37),
.B2(n_33),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_78),
.A2(n_87),
.B1(n_95),
.B2(n_104),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_20),
.B1(n_32),
.B2(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_84),
.B(n_92),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_15),
.B1(n_35),
.B2(n_22),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_20),
.B1(n_35),
.B2(n_15),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_33),
.B1(n_19),
.B2(n_22),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_98),
.B(n_100),
.C(n_103),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_42),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_44),
.A2(n_34),
.B1(n_29),
.B2(n_31),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_28),
.B1(n_38),
.B2(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_4),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_48),
.A2(n_52),
.B1(n_64),
.B2(n_60),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_8),
.B1(n_10),
.B2(n_2),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_28),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_39),
.B(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_17),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_39),
.B(n_28),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_28),
.B1(n_38),
.B2(n_17),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_17),
.Y(n_145)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_121),
.B(n_123),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_131),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_38),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_28),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_142),
.Y(n_175)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_130),
.B(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_110),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_38),
.B(n_17),
.C(n_3),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_5),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_90),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_136),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_80),
.B(n_38),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_146),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_8),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_163),
.B1(n_172),
.B2(n_74),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_75),
.B(n_109),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_109),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_70),
.B(n_8),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_154),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_4),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_170),
.B1(n_74),
.B2(n_117),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_4),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_164),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_82),
.B(n_5),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_83),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_11),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_171),
.Y(n_187)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_11),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_97),
.B1(n_89),
.B2(n_86),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_177),
.A2(n_178),
.B1(n_192),
.B2(n_169),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_97),
.B1(n_72),
.B2(n_86),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_182),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_5),
.B(n_9),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_196),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_125),
.A2(n_162),
.B(n_134),
.C(n_143),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_72),
.B1(n_106),
.B2(n_119),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_124),
.C(n_136),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_206),
.C(n_212),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_125),
.A2(n_76),
.B1(n_96),
.B2(n_114),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_204),
.B1(n_210),
.B2(n_158),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_96),
.B1(n_114),
.B2(n_88),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_149),
.A2(n_10),
.B1(n_11),
.B2(n_0),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_169),
.B1(n_165),
.B2(n_148),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_10),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_170),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_186),
.B1(n_214),
.B2(n_195),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_130),
.B(n_1),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_148),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_149),
.A2(n_139),
.B(n_126),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_196),
.C(n_210),
.Y(n_251)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_232),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_221),
.A2(n_227),
.B1(n_239),
.B2(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_222),
.B(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_137),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_229),
.B(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_137),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_261),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_193),
.B(n_128),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_238),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_165),
.B1(n_135),
.B2(n_153),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_144),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_155),
.B1(n_129),
.B2(n_132),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_179),
.B(n_211),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_229),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_158),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_185),
.B1(n_199),
.B2(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_188),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_256),
.B(n_258),
.C(n_221),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_175),
.A2(n_193),
.B1(n_181),
.B2(n_219),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_178),
.A2(n_183),
.B1(n_201),
.B2(n_192),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_207),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_175),
.A2(n_181),
.B1(n_218),
.B2(n_178),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_184),
.A2(n_175),
.B1(n_216),
.B2(n_181),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_195),
.A2(n_214),
.B1(n_211),
.B2(n_207),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_208),
.B1(n_198),
.B2(n_194),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_258),
.B1(n_235),
.B2(n_245),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_191),
.B1(n_186),
.B2(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_218),
.B(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_191),
.B(n_180),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_269),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_265),
.A2(n_268),
.B(n_280),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_179),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_266),
.B(n_274),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_230),
.C(n_249),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g320 ( 
.A1(n_278),
.A2(n_294),
.B1(n_292),
.B2(n_280),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_247),
.A3(n_253),
.B1(n_250),
.B2(n_223),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_251),
.B1(n_227),
.B2(n_225),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_270),
.B1(n_279),
.B2(n_274),
.Y(n_321)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_223),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_288),
.B(n_289),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_234),
.C(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_293),
.C(n_266),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_232),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_290),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_224),
.A2(n_226),
.B(n_234),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_232),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_260),
.B(n_231),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_268),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_261),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_278),
.B(n_292),
.C(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_224),
.B1(n_236),
.B2(n_241),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_300),
.B1(n_294),
.B2(n_272),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_299),
.B(n_307),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_238),
.B1(n_228),
.B2(n_237),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_237),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_220),
.Y(n_304)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_305),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_220),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_308),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_310),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_265),
.B(n_289),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_311),
.A2(n_320),
.B1(n_306),
.B2(n_296),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_307),
.Y(n_330)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_314),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_264),
.B(n_271),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_315),
.B(n_305),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_317),
.C(n_318),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_273),
.C(n_291),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_293),
.C(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_279),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_319),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_294),
.B1(n_267),
.B2(n_262),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_283),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_322),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

AOI22x1_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_294),
.B1(n_268),
.B2(n_267),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_308),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_338),
.B1(n_310),
.B2(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_315),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_333),
.B(n_337),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_299),
.B1(n_300),
.B2(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_306),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_297),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_344),
.C(n_321),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_323),
.C(n_318),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_348),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_351),
.B1(n_326),
.B2(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_353),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_352),
.B(n_356),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_302),
.C(n_314),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_313),
.B1(n_301),
.B2(n_298),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_342),
.B1(n_324),
.B2(n_331),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_301),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_361),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_298),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_328),
.B(n_332),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_351),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_366),
.A2(n_354),
.B1(n_334),
.B2(n_349),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_368),
.B(n_371),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_346),
.A2(n_341),
.B1(n_327),
.B2(n_331),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_372),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_341),
.B(n_342),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_334),
.C(n_324),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_354),
.B1(n_352),
.B2(n_358),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_348),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_376),
.B(n_379),
.Y(n_384)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_356),
.C(n_350),
.Y(n_379)
);

NAND4xp25_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_373),
.C(n_369),
.D(n_366),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_375),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_385),
.A2(n_387),
.B(n_383),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_367),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_386),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_365),
.Y(n_387)
);

OAI321xp33_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_364),
.A3(n_378),
.B1(n_385),
.B2(n_377),
.C(n_382),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_389),
.B(n_380),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_391),
.A2(n_379),
.B(n_363),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_392),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_393),
.A2(n_345),
.B1(n_370),
.B2(n_376),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_363),
.C(n_361),
.Y(n_395)
);


endmodule