module fake_jpeg_24684_n_73 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_37),
.B(n_0),
.Y(n_46)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_1),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_48),
.B1(n_11),
.B2(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_36),
.B1(n_34),
.B2(n_5),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_63),
.B1(n_59),
.B2(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_24),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

AO221x1_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_30),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_31),
.Y(n_73)
);


endmodule