module fake_jpeg_1899_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_0),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_68),
.B1(n_71),
.B2(n_69),
.Y(n_82)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_56),
.B1(n_57),
.B2(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_52),
.B1(n_58),
.B2(n_44),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_58),
.C(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_43),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_62),
.A3(n_43),
.B1(n_61),
.B2(n_50),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_84),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_52),
.B1(n_60),
.B2(n_46),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_1),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_45),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_25),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_70),
.C(n_19),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_86),
.C(n_78),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_2),
.CI(n_5),
.CON(n_102),
.SN(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_13),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_123)
);

OR2x4_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_11),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_14),
.B(n_15),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_26),
.B1(n_41),
.B2(n_40),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_106),
.B(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_22),
.C(n_39),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_127),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_120),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_123),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_15),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_16),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_98),
.C(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_139),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_102),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_102),
.B(n_21),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_154),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_20),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_143),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_142),
.B(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.C(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_130),
.C(n_134),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_130),
.C(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_145),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_156),
.C(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_141),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_166),
.B(n_148),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_164),
.B(n_141),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_145),
.B(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_136),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_37),
.C(n_38),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_42),
.Y(n_175)
);


endmodule