module fake_jpeg_9672_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_28),
.B1(n_17),
.B2(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_25),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_36),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_66),
.C(n_84),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_35),
.C(n_21),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_0),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_13),
.C(n_12),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_70),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_74),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_31),
.B(n_22),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_86),
.B(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_38),
.B1(n_41),
.B2(n_33),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_79),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_33),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_17),
.B1(n_16),
.B2(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_94),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_67),
.B(n_64),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_105),
.B(n_60),
.Y(n_119)
);

XNOR2x2_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_61),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_97),
.B1(n_72),
.B2(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_110),
.B1(n_112),
.B2(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_69),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_3),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_118),
.B1(n_128),
.B2(n_134),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_123),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_121),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_61),
.B(n_71),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_107),
.B(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_5),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_88),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_81),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_87),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_111),
.A3(n_103),
.B1(n_105),
.B2(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_88),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_133),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_151),
.B(n_152),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_101),
.B1(n_110),
.B2(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_117),
.C(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_165),
.C(n_142),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_118),
.B(n_120),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_163),
.B(n_136),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_138),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OA21x2_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_137),
.B(n_144),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_93),
.A3(n_146),
.B1(n_137),
.B2(n_142),
.C1(n_123),
.C2(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_124),
.C(n_129),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_128),
.B1(n_147),
.B2(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_177),
.B1(n_164),
.B2(n_162),
.Y(n_183)
);

AOI31xp67_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_155),
.A3(n_165),
.B(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_175),
.C(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_95),
.C(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_145),
.B1(n_125),
.B2(n_95),
.Y(n_177)
);

AOI21x1_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_166),
.B(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_183),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_166),
.B(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_186),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_182),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_153),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_153),
.B(n_8),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_169),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_176),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.C(n_192),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_196),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_185),
.B(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_5),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_195),
.C(n_9),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_8),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_199),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_200),
.B(n_9),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_201),
.Y(n_204)
);


endmodule