module fake_jpeg_27064_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_52),
.B1(n_59),
.B2(n_34),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_51),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_19),
.B1(n_32),
.B2(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_1),
.B(n_2),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_45),
.B(n_2),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_75),
.B1(n_40),
.B2(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_38),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_68),
.C(n_41),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_79),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_34),
.C(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_80),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_36),
.B1(n_37),
.B2(n_34),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_60),
.A3(n_58),
.B1(n_44),
.B2(n_52),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_28),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_81),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_31),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_41),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_40),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_36),
.B1(n_59),
.B2(n_47),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_47),
.B1(n_46),
.B2(n_48),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_106),
.B1(n_110),
.B2(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_97),
.B1(n_109),
.B2(n_82),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_104),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_36),
.B1(n_48),
.B2(n_46),
.Y(n_97)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_46),
.B1(n_17),
.B2(n_26),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_116),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_41),
.B1(n_27),
.B2(n_22),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_61),
.Y(n_118)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_41),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_68),
.C(n_70),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_127),
.C(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_134),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_67),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_112),
.C(n_117),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_65),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_71),
.C(n_102),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_62),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_88),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_100),
.B1(n_94),
.B2(n_80),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_87),
.C(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_16),
.B1(n_29),
.B2(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_143),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_88),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_31),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_98),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_85),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_115),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_176),
.B(n_131),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_162),
.C(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_86),
.B1(n_81),
.B2(n_64),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_171),
.B1(n_174),
.B2(n_126),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_100),
.B1(n_86),
.B2(n_74),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_124),
.B1(n_138),
.B2(n_56),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_168),
.B1(n_134),
.B2(n_124),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_98),
.B1(n_72),
.B2(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_126),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_96),
.B(n_107),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_177),
.B(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_99),
.C(n_76),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_173),
.C(n_178),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_31),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_31),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_172),
.C(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_94),
.B1(n_73),
.B2(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_179),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_137),
.C(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_99),
.C(n_114),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_17),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_175),
.B(n_23),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_27),
.B(n_22),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_1),
.B(n_3),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_114),
.C(n_54),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_147),
.B1(n_152),
.B2(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_193),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_195),
.B1(n_201),
.B2(n_208),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_199),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_141),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_135),
.B(n_140),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_162),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_30),
.B(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_174),
.B(n_28),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_3),
.C(n_5),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_25),
.C(n_21),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_168),
.C(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_210),
.B1(n_3),
.B2(n_4),
.Y(n_234)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_218),
.B1(n_229),
.B2(n_210),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_225),
.C(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_172),
.B1(n_148),
.B2(n_160),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_160),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_164),
.C(n_25),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_185),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_15),
.C(n_14),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_13),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_13),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_235),
.C(n_199),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_204),
.B(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_180),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_237),
.B(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_242),
.B(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_209),
.B1(n_208),
.B2(n_193),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_240),
.B1(n_244),
.B2(n_251),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_186),
.B1(n_182),
.B2(n_187),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_210),
.B1(n_194),
.B2(n_202),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_195),
.B(n_200),
.C(n_181),
.Y(n_245)
);

OAI22x1_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_188),
.B1(n_206),
.B2(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_254),
.B(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_203),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_190),
.B1(n_201),
.B2(n_192),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_211),
.B1(n_184),
.B2(n_189),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_184),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_225),
.C(n_231),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_262),
.C(n_264),
.Y(n_273)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_249),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_183),
.C(n_198),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_259),
.B(n_270),
.Y(n_282)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_215),
.B(n_243),
.C(n_218),
.D(n_220),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_243),
.C(n_252),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_205),
.C(n_207),
.Y(n_262)
);

BUFx12f_ASAP7_75t_SL g263 ( 
.A(n_245),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_240),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_222),
.C(n_233),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_235),
.C(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_6),
.C(n_7),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_196),
.B1(n_203),
.B2(n_6),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_258),
.B1(n_261),
.B2(n_266),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_260),
.B(n_9),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_242),
.B1(n_239),
.B2(n_251),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_285),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_203),
.B1(n_252),
.B2(n_13),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_283),
.B1(n_286),
.B2(n_285),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_3),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_5),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_284),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_267),
.B1(n_270),
.B2(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_8),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_8),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_257),
.C(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_9),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_9),
.B(n_10),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_281),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_273),
.C(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_284),
.B1(n_275),
.B2(n_11),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_9),
.B(n_10),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_10),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.C(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_10),
.C(n_11),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_292),
.C(n_299),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_300),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_300),
.B(n_308),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

AOI221xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_310),
.B1(n_316),
.B2(n_313),
.C(n_317),
.Y(n_319)
);

AOI211xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_309),
.B(n_303),
.C(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_11),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_11),
.C(n_12),
.Y(n_322)
);


endmodule