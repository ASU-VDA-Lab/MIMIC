module real_jpeg_4082_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_0),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_0),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_0),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_1),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_1),
.A2(n_150),
.B1(n_198),
.B2(n_267),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_1),
.A2(n_72),
.B1(n_267),
.B2(n_388),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g444 ( 
.A1(n_1),
.A2(n_267),
.B1(n_324),
.B2(n_445),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_2),
.Y(n_333)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_2),
.Y(n_348)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_2),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_2),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_91),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_3),
.A2(n_91),
.B1(n_119),
.B2(n_178),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_3),
.A2(n_91),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_4),
.Y(n_327)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_6),
.A2(n_56),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_6),
.A2(n_56),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_6),
.A2(n_56),
.B1(n_271),
.B2(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_7),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_7),
.B(n_116),
.C(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_7),
.B(n_77),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_159),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_7),
.B(n_96),
.Y(n_255)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_99),
.B1(n_105),
.B2(n_127),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_10),
.A2(n_99),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_10),
.A2(n_99),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_11),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_11),
.A2(n_199),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_11),
.A2(n_96),
.B1(n_199),
.B2(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_11),
.A2(n_52),
.B1(n_199),
.B2(n_352),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_105),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_13),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_13),
.A2(n_158),
.B1(n_188),
.B2(n_192),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_13),
.A2(n_158),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_13),
.A2(n_158),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_15),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_15),
.A2(n_177),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_15),
.A2(n_177),
.B1(n_293),
.B2(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_15),
.A2(n_55),
.B1(n_177),
.B2(n_396),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_16),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_16),
.A2(n_64),
.B1(n_165),
.B2(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_16),
.A2(n_64),
.B1(n_127),
.B2(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_16),
.A2(n_64),
.B1(n_272),
.B2(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_521),
.B(n_524),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_139),
.B(n_520),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_135),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_27),
.B(n_135),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_128),
.C(n_132),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_28),
.A2(n_29),
.B1(n_516),
.B2(n_517),
.Y(n_515)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_65),
.C(n_100),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_30),
.B(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_31),
.A2(n_57),
.B1(n_59),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_31),
.A2(n_57),
.B1(n_129),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_31),
.A2(n_350),
.B(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_31),
.A2(n_41),
.B1(n_395),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_31),
.A2(n_51),
.B1(n_57),
.B2(n_493),
.Y(n_492)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_32),
.A2(n_346),
.B(n_349),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_32),
.B(n_351),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_32),
.A2(n_58),
.B(n_523),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_41),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_39),
.Y(n_354)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_41),
.B(n_154),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_50),
.Y(n_41)
);

OAI32xp33_ASAP7_75t_L g317 ( 
.A1(n_42),
.A2(n_318),
.A3(n_321),
.B1(n_325),
.B2(n_330),
.Y(n_317)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_45),
.Y(n_273)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_46),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_46),
.Y(n_261)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_49),
.Y(n_388)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_57),
.A2(n_419),
.B(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_58),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_58),
.B(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_65),
.A2(n_100),
.B1(n_101),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_65),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_66),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_66),
.A2(n_92),
.B1(n_292),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_66),
.A2(n_92),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_66),
.A2(n_85),
.B1(n_92),
.B2(n_497),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_67)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_68),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_71),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_76),
.Y(n_329)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_76),
.Y(n_393)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_76),
.Y(n_432)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_77),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_77),
.A2(n_133),
.B1(n_297),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_77),
.A2(n_133),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_80),
.Y(n_384)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_81),
.Y(n_380)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_92),
.B(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_92),
.A2(n_292),
.B(n_296),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_97),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_100),
.A2(n_101),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_100),
.B(n_492),
.C(n_495),
.Y(n_503)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_115),
.B(n_126),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_149),
.B(n_155),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_102),
.A2(n_196),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_102),
.A2(n_155),
.B(n_246),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_102),
.A2(n_245),
.B1(n_362),
.B2(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_103),
.B(n_156),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_103),
.A2(n_159),
.B1(n_376),
.B2(n_381),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_103),
.A2(n_159),
.B1(n_381),
.B2(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_103),
.A2(n_159),
.B1(n_401),
.B2(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx5_ASAP7_75t_SL g249 ( 
.A(n_112),
.Y(n_249)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_115),
.A2(n_196),
.B(n_202),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_115),
.A2(n_202),
.B(n_362),
.Y(n_361)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_126),
.Y(n_435)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_127),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_128),
.B(n_132),
.Y(n_517)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_133),
.A2(n_252),
.B(n_256),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_133),
.B(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_133),
.A2(n_256),
.B(n_460),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_135),
.B(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_135),
.B(n_522),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_136),
.Y(n_523)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_514),
.B(n_519),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_486),
.B(n_511),
.Y(n_140)
);

OAI311xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_365),
.A3(n_462),
.B1(n_480),
.C1(n_485),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_311),
.B(n_364),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_283),
.B(n_310),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_239),
.B(n_282),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_205),
.B(n_238),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_170),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_147),
.B(n_170),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_160),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_148),
.A2(n_160),
.B1(n_161),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_148),
.Y(n_236)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_152),
.B(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_152),
.Y(n_403)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g402 ( 
.A(n_153),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_180),
.B(n_185),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_154),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_154),
.B(n_331),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_154),
.A2(n_330),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_193),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_171),
.B(n_194),
.C(n_204),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_180),
.B(n_185),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_180),
.A2(n_211),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_180),
.A2(n_234),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_180),
.A2(n_372),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_181),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_181),
.A2(n_265),
.B1(n_301),
.B2(n_307),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_181),
.A2(n_338),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_190),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_203),
.B2(n_204),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_229),
.B(n_237),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_215),
.B(n_228),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_227),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_227),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_226),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_218),
.Y(n_374)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_264),
.B(n_269),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_235),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_241),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_262),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_250),
.C(n_262),
.Y(n_284)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_271),
.A3(n_274),
.B1(n_276),
.B2(n_280),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_275),
.Y(n_377)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_284),
.B(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_309),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_289),
.C(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_299),
.C(n_300),
.Y(n_340)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_307),
.Y(n_405)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_312),
.B(n_313),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_343),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_314)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_334),
.B2(n_335),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_317),
.B(n_334),
.Y(n_458)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_340),
.B(n_341),
.C(n_343),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_355),
.B2(n_363),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_344),
.B(n_356),
.C(n_361),
.Y(n_471)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_355),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_SL g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_448),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_366),
.A2(n_448),
.B(n_481),
.C(n_484),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_422),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_367),
.B(n_422),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_398),
.C(n_407),
.Y(n_367)
);

FAx1_ASAP7_75t_SL g461 ( 
.A(n_368),
.B(n_398),
.CI(n_407),
.CON(n_461),
.SN(n_461)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_385),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_386),
.C(n_394),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_370),
.B(n_375),
.Y(n_454)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_376),
.Y(n_410)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_389),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_404),
.B2(n_406),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_404),
.A2(n_406),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_404),
.A2(n_439),
.B(n_442),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_417),
.C(n_420),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_409),
.B(n_411),
.Y(n_470)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_420),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_426),
.C(n_437),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_437),
.B2(n_438),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_433),
.B(n_436),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_434),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_436),
.B(n_489),
.CI(n_490),
.CON(n_488),
.SN(n_488)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_436),
.B(n_489),
.C(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_447),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_454),
.C(n_455),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_450),
.A2(n_451),
.B1(n_454),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_473),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_461),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_475),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_482),
.B(n_483),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_472),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.C(n_471),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_478),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_470),
.B1(n_471),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_477),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_500),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_499),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_499),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_488),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_492),
.B1(n_494),
.B2(n_498),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_492),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_502),
.C(n_506),
.Y(n_518)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_494),
.Y(n_498)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_510),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_510),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_518),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_518),
.Y(n_519)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);


endmodule