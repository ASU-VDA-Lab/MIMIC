module real_aes_313_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_848, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_848;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g580 ( .A(n_0), .B(n_154), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g830 ( .A1(n_2), .A2(n_11), .B1(n_831), .B2(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_2), .Y(n_832) );
INVx1_ASAP7_75t_L g161 ( .A(n_3), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_4), .B(n_514), .Y(n_540) );
NAND2xp33_ASAP7_75t_SL g599 ( .A(n_5), .B(n_160), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_6), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g592 ( .A(n_7), .Y(n_592) );
INVx1_ASAP7_75t_L g210 ( .A(n_8), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_10), .Y(n_201) );
AOI222xp33_ASAP7_75t_SL g104 ( .A1(n_11), .A2(n_105), .B1(n_120), .B2(n_818), .C1(n_820), .C2(n_838), .Y(n_104) );
AND2x2_ASAP7_75t_L g538 ( .A(n_11), .B(n_188), .Y(n_538) );
INVxp67_ASAP7_75t_L g831 ( .A(n_11), .Y(n_831) );
INVx2_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
AOI221x1_ASAP7_75t_L g595 ( .A1(n_15), .A2(n_167), .B1(n_516), .B2(n_596), .C(n_598), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_16), .B(n_514), .Y(n_561) );
INVx1_ASAP7_75t_L g815 ( .A(n_17), .Y(n_815) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
INVx1_ASAP7_75t_L g152 ( .A(n_19), .Y(n_152) );
INVx1_ASAP7_75t_SL g271 ( .A(n_20), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_21), .B(n_146), .Y(n_244) );
AOI33xp33_ASAP7_75t_L g220 ( .A1(n_22), .A2(n_53), .A3(n_140), .B1(n_181), .B2(n_221), .B3(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_23), .A2(n_516), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_24), .B(n_154), .Y(n_543) );
AOI221xp5_ASAP7_75t_SL g570 ( .A1(n_25), .A2(n_42), .B1(n_514), .B2(n_516), .C(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g195 ( .A(n_26), .Y(n_195) );
OAI22x1_ASAP7_75t_R g806 ( .A1(n_27), .A2(n_51), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_27), .Y(n_808) );
OR2x2_ASAP7_75t_L g134 ( .A(n_28), .B(n_92), .Y(n_134) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_28), .A2(n_92), .B(n_135), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_29), .B(n_157), .Y(n_565) );
INVxp67_ASAP7_75t_L g594 ( .A(n_30), .Y(n_594) );
AND2x2_ASAP7_75t_L g535 ( .A(n_31), .B(n_187), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_32), .B(n_172), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_33), .A2(n_516), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_34), .B(n_157), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_35), .A2(n_52), .B1(n_357), .B2(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_35), .Y(n_827) );
AND2x2_ASAP7_75t_L g160 ( .A(n_36), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g176 ( .A(n_36), .B(n_143), .Y(n_176) );
INVx1_ASAP7_75t_L g180 ( .A(n_36), .Y(n_180) );
OR2x6_ASAP7_75t_L g116 ( .A(n_37), .B(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_38), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_39), .B(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_40), .A2(n_133), .B1(n_168), .B2(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_41), .B(n_246), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_43), .A2(n_84), .B1(n_178), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_44), .B(n_146), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_45), .B(n_154), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_46), .B(n_207), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_47), .B(n_146), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_48), .Y(n_241) );
AND2x2_ASAP7_75t_L g583 ( .A(n_49), .B(n_187), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_50), .B(n_187), .Y(n_574) );
INVx1_ASAP7_75t_L g807 ( .A(n_51), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_52), .Y(n_357) );
HB1xp67_ASAP7_75t_SL g428 ( .A(n_52), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_54), .B(n_146), .Y(n_185) );
OAI22x1_ASAP7_75t_R g825 ( .A1(n_55), .A2(n_826), .B1(n_828), .B2(n_829), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_55), .Y(n_829) );
INVx1_ASAP7_75t_L g141 ( .A(n_56), .Y(n_141) );
INVx1_ASAP7_75t_L g148 ( .A(n_56), .Y(n_148) );
AND2x2_ASAP7_75t_L g186 ( .A(n_57), .B(n_187), .Y(n_186) );
AOI221xp5_ASAP7_75t_L g208 ( .A1(n_58), .A2(n_77), .B1(n_172), .B2(n_178), .C(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_59), .B(n_172), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_60), .B(n_514), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_61), .B(n_168), .Y(n_203) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_62), .B(n_803), .Y(n_802) );
AOI21xp5_ASAP7_75t_SL g230 ( .A1(n_63), .A2(n_178), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g526 ( .A(n_64), .B(n_187), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_65), .B(n_157), .Y(n_581) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_67), .B(n_154), .Y(n_524) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_68), .B(n_188), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_69), .A2(n_516), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g184 ( .A(n_70), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_71), .B(n_157), .Y(n_544) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_72), .B(n_207), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_73), .A2(n_178), .B(n_183), .Y(n_177) );
INVx1_ASAP7_75t_L g143 ( .A(n_74), .Y(n_143) );
INVx1_ASAP7_75t_L g150 ( .A(n_74), .Y(n_150) );
AOI22x1_ASAP7_75t_L g803 ( .A1(n_75), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_75), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_76), .B(n_172), .Y(n_223) );
AND2x2_ASAP7_75t_L g273 ( .A(n_78), .B(n_167), .Y(n_273) );
INVx1_ASAP7_75t_L g144 ( .A(n_79), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_80), .A2(n_178), .B(n_270), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_81), .A2(n_178), .B(n_215), .C(n_243), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_82), .A2(n_87), .B1(n_172), .B2(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_83), .B(n_514), .Y(n_525) );
INVx1_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
AND2x2_ASAP7_75t_SL g228 ( .A(n_86), .B(n_167), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_88), .A2(n_178), .B1(n_218), .B2(n_219), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_89), .B(n_154), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_90), .B(n_154), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_91), .A2(n_516), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g232 ( .A(n_93), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_94), .B(n_157), .Y(n_523) );
AND2x2_ASAP7_75t_L g224 ( .A(n_95), .B(n_167), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_96), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_97), .B(n_514), .Y(n_582) );
INVxp67_ASAP7_75t_L g597 ( .A(n_98), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_99), .B(n_157), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_100), .A2(n_516), .B(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g111 ( .A(n_101), .Y(n_111) );
BUFx2_ASAP7_75t_SL g844 ( .A(n_101), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_102), .B(n_146), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_103), .B(n_837), .Y(n_836) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_SL g819 ( .A(n_109), .B(n_111), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_109), .A2(n_842), .B(n_845), .Y(n_841) );
INVx2_ASAP7_75t_L g835 ( .A(n_112), .Y(n_835) );
INVx1_ASAP7_75t_SL g837 ( .A(n_112), .Y(n_837) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g846 ( .A(n_113), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x6_ASAP7_75t_SL g504 ( .A(n_114), .B(n_116), .Y(n_504) );
OR2x6_ASAP7_75t_SL g800 ( .A(n_114), .B(n_115), .Y(n_800) );
OR2x2_ASAP7_75t_L g817 ( .A(n_114), .B(n_116), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_809), .Y(n_121) );
NAND2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_801), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_501), .B1(n_505), .B2(n_798), .Y(n_123) );
INVx1_ASAP7_75t_L g812 ( .A(n_124), .Y(n_812) );
AOI211x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_357), .B(n_358), .C(n_498), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND4x1_ASAP7_75t_L g498 ( .A(n_126), .B(n_359), .C(n_499), .D(n_500), .Y(n_498) );
NAND3x1_ASAP7_75t_L g823 ( .A(n_126), .B(n_359), .C(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_325), .Y(n_126) );
AOI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_247), .B(n_259), .C(n_301), .Y(n_127) );
OAI21xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_162), .B(n_225), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_130), .A2(n_248), .B(n_253), .C(n_258), .Y(n_247) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_130), .B(n_379), .Y(n_378) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_130), .B(n_398), .Y(n_469) );
AND2x2_ASAP7_75t_L g488 ( .A(n_130), .B(n_227), .Y(n_488) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx3_ASAP7_75t_L g264 ( .A(n_131), .Y(n_264) );
AND2x2_ASAP7_75t_L g336 ( .A(n_131), .B(n_265), .Y(n_336) );
AND2x2_ASAP7_75t_L g341 ( .A(n_131), .B(n_236), .Y(n_341) );
NOR2x1_ASAP7_75t_SL g457 ( .A(n_131), .B(n_227), .Y(n_457) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_133), .B(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_133), .A2(n_230), .B(n_234), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_133), .A2(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_133), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_133), .B(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_133), .B(n_597), .Y(n_596) );
NOR3xp33_ASAP7_75t_L g598 ( .A(n_133), .B(n_145), .C(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_134), .B(n_135), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_151), .B(n_158), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B1(n_144), .B2(n_145), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_159), .B(n_184), .C(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_139), .A2(n_159), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_139), .A2(n_159), .B(n_232), .C(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g246 ( .A(n_139), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_139), .A2(n_159), .B(n_271), .C(n_272), .Y(n_270) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x2_ASAP7_75t_L g173 ( .A(n_140), .B(n_174), .Y(n_173) );
INVxp33_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g157 ( .A(n_141), .B(n_149), .Y(n_157) );
AND2x2_ASAP7_75t_L g182 ( .A(n_141), .B(n_161), .Y(n_182) );
INVx3_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g154 ( .A(n_143), .B(n_147), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_145), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g514 ( .A(n_146), .B(n_160), .Y(n_514) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B1(n_155), .B2(n_156), .Y(n_151) );
INVxp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVxp67_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g218 ( .A(n_159), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_159), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_159), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_159), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_159), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_159), .A2(n_564), .B(n_565), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_159), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_159), .A2(n_580), .B(n_581), .Y(n_579) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_205), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_164), .B(n_306), .Y(n_372) );
AND2x2_ASAP7_75t_L g489 ( .A(n_164), .B(n_330), .Y(n_489) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_189), .Y(n_164) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_165), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g278 ( .A(n_165), .Y(n_278) );
AND2x2_ASAP7_75t_L g286 ( .A(n_165), .B(n_287), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_165), .B(n_189), .Y(n_424) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_170), .B(n_186), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_166), .A2(n_167), .B1(n_192), .B2(n_197), .Y(n_191) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_166), .A2(n_170), .B(n_186), .Y(n_309) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_168), .B(n_200), .Y(n_199) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_168), .A2(n_577), .B(n_583), .Y(n_576) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx4f_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_177), .Y(n_170) );
INVx1_ASAP7_75t_L g204 ( .A(n_172), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_172), .A2(n_178), .B1(n_591), .B2(n_593), .Y(n_590) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_175), .Y(n_172) );
INVx1_ASAP7_75t_L g239 ( .A(n_173), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
BUFx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x6_ASAP7_75t_L g516 ( .A(n_176), .B(n_182), .Y(n_516) );
INVxp67_ASAP7_75t_L g202 ( .A(n_178), .Y(n_202) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_182), .Y(n_178) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_187), .Y(n_266) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_187), .A2(n_570), .B(n_574), .Y(n_569) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g376 ( .A(n_189), .B(n_214), .Y(n_376) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x4_ASAP7_75t_L g251 ( .A(n_190), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
INVx1_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_190), .B(n_309), .Y(n_333) );
AND2x2_ASAP7_75t_L g382 ( .A(n_190), .B(n_206), .Y(n_382) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_198), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g337 ( .A(n_205), .B(n_332), .Y(n_337) );
AND2x2_ASAP7_75t_L g393 ( .A(n_205), .B(n_276), .Y(n_393) );
AND2x2_ASAP7_75t_L g408 ( .A(n_205), .B(n_322), .Y(n_408) );
AND2x2_ASAP7_75t_L g445 ( .A(n_205), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g461 ( .A(n_205), .Y(n_461) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_213), .Y(n_205) );
INVx2_ASAP7_75t_L g252 ( .A(n_206), .Y(n_252) );
INVx1_ASAP7_75t_L g257 ( .A(n_206), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_206), .B(n_288), .Y(n_291) );
INVx1_ASAP7_75t_L g305 ( .A(n_206), .Y(n_305) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_206), .Y(n_315) );
INVxp67_ASAP7_75t_L g331 ( .A(n_206), .Y(n_331) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_212), .Y(n_206) );
INVx2_ASAP7_75t_SL g215 ( .A(n_207), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_207), .A2(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
AND2x4_ASAP7_75t_L g277 ( .A(n_214), .B(n_278), .Y(n_277) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_214) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_288) );
AOI21x1_ASAP7_75t_L g511 ( .A1(n_215), .A2(n_512), .B(n_517), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_217), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g258 ( .A(n_225), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_225), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_226), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_226), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_226), .B(n_294), .Y(n_437) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_226), .Y(n_475) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_235), .Y(n_226) );
INVx2_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_227), .B(n_236), .Y(n_311) );
INVx4_ASAP7_75t_L g319 ( .A(n_227), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_227), .B(n_295), .Y(n_355) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_227), .Y(n_368) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AND2x4_ASAP7_75t_L g346 ( .A(n_235), .B(n_319), .Y(n_346) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g297 ( .A(n_236), .B(n_264), .Y(n_297) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_236), .Y(n_318) );
INVx2_ASAP7_75t_L g367 ( .A(n_236), .Y(n_367) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .C(n_241), .Y(n_238) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_249), .B(n_254), .Y(n_356) );
NAND2x1_ASAP7_75t_SL g470 ( .A(n_249), .B(n_251), .Y(n_470) );
OR2x2_ASAP7_75t_L g349 ( .A(n_250), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g452 ( .A(n_250), .Y(n_452) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g342 ( .A(n_251), .B(n_277), .Y(n_342) );
AND2x2_ASAP7_75t_L g458 ( .A(n_251), .B(n_451), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_253), .A2(n_467), .B1(n_470), .B2(n_471), .C(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_254), .A2(n_411), .B1(n_413), .B2(n_415), .Y(n_410) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_255), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g324 ( .A(n_255), .Y(n_324) );
BUFx2_ASAP7_75t_L g405 ( .A(n_255), .Y(n_405) );
AND2x2_ASAP7_75t_L g375 ( .A(n_256), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_260), .B(n_279), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_274), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g348 ( .A(n_263), .Y(n_348) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_263), .B(n_474), .C(n_475), .D(n_476), .Y(n_473) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
AND2x2_ASAP7_75t_L g366 ( .A(n_264), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
INVx2_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_265), .Y(n_340) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_265), .Y(n_380) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_273), .Y(n_265) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_266), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_266), .A2(n_529), .B(n_535), .Y(n_528) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_266), .A2(n_529), .B(n_535), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g487 ( .A(n_275), .Y(n_487) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
AND2x2_ASAP7_75t_L g381 ( .A(n_277), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g481 ( .A(n_277), .B(n_482), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_289), .B2(n_292), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_281), .B(n_346), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_281), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g462 ( .A(n_281), .B(n_440), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_281), .A2(n_317), .B(n_439), .Y(n_492) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_282), .B(n_366), .Y(n_403) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_282), .Y(n_419) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g289 ( .A(n_285), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
AND2x2_ASAP7_75t_L g330 ( .A(n_287), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g451 ( .A(n_287), .B(n_308), .Y(n_451) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_288), .B(n_309), .Y(n_350) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g426 ( .A(n_291), .B(n_333), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_298), .Y(n_292) );
INVx1_ASAP7_75t_L g407 ( .A(n_293), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g302 ( .A(n_294), .B(n_303), .C(n_307), .Y(n_302) );
AND2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g374 ( .A(n_294), .B(n_317), .Y(n_374) );
AND2x2_ASAP7_75t_L g456 ( .A(n_294), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g482 ( .A(n_294), .Y(n_482) );
INVx1_ASAP7_75t_L g496 ( .A(n_294), .Y(n_496) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g299 ( .A(n_297), .B(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g455 ( .A(n_297), .Y(n_455) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g495 ( .A(n_299), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g398 ( .A(n_300), .Y(n_398) );
AO22x1_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_310), .B1(n_312), .B2(n_320), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_304), .B(n_308), .Y(n_388) );
INVx3_ASAP7_75t_L g422 ( .A(n_304), .Y(n_422) );
BUFx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx3_ASAP7_75t_L g322 ( .A(n_308), .Y(n_322) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g400 ( .A(n_309), .B(n_315), .Y(n_400) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_309), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g351 ( .A1(n_310), .A2(n_352), .A3(n_354), .B(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_311), .A2(n_328), .B1(n_334), .B2(n_337), .Y(n_327) );
AND2x2_ASAP7_75t_L g411 ( .A(n_311), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g418 ( .A(n_311), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_317), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_SL g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g347 ( .A(n_319), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_319), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g442 ( .A(n_322), .B(n_382), .Y(n_442) );
INVx1_ASAP7_75t_L g477 ( .A(n_322), .Y(n_477) );
AND2x2_ASAP7_75t_L g427 ( .A(n_323), .B(n_366), .Y(n_427) );
BUFx2_ASAP7_75t_L g472 ( .A(n_323), .Y(n_472) );
AND2x2_ASAP7_75t_L g415 ( .A(n_324), .B(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_343), .C(n_351), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_327), .B(n_338), .Y(n_326) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g404 ( .A(n_330), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_336), .B(n_346), .Y(n_369) );
AND2x2_ASAP7_75t_L g391 ( .A(n_336), .B(n_368), .Y(n_391) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_336), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
AND2x2_ASAP7_75t_L g494 ( .A(n_339), .B(n_368), .Y(n_494) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g468 ( .A(n_340), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g385 ( .A(n_341), .Y(n_385) );
AND2x2_ASAP7_75t_L g485 ( .A(n_341), .B(n_368), .Y(n_485) );
AOI21xp33_ASAP7_75t_R g343 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_345), .B(n_449), .Y(n_448) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_346), .Y(n_353) );
INVx1_ASAP7_75t_L g416 ( .A(n_350), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_352), .A2(n_370), .B1(n_384), .B2(n_386), .Y(n_383) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g384 ( .A(n_355), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_357), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_357), .B(n_464), .Y(n_463) );
NOR2xp67_ASAP7_75t_SL g499 ( .A(n_357), .B(n_430), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_428), .B(n_429), .C(n_463), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_394), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_383), .C(n_389), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_370), .B(n_373), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_365), .A2(n_404), .B1(n_407), .B2(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g441 ( .A(n_367), .Y(n_441) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g433 ( .A(n_372), .B(n_422), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_377), .B2(n_381), .Y(n_373) );
INVx1_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
AND2x4_ASAP7_75t_L g399 ( .A(n_376), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_381), .A2(n_391), .B1(n_439), .B2(n_442), .Y(n_438) );
INVxp67_ASAP7_75t_L g483 ( .A(n_382), .Y(n_483) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_385), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVxp33_ASAP7_75t_L g497 ( .A(n_388), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_409), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_406), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_401), .B2(n_404), .Y(n_396) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_410), .B(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_425), .B2(n_427), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g824 ( .A(n_431), .B(n_465), .Y(n_824) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_443), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_438), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_444), .B(n_448), .C(n_453), .D(n_459), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g486 ( .A(n_451), .B(n_487), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_458), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g500 ( .A(n_464), .Y(n_500) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR3x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_478), .C(n_490), .Y(n_465) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_483), .B(n_484), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_488), .B2(n_489), .Y(n_484) );
INVx1_ASAP7_75t_L g491 ( .A(n_489), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_493), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_497), .Y(n_493) );
CKINVDCx6p67_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
CKINVDCx11_ASAP7_75t_R g813 ( .A(n_502), .Y(n_813) );
INVx3_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g811 ( .A(n_505), .Y(n_811) );
AND3x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_669), .C(n_743), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_611), .C(n_642), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_547), .B(n_556), .C(n_584), .Y(n_507) );
AOI21x1_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_527), .B(n_545), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_509), .A2(n_645), .B1(n_651), .B2(n_654), .Y(n_644) );
AND2x2_ASAP7_75t_L g778 ( .A(n_509), .B(n_549), .Y(n_778) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
BUFx2_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
AND2x2_ASAP7_75t_L g637 ( .A(n_510), .B(n_519), .Y(n_637) );
AND2x2_ASAP7_75t_L g708 ( .A(n_510), .B(n_555), .Y(n_708) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_511), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
AND2x4_ASAP7_75t_L g601 ( .A(n_518), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g546 ( .A(n_519), .B(n_537), .Y(n_546) );
OR2x2_ASAP7_75t_L g554 ( .A(n_519), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g606 ( .A(n_519), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g653 ( .A(n_519), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_519), .B(n_555), .Y(n_661) );
AND2x2_ASAP7_75t_L g698 ( .A(n_519), .B(n_602), .Y(n_698) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_519), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_519), .B(n_536), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVx2_ASAP7_75t_L g640 ( .A(n_527), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_527), .B(n_601), .Y(n_696) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_527), .Y(n_797) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_536), .Y(n_527) );
AND2x2_ASAP7_75t_L g545 ( .A(n_528), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g622 ( .A(n_528), .B(n_537), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_528), .B(n_653), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
AND2x2_ASAP7_75t_L g689 ( .A(n_536), .B(n_606), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_536), .B(n_601), .Y(n_745) );
INVx5_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g550 ( .A(n_537), .Y(n_550) );
AND2x2_ASAP7_75t_L g616 ( .A(n_537), .B(n_607), .Y(n_616) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_537), .Y(n_636) );
AND2x4_ASAP7_75t_L g643 ( .A(n_537), .B(n_555), .Y(n_643) );
AND2x2_ASAP7_75t_SL g790 ( .A(n_537), .B(n_602), .Y(n_790) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g769 ( .A(n_545), .Y(n_769) );
INVx1_ASAP7_75t_L g711 ( .A(n_546), .Y(n_711) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g633 ( .A(n_550), .B(n_554), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_550), .B(n_602), .Y(n_726) );
AND2x2_ASAP7_75t_L g728 ( .A(n_550), .B(n_553), .Y(n_728) );
AOI32xp33_ASAP7_75t_L g794 ( .A1(n_550), .A2(n_610), .A3(n_765), .B1(n_795), .B2(n_797), .Y(n_794) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g620 ( .A(n_552), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g738 ( .A(n_552), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g761 ( .A(n_552), .B(n_622), .Y(n_761) );
AND2x2_ASAP7_75t_L g788 ( .A(n_552), .B(n_689), .Y(n_788) );
AND2x2_ASAP7_75t_L g714 ( .A(n_553), .B(n_602), .Y(n_714) );
AND2x2_ASAP7_75t_L g789 ( .A(n_553), .B(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g607 ( .A(n_555), .Y(n_607) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_567), .Y(n_557) );
NOR2x1p5_ASAP7_75t_L g647 ( .A(n_558), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
OR2x2_ASAP7_75t_L g693 ( .A(n_558), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_559), .B(n_589), .Y(n_610) );
AND2x4_ASAP7_75t_L g626 ( .A(n_559), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g657 ( .A(n_559), .B(n_569), .Y(n_657) );
OR2x2_ASAP7_75t_L g682 ( .A(n_559), .B(n_631), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_559), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_559), .B(n_569), .Y(n_717) );
INVx2_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
AND2x2_ASAP7_75t_L g748 ( .A(n_559), .B(n_588), .Y(n_748) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_559), .Y(n_772) );
INVx1_ASAP7_75t_L g777 ( .A(n_559), .Y(n_777) );
OR2x6_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
AND2x2_ASAP7_75t_L g641 ( .A(n_567), .B(n_626), .Y(n_641) );
AND2x2_ASAP7_75t_L g662 ( .A(n_567), .B(n_610), .Y(n_662) );
INVx1_ASAP7_75t_L g694 ( .A(n_567), .Y(n_694) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_575), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g587 ( .A(n_569), .Y(n_587) );
INVx2_ASAP7_75t_L g631 ( .A(n_569), .Y(n_631) );
BUFx3_ASAP7_75t_L g648 ( .A(n_569), .Y(n_648) );
AND2x2_ASAP7_75t_L g687 ( .A(n_569), .B(n_575), .Y(n_687) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_569), .Y(n_785) );
INVx2_ASAP7_75t_L g600 ( .A(n_575), .Y(n_600) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
INVx1_ASAP7_75t_L g625 ( .A(n_575), .Y(n_625) );
OR2x2_ASAP7_75t_L g630 ( .A(n_575), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g650 ( .A(n_575), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_575), .B(n_627), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_575), .B(n_733), .Y(n_732) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_601), .B(n_603), .Y(n_584) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_586), .B(n_588), .Y(n_585) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_586), .Y(n_793) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_587), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_587), .B(n_625), .Y(n_667) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_587), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_588), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_588), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g723 ( .A(n_588), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_588), .A2(n_728), .B1(n_729), .B2(n_734), .C(n_737), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_588), .B(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .Y(n_588) );
INVx3_ASAP7_75t_L g627 ( .A(n_589), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_589), .B(n_631), .Y(n_731) );
AND2x2_ASAP7_75t_L g760 ( .A(n_589), .B(n_733), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_589), .B(n_792), .Y(n_791) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_595), .Y(n_589) );
AND2x2_ASAP7_75t_L g668 ( .A(n_601), .B(n_643), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_601), .A2(n_621), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g605 ( .A(n_602), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g614 ( .A(n_602), .Y(n_614) );
OR2x2_ASAP7_75t_L g660 ( .A(n_602), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_602), .B(n_643), .Y(n_752) );
OR2x2_ASAP7_75t_L g784 ( .A(n_602), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g796 ( .A(n_602), .B(n_702), .Y(n_796) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx2_ASAP7_75t_L g674 ( .A(n_605), .Y(n_674) );
INVx3_ASAP7_75t_SL g740 ( .A(n_606), .Y(n_740) );
INVxp67_ASAP7_75t_L g690 ( .A(n_608), .Y(n_690) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g612 ( .A1(n_610), .A2(n_613), .A3(n_617), .B1(n_620), .B2(n_623), .C1(n_628), .C2(n_632), .Y(n_612) );
INVx1_ASAP7_75t_SL g701 ( .A(n_610), .Y(n_701) );
AND2x4_ASAP7_75t_L g786 ( .A(n_610), .B(n_673), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_634), .Y(n_611) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OR2x2_ASAP7_75t_L g639 ( .A(n_614), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g735 ( .A(n_614), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g763 ( .A(n_614), .B(n_616), .Y(n_763) );
AOI32xp33_ASAP7_75t_L g764 ( .A1(n_614), .A2(n_615), .A3(n_765), .B1(n_767), .B2(n_770), .Y(n_764) );
OR2x2_ASAP7_75t_L g768 ( .A(n_614), .B(n_661), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_615), .B(n_640), .C(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_SL g744 ( .A1(n_615), .A2(n_681), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g747 ( .A(n_618), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_622), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g670 ( .A1(n_626), .A2(n_630), .A3(n_639), .B1(n_671), .B2(n_674), .C1(n_675), .C2(n_676), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_626), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_626), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g649 ( .A(n_627), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g681 ( .A(n_627), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_627), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g742 ( .A(n_630), .Y(n_742) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_631), .Y(n_673) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B(n_641), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_637), .B(n_685), .Y(n_684) );
AOI322xp5_ASAP7_75t_SL g779 ( .A1(n_637), .A2(n_643), .A3(n_760), .B1(n_778), .B2(n_780), .C1(n_783), .C2(n_786), .Y(n_779) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_658), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_643), .B(n_653), .Y(n_675) );
INVx2_ASAP7_75t_SL g685 ( .A(n_643), .Y(n_685) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_SL g710 ( .A(n_649), .Y(n_710) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_650), .Y(n_680) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g755 ( .A(n_656), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g709 ( .A(n_657), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_663), .B2(n_668), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR4xp75_ASAP7_75t_L g669 ( .A(n_670), .B(n_683), .C(n_703), .D(n_719), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_678), .B(n_681), .Y(n_677) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_681), .A2(n_758), .B1(n_761), .B2(n_762), .Y(n_757) );
OR2x2_ASAP7_75t_L g722 ( .A(n_682), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g766 ( .A(n_682), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_683) );
INVx2_ASAP7_75t_L g702 ( .A(n_687), .Y(n_702) );
AND2x2_ASAP7_75t_L g759 ( .A(n_687), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B1(n_697), .B2(n_699), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g754 ( .A(n_698), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_699), .A2(n_705), .B1(n_721), .B2(n_724), .Y(n_720) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_709), .B1(n_711), .B2(n_712), .C(n_848), .Y(n_703) );
AND2x2_ASAP7_75t_SL g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g771 ( .A(n_710), .B(n_772), .Y(n_771) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g756 ( .A(n_718), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B(n_741), .Y(n_737) );
NOR3xp33_ASAP7_75t_SL g743 ( .A(n_744), .B(n_749), .C(n_773), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_764), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .B(n_755), .C(n_757), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_L g765 ( .A(n_756), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
NAND4xp25_ASAP7_75t_SL g773 ( .A(n_774), .B(n_779), .C(n_787), .D(n_794), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_778), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
OAI21xp5_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_789), .B(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx11_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
OAI22x1_ASAP7_75t_L g810 ( .A1(n_800), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AOI21xp33_ASAP7_75t_L g809 ( .A1(n_802), .A2(n_810), .B(n_814), .Y(n_809) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_835), .B(n_836), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_830), .B1(n_833), .B2(n_834), .Y(n_821) );
INVx2_ASAP7_75t_L g834 ( .A(n_822), .Y(n_834) );
XNOR2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_826), .Y(n_828) );
INVx1_ASAP7_75t_L g833 ( .A(n_830), .Y(n_833) );
INVx1_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
CKINVDCx11_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
CKINVDCx8_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
endmodule