module real_jpeg_23788_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_0),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_48),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_46),
.Y(n_147)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_3),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_32),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_51),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_3),
.B(n_48),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_51),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_6),
.B(n_66),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_233),
.Y(n_273)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_8),
.B(n_48),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_8),
.B(n_51),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_32),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_8),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_8),
.B(n_66),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_8),
.B(n_89),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_51),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_9),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_32),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_9),
.B(n_46),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_9),
.B(n_66),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_46),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_66),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_10),
.B(n_48),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_10),
.B(n_32),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_10),
.B(n_89),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_12),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_12),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_32),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_51),
.Y(n_280)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_14),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_14),
.B(n_51),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_14),
.B(n_48),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_14),
.B(n_46),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_14),
.B(n_66),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_16),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_16),
.B(n_32),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_16),
.B(n_51),
.Y(n_294)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_17),
.Y(n_112)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_17),
.Y(n_176)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_150),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_21),
.B(n_77),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_54),
.C(n_70),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_44),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_23),
.B(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_29),
.C(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_26),
.B(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_29),
.A2(n_37),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_29),
.B(n_79),
.C(n_82),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_31),
.B(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_35),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_39),
.C(n_40),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_38),
.B(n_44),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_39),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_40),
.A2(n_41),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_44),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.CI(n_50),
.CON(n_44),
.SN(n_44)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_47),
.C(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_51),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_56),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_62),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_69),
.B1(n_75),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_74),
.C(n_76),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_72),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_84),
.C(n_85),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_82),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_85),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_85),
.SN(n_85)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_87),
.C(n_88),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_90),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.C(n_108),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_91),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_92),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_94),
.B(n_100),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_97),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_104),
.B(n_108),
.Y(n_328)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.C(n_120),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_109),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_117),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_110),
.B(n_117),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_113),
.B(n_304),
.Y(n_303)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_115),
.B(n_217),
.Y(n_277)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_119),
.B(n_120),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_136),
.B2(n_137),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_148),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_330),
.C(n_331),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_320),
.C(n_321),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_306),
.C(n_307),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_283),
.C(n_284),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_253),
.C(n_254),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_227),
.C(n_228),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_188),
.C(n_200),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_171),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_166),
.C(n_171),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_161),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_167),
.B(n_169),
.C(n_170),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_172),
.B(n_180),
.C(n_181),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_187),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_199),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_193),
.B1(n_199),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_223),
.C(n_224),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_214),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.C(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_242),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_243),
.C(n_252),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_237),
.C(n_238),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_232),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_236),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_238),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.CI(n_241),
.CON(n_238),
.SN(n_238)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_251),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_249),
.C(n_251),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.C(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_265),
.C(n_268),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_260),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.CI(n_263),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_276),
.C(n_281),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_302),
.C(n_303),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_298),
.B2(n_305),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_299),
.C(n_300),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_318),
.B2(n_319),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.C(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_315),
.C(n_316),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.C(n_329),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_327),
.B2(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);


endmodule