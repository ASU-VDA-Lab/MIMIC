module fake_ibex_1558_n_1042 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1042);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1042;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_469;
wire n_323;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_439;
wire n_262;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_506;
wire n_444;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_951;
wire n_272;
wire n_881;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_874;
wire n_816;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_76),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_12),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_153),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_131),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_49),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_6),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_47),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_17),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_140),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_132),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_30),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_23),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_156),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_152),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_104),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_51),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_78),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_133),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_39),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_62),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_149),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_101),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_151),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_67),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_57),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_85),
.B(n_174),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_43),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_62),
.B(n_197),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_117),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_162),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_186),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_123),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_58),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_69),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_18),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_138),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_184),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_113),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_98),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_141),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_167),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_99),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_171),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_64),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_102),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_116),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_79),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_65),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_164),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_176),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_106),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_86),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_175),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_107),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_143),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_59),
.Y(n_299)
);

BUFx8_ASAP7_75t_SL g300 ( 
.A(n_48),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_19),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_35),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_115),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_168),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_127),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_84),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_129),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_56),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_146),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_188),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_91),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_180),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_55),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_51),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_103),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_136),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_95),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_97),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_114),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_21),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_19),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_41),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_137),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_3),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_61),
.B(n_20),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_74),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_33),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_232),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_230),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_224),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_271),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_230),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_224),
.Y(n_343)
);

OAI22x1_ASAP7_75t_R g344 ( 
.A1(n_212),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_5),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

CKINVDCx6p67_ASAP7_75t_R g350 ( 
.A(n_324),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_236),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_243),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_199),
.A2(n_68),
.B(n_66),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_270),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_199),
.A2(n_71),
.B(n_70),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_9),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_251),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_244),
.B(n_10),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_227),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_269),
.B(n_11),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_258),
.B(n_72),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_300),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_276),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_201),
.B(n_77),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g377 ( 
.A1(n_207),
.A2(n_108),
.B(n_193),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_207),
.A2(n_109),
.B(n_191),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_13),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_219),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_300),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_221),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_257),
.B(n_13),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_209),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_237),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_238),
.B(n_15),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_241),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_273),
.B(n_17),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_259),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_261),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_266),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_236),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_257),
.B(n_22),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_285),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_204),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_213),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_215),
.A2(n_112),
.B(n_187),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_25),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_216),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_293),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_217),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_247),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_277),
.B(n_27),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_223),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g408 ( 
.A1(n_228),
.A2(n_111),
.B(n_185),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_293),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_231),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_233),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_293),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_203),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_235),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_240),
.Y(n_415)
);

BUFx12f_ASAP7_75t_L g416 ( 
.A(n_209),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_206),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_249),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_391),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_211),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_417),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_334),
.B(n_409),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_389),
.B(n_254),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_389),
.B(n_256),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_384),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_335),
.A2(n_212),
.B1(n_242),
.B2(n_214),
.Y(n_435)
);

AND3x2_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_308),
.C(n_283),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_384),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_345),
.B(n_220),
.Y(n_441)
);

AO21x2_ASAP7_75t_L g442 ( 
.A1(n_357),
.A2(n_272),
.B(n_265),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_397),
.B(n_275),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_345),
.B(n_225),
.Y(n_445)
);

NOR2x1p5_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_312),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

BUFx6f_ASAP7_75t_SL g449 ( 
.A(n_366),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_341),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_346),
.B(n_279),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_341),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_366),
.Y(n_455)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

AO21x2_ASAP7_75t_L g457 ( 
.A1(n_357),
.A2(n_281),
.B(n_280),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_337),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_338),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_406),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_358),
.B(n_198),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_399),
.B(n_284),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_338),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_358),
.A2(n_327),
.B1(n_329),
.B2(n_319),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_399),
.B(n_287),
.Y(n_468)
);

CKINVDCx6p67_ASAP7_75t_R g469 ( 
.A(n_416),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_407),
.B(n_288),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_342),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_349),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_336),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_407),
.B(n_289),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_419),
.B(n_292),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_347),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_337),
.Y(n_477)
);

INVx8_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_352),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_356),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_343),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_349),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_356),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_354),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_419),
.B(n_295),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_369),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_359),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_402),
.B(n_411),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_402),
.B(n_296),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_378),
.A2(n_313),
.B(n_310),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_363),
.B(n_412),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_373),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_383),
.A2(n_394),
.B1(n_373),
.B2(n_382),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_412),
.B(n_282),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_402),
.B(n_317),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_403),
.B(n_302),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

BUFx6f_ASAP7_75t_SL g505 ( 
.A(n_404),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_383),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_403),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_411),
.B(n_200),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_360),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_403),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_381),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_415),
.B(n_202),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_404),
.B(n_305),
.Y(n_514)
);

AOI21x1_ASAP7_75t_L g515 ( 
.A1(n_378),
.A2(n_332),
.B(n_322),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_355),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_344),
.Y(n_518)
);

AND3x2_ASAP7_75t_L g519 ( 
.A(n_339),
.B(n_260),
.C(n_242),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_380),
.B(n_205),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_385),
.B(n_208),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_418),
.B(n_210),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_387),
.B(n_218),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_353),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_351),
.A2(n_214),
.B1(n_299),
.B2(n_301),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_445),
.B(n_390),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_441),
.B(n_386),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_495),
.A2(n_252),
.B1(n_253),
.B2(n_247),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_410),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_424),
.B(n_405),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_483),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_460),
.B(n_447),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_462),
.B(n_492),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_477),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

A2O1A1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_426),
.A2(n_422),
.B(n_429),
.C(n_423),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_493),
.A2(n_253),
.B1(n_290),
.B2(n_252),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_510),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_425),
.B(n_392),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_481),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_520),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_516),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_424),
.B(n_370),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_435),
.A2(n_301),
.B1(n_325),
.B2(n_307),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_465),
.B(n_331),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_370),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_453),
.B(n_371),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_521),
.B(n_372),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_453),
.B(n_374),
.Y(n_553)
);

BUFx5_ASAP7_75t_L g554 ( 
.A(n_524),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_427),
.A2(n_377),
.B(n_353),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_372),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_462),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_443),
.B(n_353),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_493),
.A2(n_290),
.B1(n_303),
.B2(n_304),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_421),
.B(n_376),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_476),
.B(n_372),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_479),
.B(n_299),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_448),
.B(n_450),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_452),
.B(n_377),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_486),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_473),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_432),
.B(n_365),
.Y(n_567)
);

BUFx8_ASAP7_75t_L g568 ( 
.A(n_512),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_226),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_451),
.A2(n_304),
.B1(n_306),
.B2(n_263),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_494),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_438),
.B(n_229),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_484),
.B(n_27),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_498),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_523),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_446),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_433),
.B(n_222),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_496),
.B(n_234),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_503),
.B(n_239),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_469),
.B(n_245),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_428),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_449),
.A2(n_309),
.B1(n_248),
.B2(n_250),
.Y(n_586)
);

NOR2xp67_ASAP7_75t_L g587 ( 
.A(n_459),
.B(n_28),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_456),
.B(n_400),
.Y(n_589)
);

BUFx6f_ASAP7_75t_SL g590 ( 
.A(n_497),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_437),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_436),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_467),
.A2(n_314),
.B1(n_262),
.B2(n_264),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_455),
.B(n_268),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_456),
.B(n_274),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_420),
.B(n_286),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_431),
.B(n_291),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_444),
.B(n_294),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_444),
.B(n_298),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_487),
.B(n_29),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_497),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_464),
.B(n_311),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_464),
.B(n_315),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_507),
.B(n_320),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_468),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_511),
.B(n_321),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_470),
.B(n_323),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_474),
.B(n_328),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_463),
.B(n_408),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_437),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_475),
.B(n_361),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_485),
.B(n_408),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_490),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_497),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_461),
.A2(n_375),
.B(n_368),
.C(n_367),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_504),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_466),
.B(n_361),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_499),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_428),
.B1(n_478),
.B2(n_518),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_558),
.A2(n_457),
.B(n_442),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_558),
.A2(n_564),
.B(n_555),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_543),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_530),
.A2(n_525),
.B1(n_519),
.B2(n_515),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_564),
.A2(n_457),
.B(n_442),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_563),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_531),
.B(n_471),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_531),
.B(n_472),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_613),
.A2(n_491),
.B(n_522),
.Y(n_634)
);

AND2x2_ASAP7_75t_SL g635 ( 
.A(n_539),
.B(n_508),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_526),
.B(n_482),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_599),
.B(n_488),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_535),
.A2(n_538),
.B(n_553),
.C(n_551),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_563),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_527),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_599),
.B(n_502),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_545),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_547),
.B(n_513),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_541),
.A2(n_534),
.B(n_573),
.C(n_544),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_560),
.B(n_29),
.Y(n_645)
);

BUFx12f_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_532),
.B(n_31),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_589),
.A2(n_489),
.B(n_509),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_534),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_566),
.B(n_31),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_540),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_590),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_580),
.B(n_32),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_579),
.B(n_34),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_592),
.B(n_36),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_37),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_562),
.B(n_38),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_528),
.B(n_39),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_546),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_569),
.B(n_40),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_572),
.B(n_40),
.Y(n_661)
);

AND2x2_ASAP7_75t_SL g662 ( 
.A(n_559),
.B(n_42),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_593),
.B(n_44),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_593),
.B(n_45),
.Y(n_665)
);

BUFx4f_ASAP7_75t_L g666 ( 
.A(n_601),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_571),
.B(n_46),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_548),
.B(n_49),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_568),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_50),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_575),
.B(n_52),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_550),
.B(n_53),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_529),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_552),
.B(n_53),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_556),
.B(n_54),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_590),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g680 ( 
.A1(n_612),
.A2(n_621),
.B(n_615),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_606),
.A2(n_517),
.B(n_454),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_548),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

AO22x1_ASAP7_75t_L g684 ( 
.A1(n_611),
.A2(n_616),
.B1(n_588),
.B2(n_581),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_582),
.B(n_57),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_577),
.B(n_58),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_614),
.A2(n_60),
.B(n_61),
.C(n_63),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_598),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_620),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_584),
.B(n_83),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_622),
.A2(n_90),
.B(n_92),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_586),
.B(n_100),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_536),
.Y(n_694)
);

BUFx8_ASAP7_75t_L g695 ( 
.A(n_537),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_587),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_600),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_585),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_594),
.B(n_147),
.Y(n_699)
);

NOR2x1p5_ASAP7_75t_L g700 ( 
.A(n_619),
.B(n_150),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_602),
.A2(n_154),
.B(n_155),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_604),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_549),
.B(n_179),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_608),
.A2(n_609),
.B(n_618),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_542),
.A2(n_163),
.B(n_165),
.C(n_166),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_170),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_585),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_640),
.B(n_631),
.Y(n_708)
);

AO31x2_ASAP7_75t_L g709 ( 
.A1(n_630),
.A2(n_617),
.A3(n_583),
.B(n_603),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_639),
.B(n_607),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_664),
.A2(n_554),
.B1(n_597),
.B2(n_605),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_649),
.B(n_596),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_642),
.Y(n_713)
);

BUFx2_ASAP7_75t_R g714 ( 
.A(n_671),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_646),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_638),
.B(n_673),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_650),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_632),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_669),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_647),
.B(n_657),
.Y(n_720)
);

OAI21x1_ASAP7_75t_SL g721 ( 
.A1(n_701),
.A2(n_704),
.B(n_661),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_633),
.B(n_636),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_656),
.B(n_637),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_652),
.B(n_679),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_641),
.B(n_693),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_651),
.B(n_628),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_645),
.A2(n_678),
.B1(n_677),
.B2(n_675),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_695),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_695),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_682),
.B(n_662),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_668),
.B(n_666),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_648),
.A2(n_681),
.B(n_680),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_670),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_665),
.B1(n_663),
.B2(n_688),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_658),
.B(n_683),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_660),
.B(n_654),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_690),
.B(n_623),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_667),
.B(n_672),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_674),
.B(n_685),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_684),
.B(n_703),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_655),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_676),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_698),
.B(n_707),
.Y(n_744)
);

AOI211x1_ASAP7_75t_L g745 ( 
.A1(n_643),
.A2(n_697),
.B(n_696),
.C(n_653),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_659),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_692),
.B(n_699),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_626),
.B(n_629),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_700),
.A2(n_702),
.B1(n_707),
.B2(n_698),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_689),
.A2(n_705),
.A3(n_687),
.B(n_691),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_706),
.B(n_686),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_694),
.Y(n_752)
);

AO31x2_ASAP7_75t_L g753 ( 
.A1(n_624),
.A2(n_630),
.A3(n_610),
.B(n_625),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_631),
.B(n_639),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_639),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_631),
.B(n_639),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_625),
.A2(n_630),
.B(n_624),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_646),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_625),
.A2(n_630),
.B(n_624),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_625),
.A2(n_630),
.B(n_624),
.Y(n_761)
);

AOI21xp33_ASAP7_75t_L g762 ( 
.A1(n_644),
.A2(n_638),
.B(n_663),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_631),
.B(n_639),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_631),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_631),
.B(n_639),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_666),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_646),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_662),
.B(n_576),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_624),
.A2(n_630),
.B(n_634),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_631),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_666),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_631),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_644),
.A2(n_639),
.B(n_631),
.C(n_638),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_625),
.A2(n_630),
.B(n_624),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_646),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_666),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_624),
.A2(n_630),
.B(n_634),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_624),
.A2(n_630),
.B(n_634),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_640),
.B(n_527),
.Y(n_782)
);

OAI21x1_ASAP7_75t_SL g783 ( 
.A1(n_644),
.A2(n_639),
.B(n_631),
.Y(n_783)
);

NAND3x1_ASAP7_75t_L g784 ( 
.A(n_668),
.B(n_351),
.C(n_539),
.Y(n_784)
);

OA22x2_ASAP7_75t_L g785 ( 
.A1(n_682),
.A2(n_539),
.B1(n_559),
.B2(n_530),
.Y(n_785)
);

AO31x2_ASAP7_75t_L g786 ( 
.A1(n_624),
.A2(n_630),
.A3(n_610),
.B(n_625),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_630),
.B(n_634),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_662),
.B(n_576),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_631),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_646),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_631),
.B(n_639),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_624),
.A2(n_630),
.A3(n_610),
.B(n_625),
.Y(n_793)
);

OAI21x1_ASAP7_75t_SL g794 ( 
.A1(n_644),
.A2(n_639),
.B(n_631),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_644),
.B(n_610),
.C(n_656),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_631),
.B(n_639),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_631),
.B(n_639),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_646),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_631),
.B(n_639),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_631),
.B(n_639),
.Y(n_801)
);

AOI21xp33_ASAP7_75t_L g802 ( 
.A1(n_644),
.A2(n_638),
.B(n_663),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_631),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_631),
.A2(n_639),
.B1(n_449),
.B2(n_493),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_627),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_631),
.A2(n_639),
.B1(n_664),
.B2(n_644),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_730),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_764),
.A2(n_803),
.B1(n_718),
.B2(n_772),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_777),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_729),
.Y(n_810)
);

OA21x2_ASAP7_75t_L g811 ( 
.A1(n_769),
.A2(n_781),
.B(n_780),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_755),
.B(n_757),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_718),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_763),
.B(n_765),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_769),
.A2(n_781),
.B(n_780),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_787),
.A2(n_760),
.B(n_758),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_733),
.A2(n_776),
.B(n_761),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_756),
.A2(n_772),
.B1(n_806),
.B2(n_778),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_768),
.B(n_788),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_731),
.A2(n_785),
.B1(n_806),
.B2(n_795),
.Y(n_820)
);

AOI22x1_ASAP7_75t_L g821 ( 
.A1(n_749),
.A2(n_721),
.B1(n_794),
.B2(n_783),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_713),
.B(n_725),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_796),
.A2(n_775),
.B(n_756),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_800),
.B(n_792),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_719),
.Y(n_825)
);

NOR2x1_ASAP7_75t_R g826 ( 
.A(n_767),
.B(n_791),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_728),
.B(n_800),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_797),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_728),
.B(n_789),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_722),
.A2(n_798),
.B1(n_801),
.B2(n_720),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_710),
.A2(n_802),
.B(n_762),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_770),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_762),
.A2(n_802),
.B(n_712),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_715),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_773),
.Y(n_835)
);

CKINVDCx14_ASAP7_75t_R g836 ( 
.A(n_799),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_714),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_728),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_790),
.Y(n_839)
);

AO32x2_ASAP7_75t_L g840 ( 
.A1(n_727),
.A2(n_711),
.A3(n_745),
.B1(n_752),
.B2(n_786),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_732),
.B(n_782),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_738),
.A2(n_735),
.B1(n_745),
.B2(n_804),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_716),
.B(n_726),
.Y(n_843)
);

INVx6_ASAP7_75t_L g844 ( 
.A(n_767),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_744),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_708),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_737),
.A2(n_740),
.B(n_739),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_759),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_791),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_753),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_724),
.B(n_779),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_717),
.A2(n_723),
.B1(n_751),
.B2(n_736),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_741),
.A2(n_784),
.B1(n_734),
.B2(n_746),
.Y(n_853)
);

OAI221xp5_ASAP7_75t_L g854 ( 
.A1(n_747),
.A2(n_742),
.B1(n_771),
.B2(n_766),
.C(n_748),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_753),
.A2(n_793),
.B(n_786),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_805),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_709),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_743),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_750),
.A2(n_774),
.B(n_796),
.Y(n_859)
);

OA21x2_ASAP7_75t_L g860 ( 
.A1(n_750),
.A2(n_780),
.B(n_769),
.Y(n_860)
);

AO21x2_ASAP7_75t_L g861 ( 
.A1(n_769),
.A2(n_781),
.B(n_780),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_728),
.B(n_646),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_774),
.A2(n_796),
.B(n_644),
.Y(n_863)
);

CKINVDCx11_ASAP7_75t_R g864 ( 
.A(n_777),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_774),
.A2(n_796),
.B(n_644),
.Y(n_865)
);

INVx3_ASAP7_75t_SL g866 ( 
.A(n_715),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_731),
.A2(n_682),
.B1(n_662),
.B2(n_785),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_731),
.A2(n_682),
.B1(n_662),
.B2(n_785),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_730),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_718),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_754),
.B(n_576),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_769),
.A2(n_781),
.B(n_780),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_715),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_718),
.A2(n_764),
.B1(n_803),
.B2(n_722),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_850),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_845),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_829),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_813),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_855),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_827),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_845),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_813),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_870),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_858),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_829),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_870),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_856),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_856),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_858),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_822),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_864),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_823),
.B(n_824),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_847),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_832),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_828),
.B(n_830),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_851),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_871),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_835),
.Y(n_898)
);

INVxp33_ASAP7_75t_L g899 ( 
.A(n_826),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_812),
.B(n_814),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_863),
.A2(n_865),
.B(n_833),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_843),
.B(n_831),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_820),
.B(n_818),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_853),
.A2(n_874),
.B(n_842),
.C(n_854),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_840),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_867),
.A2(n_868),
.B1(n_820),
.B2(n_846),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_818),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_816),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_857),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_907),
.B(n_860),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_895),
.B(n_859),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_SL g912 ( 
.A1(n_895),
.A2(n_821),
.B1(n_837),
.B2(n_839),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_875),
.B(n_860),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_890),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_909),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_902),
.B(n_903),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_887),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_887),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_878),
.B(n_861),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_902),
.B(n_808),
.Y(n_920)
);

INVx4_ASAP7_75t_R g921 ( 
.A(n_877),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_903),
.B(n_808),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_901),
.B(n_852),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_905),
.B(n_872),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_901),
.B(n_852),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_893),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_888),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

NOR2x1_ASAP7_75t_L g929 ( 
.A(n_877),
.B(n_885),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_900),
.B(n_894),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_879),
.B(n_817),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_877),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_915),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_928),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_932),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_915),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_911),
.B(n_882),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_929),
.B(n_880),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_916),
.B(n_883),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_926),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_930),
.B(n_807),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_927),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_924),
.B(n_811),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_911),
.B(n_886),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_916),
.B(n_906),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_931),
.B(n_913),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_919),
.B(n_892),
.Y(n_948)
);

OAI221xp5_ASAP7_75t_L g949 ( 
.A1(n_923),
.A2(n_867),
.B1(n_868),
.B2(n_904),
.C(n_900),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_919),
.B(n_815),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_946),
.B(n_910),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_910),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_933),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_937),
.B(n_914),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_934),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_939),
.B(n_937),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_933),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_936),
.Y(n_958)
);

OR2x6_ASAP7_75t_SL g959 ( 
.A(n_944),
.B(n_922),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_944),
.B(n_917),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_939),
.B(n_918),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_940),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_950),
.B(n_918),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_935),
.B(n_884),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_935),
.B(n_884),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_935),
.B(n_921),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_946),
.B(n_910),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_946),
.B(n_935),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_940),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_953),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_951),
.B(n_946),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_959),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_955),
.Y(n_974)
);

AOI32xp33_ASAP7_75t_L g975 ( 
.A1(n_968),
.A2(n_899),
.A3(n_912),
.B1(n_941),
.B2(n_929),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_957),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_954),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_958),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_962),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_956),
.B(n_945),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_961),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_969),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_959),
.B(n_945),
.Y(n_984)
);

AOI32xp33_ASAP7_75t_L g985 ( 
.A1(n_984),
.A2(n_968),
.A3(n_912),
.B1(n_967),
.B2(n_952),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_974),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_949),
.C(n_947),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_981),
.B(n_960),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_982),
.A2(n_968),
.B1(n_949),
.B2(n_952),
.Y(n_989)
);

NOR2x1p5_ASAP7_75t_L g990 ( 
.A(n_975),
.B(n_966),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_973),
.A2(n_967),
.B(n_951),
.Y(n_991)
);

AOI21xp33_ASAP7_75t_L g992 ( 
.A1(n_978),
.A2(n_925),
.B(n_923),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_977),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_971),
.A2(n_964),
.B1(n_960),
.B2(n_922),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_971),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_974),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_970),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_970),
.B(n_942),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_976),
.B(n_943),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_990),
.A2(n_983),
.B1(n_976),
.B2(n_925),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_989),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_988),
.B(n_979),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_L g1003 ( 
.A(n_987),
.B(n_849),
.C(n_825),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_997),
.Y(n_1004)
);

NAND4xp25_ASAP7_75t_L g1005 ( 
.A(n_985),
.B(n_862),
.C(n_869),
.D(n_819),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_993),
.Y(n_1006)
);

NAND2x1_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_921),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_1000),
.B(n_1001),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_1005),
.A2(n_1007),
.B(n_985),
.Y(n_1009)
);

OAI221xp5_ASAP7_75t_L g1010 ( 
.A1(n_1006),
.A2(n_994),
.B1(n_991),
.B2(n_995),
.C(n_965),
.Y(n_1010)
);

NOR4xp25_ASAP7_75t_L g1011 ( 
.A(n_1004),
.B(n_809),
.C(n_894),
.D(n_898),
.Y(n_1011)
);

OAI321xp33_ASAP7_75t_L g1012 ( 
.A1(n_1002),
.A2(n_965),
.A3(n_920),
.B1(n_938),
.B2(n_948),
.C(n_950),
.Y(n_1012)
);

OAI211xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1000),
.A2(n_864),
.B(n_836),
.C(n_930),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1001),
.B(n_998),
.Y(n_1014)
);

AOI322xp5_ASAP7_75t_L g1015 ( 
.A1(n_1001),
.A2(n_891),
.A3(n_986),
.B1(n_996),
.B2(n_947),
.C1(n_897),
.C2(n_980),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1014),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_848),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_1010),
.B(n_834),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1011),
.A2(n_836),
.B(n_834),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_979),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_1013),
.B(n_848),
.C(n_810),
.Y(n_1021)
);

NAND3x1_ASAP7_75t_L g1022 ( 
.A(n_1019),
.B(n_1008),
.C(n_1012),
.Y(n_1022)
);

NOR4xp25_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_881),
.C(n_876),
.D(n_841),
.Y(n_1023)
);

NOR3x1_ASAP7_75t_L g1024 ( 
.A(n_1020),
.B(n_866),
.C(n_896),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_1016),
.B(n_838),
.C(n_884),
.Y(n_1025)
);

NAND4xp75_ASAP7_75t_L g1026 ( 
.A(n_1018),
.B(n_1021),
.C(n_896),
.D(n_876),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1016),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_1023),
.B(n_873),
.C(n_866),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1027),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1026),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_889),
.C(n_884),
.Y(n_1031)
);

AND2x4_ASAP7_75t_SL g1032 ( 
.A(n_1022),
.B(n_873),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_1032),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_851),
.Y(n_1034)
);

XNOR2xp5_ASAP7_75t_L g1035 ( 
.A(n_1033),
.B(n_1030),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1035),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1036),
.Y(n_1037)
);

XNOR2xp5_ASAP7_75t_L g1038 ( 
.A(n_1037),
.B(n_1034),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1038),
.Y(n_1039)
);

OA21x2_ASAP7_75t_L g1040 ( 
.A1(n_1039),
.A2(n_1029),
.B(n_1031),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_1040),
.B(n_844),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_1041),
.A2(n_844),
.B1(n_1024),
.B2(n_851),
.Y(n_1042)
);


endmodule