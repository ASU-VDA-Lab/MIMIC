module fake_jpeg_18771_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_58),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_53),
.B1(n_66),
.B2(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_79),
.B1(n_78),
.B2(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_52),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_106),
.B1(n_87),
.B2(n_72),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_67),
.B1(n_57),
.B2(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_61),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_60),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx11_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_114),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_68),
.B1(n_73),
.B2(n_70),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_63),
.B1(n_59),
.B2(n_55),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_49),
.B1(n_48),
.B2(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_120),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_51),
.B(n_18),
.C(n_19),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_20),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_17),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_16),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_25),
.B(n_43),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_132),
.B(n_133),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_0),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_128),
.C(n_1),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_21),
.C(n_41),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_112),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_117),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_14),
.B(n_39),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_139),
.C(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_141),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_142),
.CI(n_140),
.CON(n_145),
.SN(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_145),
.C(n_143),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_130),
.B(n_123),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_130),
.C(n_10),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_31),
.B(n_29),
.C(n_23),
.Y(n_150)
);

OA21x2_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_2),
.B(n_3),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_7),
.C(n_4),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_6),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_6),
.Y(n_154)
);


endmodule