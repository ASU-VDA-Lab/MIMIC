module fake_jpeg_29516_n_361 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_361);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_33),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_56),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_44),
.B(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_33),
.B1(n_22),
.B2(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_74),
.B1(n_21),
.B2(n_40),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_31),
.B1(n_35),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_31),
.B1(n_35),
.B2(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_31),
.B1(n_34),
.B2(n_30),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_33),
.B1(n_20),
.B2(n_27),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_21),
.B(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_34),
.B1(n_41),
.B2(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_22),
.B1(n_38),
.B2(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_81),
.Y(n_88)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_34),
.B1(n_41),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_41),
.B1(n_55),
.B2(n_47),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_59),
.B1(n_74),
.B2(n_67),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_103),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_46),
.C(n_56),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_91),
.C(n_50),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_51),
.B1(n_49),
.B2(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_86),
.A2(n_90),
.B1(n_93),
.B2(n_95),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_68),
.B1(n_45),
.B2(n_65),
.Y(n_131)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_53),
.C(n_47),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_22),
.B1(n_38),
.B2(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_101),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_22),
.B1(n_38),
.B2(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_102),
.A2(n_108),
.B1(n_110),
.B2(n_114),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_50),
.B1(n_78),
.B2(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_119),
.Y(n_149)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_36),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_68),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_65),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_90),
.B1(n_121),
.B2(n_65),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_151),
.Y(n_169)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_36),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_39),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_39),
.B1(n_50),
.B2(n_45),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_89),
.B1(n_109),
.B2(n_113),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_32),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_106),
.C(n_91),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_181),
.C(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_82),
.B1(n_95),
.B2(n_92),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_162),
.B1(n_177),
.B2(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_86),
.B1(n_108),
.B2(n_96),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_176),
.B1(n_166),
.B2(n_165),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_106),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_175),
.B(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_133),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_106),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_99),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_171),
.A2(n_180),
.B(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_83),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_179),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_152),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_104),
.CI(n_120),
.CON(n_174),
.SN(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_112),
.B(n_107),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_100),
.B1(n_94),
.B2(n_110),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_125),
.B1(n_147),
.B2(n_129),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_127),
.A2(n_119),
.B1(n_110),
.B2(n_80),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_116),
.B(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_111),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_32),
.B(n_1),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_80),
.B1(n_45),
.B2(n_89),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_145),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_184),
.B(n_189),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_195),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_194),
.B(n_0),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_156),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_198),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_132),
.B(n_154),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_132),
.B(n_140),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_158),
.B(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_140),
.B1(n_153),
.B2(n_130),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_197),
.B1(n_202),
.B2(n_203),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_129),
.C(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_125),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_211),
.Y(n_215)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_183),
.Y(n_201)
);

INVx11_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_153),
.B1(n_124),
.B2(n_135),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_146),
.B(n_137),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_135),
.C(n_137),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_212),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_164),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_146),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_153),
.C(n_146),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_192),
.Y(n_223)
);

INVx2_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_178),
.B(n_160),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_233),
.B(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_162),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_236),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_163),
.B(n_182),
.C(n_183),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_161),
.B(n_157),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_1),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_240),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_197),
.B1(n_184),
.B2(n_213),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_191),
.B(n_13),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_206),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_189),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_249),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_193),
.B1(n_191),
.B2(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_193),
.B1(n_229),
.B2(n_225),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_265),
.B1(n_233),
.B2(n_237),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_212),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_250),
.A2(n_252),
.B1(n_266),
.B2(n_270),
.Y(n_286)
);

XNOR2x2_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_185),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_231),
.B(n_228),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_233),
.B1(n_222),
.B2(n_218),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_207),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_255),
.C(n_267),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_198),
.Y(n_255)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_185),
.B1(n_40),
.B2(n_122),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_40),
.B1(n_45),
.B2(n_42),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_57),
.C(n_42),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_269),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_42),
.B1(n_11),
.B2(n_18),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_221),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_277),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_214),
.B(n_222),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_281),
.B(n_262),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_239),
.C(n_234),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_282),
.C(n_246),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_220),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_245),
.A2(n_216),
.B(n_217),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_215),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_215),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_216),
.B(n_219),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_261),
.B(n_264),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_254),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_220),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_219),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_251),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_291),
.B1(n_270),
.B2(n_266),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_248),
.A2(n_232),
.B1(n_243),
.B2(n_13),
.Y(n_291)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_280),
.B1(n_279),
.B2(n_297),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_249),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_296),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_280),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_265),
.B1(n_250),
.B2(n_256),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_300),
.A2(n_306),
.B1(n_289),
.B2(n_291),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_267),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_307),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_309),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_256),
.B1(n_260),
.B2(n_262),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_284),
.A2(n_269),
.B(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_8),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_271),
.B(n_8),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_279),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_299),
.A2(n_271),
.B1(n_303),
.B2(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_318),
.B1(n_300),
.B2(n_297),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_319),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_317),
.A2(n_293),
.B1(n_10),
.B2(n_14),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_272),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_278),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_323),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_322),
.B(n_302),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_298),
.A2(n_285),
.B(n_274),
.C(n_281),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_296),
.B(n_272),
.Y(n_323)
);

AOI321xp33_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_275),
.A3(n_287),
.B1(n_276),
.B2(n_288),
.C(n_14),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_6),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_331),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_324),
.A2(n_302),
.B(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_322),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_312),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.C(n_331),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_334),
.A2(n_336),
.B(n_315),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_326),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_316),
.B(n_311),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_330),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_339),
.B(n_340),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_327),
.A2(n_315),
.B(n_322),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_341),
.A2(n_345),
.B(n_346),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_342),
.B(n_15),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_322),
.B(n_326),
.Y(n_345)
);

AOI322xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_333),
.A3(n_328),
.B1(n_337),
.B2(n_57),
.C1(n_10),
.C2(n_7),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g357 ( 
.A1(n_347),
.A2(n_348),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_343),
.C2(n_352),
.Y(n_357)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_57),
.A3(n_15),
.B1(n_7),
.B2(n_4),
.C1(n_1),
.C2(n_3),
.Y(n_348)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_57),
.B(n_3),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_2),
.B(n_4),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_355),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_349),
.B(n_4),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_356),
.C(n_5),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_358),
.Y(n_361)
);


endmodule