module real_aes_11248_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_92;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_0), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_1), .B(n_56), .Y(n_596) );
AND2x2_ASAP7_75t_L g606 ( .A(n_1), .B(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_1), .Y(n_650) );
INVx1_ASAP7_75t_L g675 ( .A(n_1), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_2), .B(n_157), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_3), .B(n_140), .Y(n_188) );
INVx2_ASAP7_75t_L g521 ( .A(n_4), .Y(n_521) );
OR2x2_ASAP7_75t_L g691 ( .A(n_4), .B(n_519), .Y(n_691) );
INVx1_ASAP7_75t_L g523 ( .A(n_5), .Y(n_523) );
BUFx2_ASAP7_75t_L g530 ( .A(n_5), .Y(n_530) );
BUFx2_ASAP7_75t_L g556 ( .A(n_5), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_6), .B(n_120), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_7), .B(n_104), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_8), .B(n_104), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_9), .Y(n_492) );
AND2x2_ASAP7_75t_L g231 ( .A(n_10), .B(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_11), .Y(n_585) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_13), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_14), .B(n_124), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_15), .A2(n_33), .B1(n_572), .B2(n_579), .Y(n_571) );
INVx1_ASAP7_75t_L g677 ( .A(n_15), .Y(n_677) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_16), .Y(n_489) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_17), .B(n_172), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_18), .B(n_172), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_19), .A2(n_504), .B1(n_699), .B2(n_719), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_19), .Y(n_719) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_21), .Y(n_198) );
INVx1_ASAP7_75t_L g501 ( .A(n_22), .Y(n_501) );
INVx1_ASAP7_75t_L g519 ( .A(n_23), .Y(n_519) );
INVx1_ASAP7_75t_L g528 ( .A(n_23), .Y(n_528) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_24), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_25), .B(n_139), .Y(n_175) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_26), .A2(n_40), .B1(n_669), .B2(n_670), .C(n_672), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_26), .A2(n_44), .B1(n_695), .B2(n_697), .Y(n_694) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_27), .A2(n_47), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_28), .A2(n_114), .B(n_237), .C(n_238), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_29), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_30), .B(n_118), .Y(n_133) );
NAND2xp33_ASAP7_75t_L g158 ( .A(n_31), .B(n_152), .Y(n_158) );
AND2x6_ASAP7_75t_L g84 ( .A(n_32), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_32), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_32), .B(n_704), .Y(n_735) );
INVx1_ASAP7_75t_L g681 ( .A(n_33), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_34), .B(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_34), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_35), .B(n_218), .Y(n_217) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_36), .B(n_152), .Y(n_189) );
INVx1_ASAP7_75t_L g485 ( .A(n_37), .Y(n_485) );
INVx1_ASAP7_75t_L g85 ( .A(n_38), .Y(n_85) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_38), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_39), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g687 ( .A1(n_40), .A2(n_52), .B1(n_688), .B2(n_692), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_41), .B(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_42), .Y(n_131) );
AND2x2_ASAP7_75t_L g240 ( .A(n_43), .B(n_124), .Y(n_240) );
INVx1_ASAP7_75t_L g662 ( .A(n_44), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_45), .B(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_45), .Y(n_731) );
INVx2_ASAP7_75t_L g600 ( .A(n_46), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_48), .Y(n_174) );
NAND2xp33_ASAP7_75t_L g110 ( .A(n_49), .B(n_90), .Y(n_110) );
INVx1_ASAP7_75t_L g565 ( .A(n_50), .Y(n_565) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_50), .A2(n_655), .B(n_660), .C(n_676), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_51), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g667 ( .A(n_52), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_53), .Y(n_497) );
BUFx10_ASAP7_75t_L g713 ( .A(n_54), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_55), .B(n_89), .Y(n_215) );
INVx2_ASAP7_75t_L g607 ( .A(n_56), .Y(n_607) );
INVx1_ASAP7_75t_L g651 ( .A(n_56), .Y(n_651) );
NAND2xp33_ASAP7_75t_L g119 ( .A(n_57), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g561 ( .A(n_58), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_58), .A2(n_621), .B1(n_624), .B2(n_637), .C(n_652), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_59), .A2(n_77), .B1(n_547), .B2(n_550), .Y(n_546) );
INVx1_ASAP7_75t_L g630 ( .A(n_59), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_60), .B(n_172), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_61), .Y(n_239) );
INVx2_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_63), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_64), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_65), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_66), .B(n_143), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_67), .Y(n_184) );
INVx1_ASAP7_75t_L g230 ( .A(n_68), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_69), .Y(n_200) );
AND2x2_ASAP7_75t_L g209 ( .A(n_70), .B(n_104), .Y(n_209) );
INVx2_ASAP7_75t_L g601 ( .A(n_71), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_72), .A2(n_74), .B1(n_567), .B2(n_570), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_72), .A2(n_74), .B1(n_604), .B2(n_612), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_73), .B(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g513 ( .A(n_75), .Y(n_513) );
INVx1_ASAP7_75t_L g537 ( .A(n_75), .Y(n_537) );
BUFx3_ASAP7_75t_L g514 ( .A(n_76), .Y(n_514) );
INVx1_ASAP7_75t_L g539 ( .A(n_76), .Y(n_539) );
INVx1_ASAP7_75t_L g636 ( .A(n_77), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_95), .B(n_479), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx8_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_83), .A2(n_196), .B(n_202), .Y(n_195) );
NOR2xp67_ASAP7_75t_L g225 ( .A(n_83), .B(n_226), .Y(n_225) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
BUFx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g733 ( .A1(n_87), .A2(n_734), .B(n_735), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
INVx2_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_91), .Y(n_120) );
INVx2_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_91), .Y(n_207) );
INVx1_ASAP7_75t_L g234 ( .A(n_91), .Y(n_234) );
OAI21xp33_ASAP7_75t_L g202 ( .A1(n_92), .A2(n_203), .B(n_205), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_92), .A2(n_214), .B(n_215), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_93), .Y(n_92) );
INVx3_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_93), .A2(n_156), .B(n_158), .Y(n_155) );
BUFx2_ASAP7_75t_L g235 ( .A(n_93), .Y(n_235) );
BUFx12f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx5_ASAP7_75t_L g114 ( .A(n_94), .Y(n_114) );
INVx5_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_94), .A2(n_131), .B(n_132), .C(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
BUFx2_ASAP7_75t_SL g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NAND4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_335), .C(n_400), .D(n_450), .Y(n_98) );
NOR3x1_ASAP7_75t_L g99 ( .A(n_100), .B(n_266), .C(n_303), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_SL g100 ( .A1(n_101), .A2(n_161), .B(n_177), .C(n_241), .Y(n_100) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_101), .A2(n_281), .B(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_SL g101 ( .A(n_102), .B(n_126), .Y(n_101) );
AND2x2_ASAP7_75t_L g353 ( .A(n_102), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_102), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_103), .B(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_103), .Y(n_432) );
INVx2_ASAP7_75t_L g448 ( .A(n_103), .Y(n_448) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_108), .B(n_123), .Y(n_103) );
BUFx4f_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
INVx3_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_104), .A2(n_108), .B(n_123), .Y(n_163) );
INVx4_ASAP7_75t_L g194 ( .A(n_104), .Y(n_194) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_104), .A2(n_108), .B(n_123), .Y(n_257) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_115), .B(n_122), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_111), .B(n_113), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_113), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_113), .A2(n_188), .B(n_189), .Y(n_187) );
CKINVDCx6p67_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g201 ( .A(n_114), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B(n_121), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g199 ( .A(n_117), .B(n_200), .Y(n_199) );
INVx5_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
INVx2_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_120), .B(n_198), .Y(n_197) );
INVx2_ASAP7_75t_SL g218 ( .A(n_120), .Y(n_218) );
AOI21x1_ASAP7_75t_L g150 ( .A1(n_121), .A2(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g220 ( .A(n_121), .Y(n_220) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_122), .A2(n_130), .B(n_134), .Y(n_129) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_122), .A2(n_169), .B(n_173), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_122), .A2(n_183), .B(n_187), .Y(n_182) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_122), .A2(n_213), .B(n_216), .Y(n_212) );
BUFx5_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g311 ( .A(n_126), .Y(n_311) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_145), .Y(n_126) );
AND2x2_ASAP7_75t_L g245 ( .A(n_127), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g360 ( .A(n_127), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_127), .B(n_249), .Y(n_367) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_142), .Y(n_127) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_128), .A2(n_168), .B(n_176), .Y(n_167) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_128), .A2(n_182), .B(n_190), .Y(n_181) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_128), .A2(n_129), .B(n_142), .Y(n_253) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_128), .A2(n_168), .B(n_176), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_138), .C(n_141), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g173 ( .A1(n_136), .A2(n_141), .B(n_174), .C(n_175), .Y(n_173) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
INVx2_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_141), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g165 ( .A(n_145), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g280 ( .A(n_145), .Y(n_280) );
AND2x2_ASAP7_75t_L g329 ( .A(n_145), .B(n_167), .Y(n_329) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_160), .Y(n_146) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_147), .A2(n_212), .B(n_221), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_149), .B(n_160), .Y(n_246) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_155), .B(n_159), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_152), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
OR2x2_ASAP7_75t_L g320 ( .A(n_162), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g372 ( .A(n_162), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g382 ( .A(n_162), .B(n_376), .Y(n_382) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_SL g248 ( .A(n_163), .Y(n_248) );
BUFx2_ASAP7_75t_L g293 ( .A(n_163), .Y(n_293) );
INVx1_ASAP7_75t_SL g411 ( .A(n_163), .Y(n_411) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g291 ( .A(n_165), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g442 ( .A(n_165), .B(n_327), .Y(n_442) );
INVx2_ASAP7_75t_L g249 ( .A(n_166), .Y(n_249) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_172), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI221xp5_ASAP7_75t_SL g433 ( .A1(n_178), .A2(n_434), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_433) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
INVxp67_ASAP7_75t_L g368 ( .A(n_179), .Y(n_368) );
AND2x4_ASAP7_75t_L g371 ( .A(n_179), .B(n_348), .Y(n_371) );
OR2x2_ASAP7_75t_L g393 ( .A(n_179), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_180), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g333 ( .A(n_180), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_180), .B(n_288), .Y(n_350) );
AND2x2_ASAP7_75t_L g361 ( .A(n_180), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_180), .B(n_348), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_180), .B(n_192), .Y(n_430) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
AND2x2_ASAP7_75t_L g445 ( .A(n_181), .B(n_271), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_191), .A2(n_326), .B1(n_353), .B2(n_355), .Y(n_352) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_210), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_192), .B(n_273), .Y(n_458) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_SL g302 ( .A(n_193), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_193), .B(n_309), .Y(n_308) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_209), .Y(n_193) );
INVx3_ASAP7_75t_L g226 ( .A(n_194), .Y(n_226) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_194), .A2(n_195), .B(n_209), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_199), .B(n_201), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_198), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_198), .Y(n_502) );
NOR2xp33_ASAP7_75t_SL g205 ( .A(n_206), .B(n_208), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_206), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g431 ( .A(n_210), .Y(n_431) );
AND2x4_ASAP7_75t_L g444 ( .A(n_210), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
AND2x2_ASAP7_75t_L g261 ( .A(n_211), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g274 ( .A(n_211), .Y(n_274) );
OR2x2_ASAP7_75t_L g284 ( .A(n_211), .B(n_271), .Y(n_284) );
INVx1_ASAP7_75t_L g309 ( .A(n_211), .Y(n_309) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_211), .Y(n_334) );
INVx1_ASAP7_75t_L g362 ( .A(n_211), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_219), .B(n_220), .Y(n_216) );
INVx2_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AND2x2_ASAP7_75t_L g270 ( .A(n_223), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g343 ( .A(n_223), .B(n_302), .Y(n_343) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_240), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_236), .Y(n_227) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_231), .B(n_235), .Y(n_228) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_250), .B(n_260), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2x1_ASAP7_75t_SL g340 ( .A(n_244), .B(n_247), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_244), .A2(n_427), .B(n_429), .C(n_432), .Y(n_426) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
BUFx2_ASAP7_75t_L g461 ( .A(n_246), .Y(n_461) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_247), .Y(n_289) );
INVx1_ASAP7_75t_L g405 ( .A(n_247), .Y(n_405) );
OR2x2_ASAP7_75t_L g420 ( .A(n_247), .B(n_421), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_247), .A2(n_444), .B(n_461), .C(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_248), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g277 ( .A(n_249), .B(n_257), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_249), .B(n_280), .Y(n_297) );
INVx1_ASAP7_75t_L g322 ( .A(n_249), .Y(n_322) );
AND2x2_ASAP7_75t_L g471 ( .A(n_249), .B(n_257), .Y(n_471) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
AND2x2_ASAP7_75t_L g470 ( .A(n_251), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_SL g278 ( .A(n_252), .B(n_279), .Y(n_278) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_252), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_252), .B(n_258), .Y(n_373) );
BUFx2_ASAP7_75t_L g435 ( .A(n_252), .Y(n_435) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
INVx1_ASAP7_75t_L g328 ( .A(n_253), .Y(n_328) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
AND2x2_ASAP7_75t_L g465 ( .A(n_254), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_257), .B(n_360), .Y(n_392) );
INVx1_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g354 ( .A(n_259), .B(n_280), .Y(n_354) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g298 ( .A(n_261), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g318 ( .A(n_261), .B(n_270), .Y(n_318) );
AND2x4_ASAP7_75t_L g342 ( .A(n_261), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_261), .B(n_331), .Y(n_453) );
OR2x2_ASAP7_75t_L g273 ( .A(n_262), .B(n_274), .Y(n_273) );
BUFx3_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g316 ( .A(n_264), .B(n_284), .Y(n_316) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g395 ( .A(n_265), .B(n_271), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_275), .B1(n_281), .B2(n_289), .C(n_290), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_272), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_268), .A2(n_458), .B(n_469), .C(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_269), .A2(n_441), .B1(n_443), .B2(n_446), .Y(n_440) );
OR2x2_ASAP7_75t_L g478 ( .A(n_269), .B(n_333), .Y(n_478) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g386 ( .A(n_270), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_270), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_272), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g387 ( .A(n_273), .Y(n_387) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_273), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
AND2x4_ASAP7_75t_L g407 ( .A(n_276), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g436 ( .A(n_277), .Y(n_436) );
INVx1_ASAP7_75t_L g366 ( .A(n_279), .Y(n_366) );
AND2x4_ASAP7_75t_L g412 ( .A(n_279), .B(n_327), .Y(n_412) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g348 ( .A(n_284), .Y(n_348) );
OR2x2_ASAP7_75t_L g425 ( .A(n_284), .B(n_306), .Y(n_425) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g462 ( .A(n_286), .B(n_308), .Y(n_462) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_288), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_294), .B(n_298), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g385 ( .A(n_293), .B(n_329), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_294), .A2(n_419), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_418) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_296), .Y(n_408) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_296), .Y(n_421) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVxp67_ASAP7_75t_L g378 ( .A(n_300), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g402 ( .A1(n_300), .A2(n_318), .A3(n_403), .B1(n_406), .B2(n_407), .C1(n_409), .C2(n_413), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_300), .B(n_361), .Y(n_438) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_317), .C(n_323), .Y(n_303) );
AOI32xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .A3(n_311), .B1(n_312), .B2(n_315), .Y(n_304) );
OAI21xp33_ASAP7_75t_SL g317 ( .A1(n_305), .A2(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g428 ( .A(n_306), .Y(n_428) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g423 ( .A(n_308), .B(n_350), .Y(n_423) );
NAND2x1_ASAP7_75t_SL g404 ( .A(n_311), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
OR2x2_ASAP7_75t_L g459 ( .A(n_313), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g383 ( .A(n_314), .Y(n_383) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g355 ( .A(n_316), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_318), .A2(n_407), .B1(n_412), .B2(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g439 ( .A(n_321), .Y(n_439) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g324 ( .A(n_325), .B(n_330), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g454 ( .A(n_326), .B(n_432), .Y(n_454) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g466 ( .A(n_327), .Y(n_466) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g346 ( .A(n_329), .Y(n_346) );
AND2x2_ASAP7_75t_SL g358 ( .A(n_329), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g449 ( .A(n_329), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_330), .A2(n_384), .B1(n_441), .B2(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g369 ( .A(n_331), .Y(n_369) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_356), .C(n_379), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_351), .Y(n_337) );
OAI21xp33_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_341), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x2_ASAP7_75t_L g390 ( .A(n_345), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g463 ( .A(n_345), .Y(n_463) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g375 ( .A(n_359), .Y(n_375) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_361), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g469 ( .A(n_361), .Y(n_469) );
OAI322xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_368), .A3(n_369), .B1(n_370), .B2(n_372), .C1(n_374), .C2(n_377), .Y(n_363) );
INVx1_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g475 ( .A(n_372), .Y(n_475) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_386), .B(n_388), .Y(n_379) );
NAND4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .C(n_383), .D(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B1(n_396), .B2(n_397), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g416 ( .A(n_395), .B(n_398), .Y(n_416) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g447 ( .A(n_399), .B(n_448), .Y(n_447) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_417), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_415), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_433), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
NAND2xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_449), .Y(n_446) );
AND3x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .C(n_472), .Y(n_450) );
NAND2xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_467), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_462), .B2(n_463), .C(n_464), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g474 ( .A(n_460), .Y(n_474) );
INVx2_ASAP7_75t_L g473 ( .A(n_462), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_475), .B2(n_476), .C(n_477), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_700), .B1(n_718), .B2(n_720), .C(n_724), .Y(n_479) );
XOR2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_494), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_481) );
INVx1_ASAP7_75t_L g493 ( .A(n_482), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_489), .B2(n_490), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_485), .Y(n_488) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_489), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_504), .B2(n_699), .Y(n_494) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_503), .Y(n_496) );
INVx1_ASAP7_75t_L g503 ( .A(n_497), .Y(n_503) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g699 ( .A(n_504), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_504), .A2(n_699), .B1(n_729), .B2(n_730), .Y(n_728) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND4x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_584), .C(n_602), .D(n_686), .Y(n_505) );
NOR3xp33_ASAP7_75t_SL g506 ( .A(n_507), .B(n_524), .C(n_571), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x4_ASAP7_75t_L g549 ( .A(n_513), .B(n_539), .Y(n_549) );
INVx2_ASAP7_75t_L g583 ( .A(n_513), .Y(n_583) );
AND2x4_ASAP7_75t_L g553 ( .A(n_514), .B(n_537), .Y(n_553) );
INVx2_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g578 ( .A(n_516), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_516), .B(n_580), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
AND2x2_ASAP7_75t_L g588 ( .A(n_517), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g716 ( .A(n_517), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g557 ( .A(n_520), .B(n_528), .Y(n_557) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g527 ( .A(n_521), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g690 ( .A(n_523), .B(n_691), .Y(n_690) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_525), .A2(n_531), .B1(n_554), .B2(n_558), .Y(n_524) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g709 ( .A(n_527), .Y(n_709) );
INVx2_ASAP7_75t_L g591 ( .A(n_529), .Y(n_591) );
BUFx2_ASAP7_75t_L g685 ( .A(n_529), .Y(n_685) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_540), .B1(n_541), .B2(n_542), .C(n_546), .Y(n_531) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g560 ( .A(n_535), .Y(n_560) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g545 ( .A(n_536), .B(n_538), .Y(n_545) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_540), .A2(n_541), .B1(n_638), .B2(n_642), .C(n_646), .Y(n_637) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g564 ( .A(n_545), .Y(n_564) );
INVx2_ASAP7_75t_L g693 ( .A(n_545), .Y(n_693) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g698 ( .A(n_548), .Y(n_698) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_549), .Y(n_569) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_552), .Y(n_570) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g689 ( .A(n_553), .Y(n_689) );
INVx4_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x4_ASAP7_75t_L g587 ( .A(n_556), .B(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_561), .B1(n_562), .B2(n_565), .C(n_566), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g696 ( .A(n_560), .Y(n_696) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
INVx1_ASAP7_75t_L g711 ( .A(n_574), .Y(n_711) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g717 ( .A(n_575), .Y(n_717) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g589 ( .A(n_577), .B(n_583), .Y(n_589) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x6_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
AND2x2_ASAP7_75t_L g678 ( .A(n_593), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x6_ASAP7_75t_L g652 ( .A(n_594), .B(n_653), .Y(n_652) );
OR2x6_ASAP7_75t_L g683 ( .A(n_594), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g669 ( .A(n_597), .Y(n_669) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g611 ( .A(n_600), .Y(n_611) );
INVx2_ASAP7_75t_L g619 ( .A(n_600), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_600), .B(n_609), .Y(n_629) );
INVx1_ASAP7_75t_L g640 ( .A(n_600), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_600), .B(n_601), .Y(n_645) );
INVx1_ASAP7_75t_L g680 ( .A(n_600), .Y(n_680) );
INVx2_ASAP7_75t_L g609 ( .A(n_601), .Y(n_609) );
AND2x4_ASAP7_75t_L g618 ( .A(n_601), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g641 ( .A(n_601), .Y(n_641) );
INVx1_ASAP7_75t_L g659 ( .A(n_601), .Y(n_659) );
OAI31xp33_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_620), .A3(n_654), .B(n_685), .Y(n_602) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx2_ASAP7_75t_L g615 ( .A(n_606), .Y(n_615) );
AND2x4_ASAP7_75t_L g622 ( .A(n_606), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g674 ( .A(n_607), .Y(n_674) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g684 ( .A(n_609), .Y(n_684) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AND2x4_ASAP7_75t_L g656 ( .A(n_614), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g666 ( .A(n_617), .Y(n_666) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g635 ( .A(n_618), .Y(n_635) );
AND2x4_ASAP7_75t_L g658 ( .A(n_619), .B(n_659), .Y(n_658) );
CKINVDCx6p67_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_630), .B1(n_631), .B2(n_636), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g661 ( .A(n_626), .Y(n_661) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g653 ( .A(n_639), .Y(n_653) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx8_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_658), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_667), .C(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_681), .B2(n_682), .Y(n_676) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
CKINVDCx11_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_694), .Y(n_686) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
OR2x6_ASAP7_75t_L g692 ( .A(n_690), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g695 ( .A(n_690), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g697 ( .A(n_690), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
CKINVDCx20_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OR2x6_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .Y(n_702) );
OR2x4_ASAP7_75t_L g727 ( .A(n_703), .B(n_707), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_704), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g734 ( .A(n_704), .Y(n_734) );
INVx1_ASAP7_75t_L g723 ( .A(n_705), .Y(n_723) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI31xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .A3(n_712), .B(n_714), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx6_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B1(n_731), .B2(n_732), .Y(n_724) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx8_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_729), .Y(n_730) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
endmodule