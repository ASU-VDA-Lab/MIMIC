module fake_jpeg_20840_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_13),
.B(n_10),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_25),
.B1(n_16),
.B2(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_35),
.B1(n_24),
.B2(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_12),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_48),
.B(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_28),
.B1(n_29),
.B2(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_42),
.B1(n_47),
.B2(n_39),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_30),
.B(n_34),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_29),
.A3(n_28),
.B1(n_15),
.B2(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_38),
.B1(n_40),
.B2(n_14),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_18),
.B(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_46),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_69),
.B1(n_48),
.B2(n_11),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_58),
.C(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_49),
.B1(n_56),
.B2(n_38),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_68),
.B1(n_67),
.B2(n_19),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.C(n_22),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_10),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_82),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_83),
.B1(n_81),
.B2(n_70),
.Y(n_87)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_83),
.A3(n_22),
.B1(n_9),
.B2(n_8),
.C1(n_6),
.C2(n_1),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_85),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_2),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_4),
.B(n_5),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_4),
.Y(n_93)
);


endmodule