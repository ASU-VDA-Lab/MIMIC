module real_aes_8553_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_1), .A2(n_144), .B(n_148), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g197 ( .A(n_2), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_3), .A2(n_139), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_4), .B(n_161), .Y(n_478) );
AOI21xp33_ASAP7_75t_L g165 ( .A1(n_5), .A2(n_139), .B(n_166), .Y(n_165) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_7), .A2(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_8), .B(n_41), .Y(n_115) );
INVx1_ASAP7_75t_L g534 ( .A(n_9), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_10), .B(n_170), .Y(n_513) );
INVx1_ASAP7_75t_L g172 ( .A(n_11), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_12), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g137 ( .A(n_13), .Y(n_137) );
INVx1_ASAP7_75t_L g253 ( .A(n_14), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_15), .A2(n_156), .B(n_254), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_16), .B(n_161), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_17), .B(n_153), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_18), .B(n_139), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_19), .B(n_562), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_20), .A2(n_180), .B(n_239), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_21), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_22), .B(n_170), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_23), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_24), .B(n_170), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_25), .Y(n_458) );
INVx1_ASAP7_75t_L g484 ( .A(n_26), .Y(n_484) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_27), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_28), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_29), .B(n_170), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_30), .A2(n_105), .B1(n_116), .B2(n_760), .Y(n_104) );
INVx1_ASAP7_75t_L g559 ( .A(n_31), .Y(n_559) );
INVx1_ASAP7_75t_L g186 ( .A(n_32), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_33), .A2(n_92), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_33), .Y(n_749) );
INVx2_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_35), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_36), .A2(n_157), .B(n_239), .C(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g560 ( .A(n_37), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_38), .A2(n_144), .B(n_148), .C(n_211), .Y(n_210) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_39), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_40), .A2(n_148), .B(n_483), .C(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g184 ( .A(n_42), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_43), .A2(n_50), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_43), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_44), .A2(n_64), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_44), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_45), .A2(n_729), .B1(n_730), .B2(n_733), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_45), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_46), .A2(n_169), .B(n_215), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_47), .B(n_170), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_48), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_49), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_50), .Y(n_744) );
INVx1_ASAP7_75t_L g499 ( .A(n_51), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_52), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_53), .B(n_139), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_54), .A2(n_148), .B1(n_180), .B2(n_182), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_55), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_56), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_57), .A2(n_157), .B(n_169), .C(n_171), .Y(n_168) );
CKINVDCx14_ASAP7_75t_R g531 ( .A(n_58), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_59), .Y(n_229) );
INVx1_ASAP7_75t_L g167 ( .A(n_60), .Y(n_167) );
INVx1_ASAP7_75t_L g145 ( .A(n_61), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_62), .Y(n_735) );
INVx1_ASAP7_75t_L g136 ( .A(n_63), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_64), .Y(n_731) );
INVx1_ASAP7_75t_SL g477 ( .A(n_65), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_66), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_67), .B(n_161), .Y(n_503) );
INVx1_ASAP7_75t_L g461 ( .A(n_68), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_69), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_SL g152 ( .A1(n_70), .A2(n_153), .B(n_154), .C(n_157), .Y(n_152) );
INVxp67_ASAP7_75t_L g155 ( .A(n_71), .Y(n_155) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_73), .A2(n_139), .B(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_74), .A2(n_727), .B1(n_728), .B2(n_734), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_74), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_75), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_76), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_77), .A2(n_139), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g222 ( .A(n_78), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_79), .A2(n_247), .B(n_555), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_80), .Y(n_481) );
INVx1_ASAP7_75t_L g519 ( .A(n_81), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_82), .A2(n_144), .B(n_148), .C(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_83), .A2(n_139), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g522 ( .A(n_84), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_85), .B(n_198), .Y(n_212) );
INVx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g512 ( .A(n_87), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_88), .B(n_153), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_89), .A2(n_144), .B(n_148), .C(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g755 ( .A(n_90), .B(n_112), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_91), .A2(n_148), .B(n_460), .C(n_464), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_92), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_92), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_93), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_94), .A2(n_144), .B(n_148), .C(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_95), .Y(n_243) );
INVx1_ASAP7_75t_L g151 ( .A(n_96), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_97), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_98), .B(n_198), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_99), .B(n_132), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_100), .B(n_132), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_101), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_102), .A2(n_139), .B(n_146), .Y(n_138) );
INVx2_ASAP7_75t_L g502 ( .A(n_103), .Y(n_502) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g760 ( .A(n_106), .Y(n_760) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_109), .A2(n_113), .B1(n_118), .B2(n_735), .Y(n_117) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g121 ( .A(n_111), .Y(n_121) );
INVx2_ASAP7_75t_L g448 ( .A(n_111), .Y(n_448) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AO221x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_736), .B1(n_741), .B2(n_751), .C(n_756), .Y(n_116) );
XOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_726), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_122), .B1(n_448), .B2(n_449), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND4x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_366), .C(n_413), .D(n_433), .Y(n_124) );
NOR3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_296), .C(n_321), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_204), .B(n_256), .C(n_286), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_175), .Y(n_128) );
INVx3_ASAP7_75t_SL g338 ( .A(n_129), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_129), .B(n_269), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_129), .B(n_191), .Y(n_419) );
AND2x2_ASAP7_75t_L g442 ( .A(n_129), .B(n_308), .Y(n_442) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_163), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g260 ( .A(n_131), .B(n_164), .Y(n_260) );
INVx3_ASAP7_75t_L g273 ( .A(n_131), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_131), .B(n_163), .Y(n_278) );
OR2x2_ASAP7_75t_L g329 ( .A(n_131), .B(n_270), .Y(n_329) );
BUFx2_ASAP7_75t_L g349 ( .A(n_131), .Y(n_349) );
AND2x2_ASAP7_75t_L g359 ( .A(n_131), .B(n_270), .Y(n_359) );
AND2x2_ASAP7_75t_L g365 ( .A(n_131), .B(n_176), .Y(n_365) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_138), .B(n_160), .Y(n_131) );
INVx4_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_132), .Y(n_471) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_134), .B(n_135), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx2_ASAP7_75t_L g247 ( .A(n_139), .Y(n_247) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_140), .B(n_144), .Y(n_188) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g487 ( .A(n_141), .Y(n_487) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
INVx1_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx1_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
INVx1_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
INVx4_ASAP7_75t_SL g159 ( .A(n_144), .Y(n_159) );
BUFx3_ASAP7_75t_L g488 ( .A(n_144), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_151), .B(n_152), .C(n_159), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_147), .A2(n_159), .B(n_167), .C(n_168), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_147), .A2(n_159), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_147), .A2(n_159), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_147), .A2(n_159), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_147), .A2(n_159), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_147), .A2(n_159), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_147), .A2(n_159), .B(n_556), .C(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx3_ASAP7_75t_L g216 ( .A(n_149), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_156), .B(n_172), .Y(n_171) );
INVx5_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_156), .B(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_158), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_159), .A2(n_179), .B1(n_187), .B2(n_188), .Y(n_178) );
INVx1_ASAP7_75t_L g464 ( .A(n_159), .Y(n_464) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_161), .A2(n_165), .B(n_173), .Y(n_164) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_162), .B(n_219), .Y(n_218) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_162), .A2(n_457), .B(n_465), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_162), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_162), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_164), .B(n_270), .Y(n_284) );
INVx2_ASAP7_75t_L g294 ( .A(n_164), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_164), .B(n_273), .Y(n_307) );
OR2x2_ASAP7_75t_L g318 ( .A(n_164), .B(n_270), .Y(n_318) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_164), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g376 ( .A(n_164), .Y(n_376) );
AND2x2_ASAP7_75t_L g422 ( .A(n_164), .B(n_176), .Y(n_422) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g239 ( .A(n_170), .Y(n_239) );
INVx1_ASAP7_75t_L g203 ( .A(n_174), .Y(n_203) );
INVx2_ASAP7_75t_L g233 ( .A(n_174), .Y(n_233) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_174), .A2(n_246), .B(n_255), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_174), .A2(n_188), .B(n_481), .C(n_482), .Y(n_480) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_174), .A2(n_529), .B(n_535), .Y(n_528) );
INVx3_ASAP7_75t_SL g295 ( .A(n_175), .Y(n_295) );
OR2x2_ASAP7_75t_L g348 ( .A(n_175), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
INVx3_ASAP7_75t_L g270 ( .A(n_176), .Y(n_270) );
AND2x2_ASAP7_75t_L g337 ( .A(n_176), .B(n_192), .Y(n_337) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_176), .Y(n_405) );
AOI33xp33_ASAP7_75t_L g409 ( .A1(n_176), .A2(n_338), .A3(n_345), .B1(n_354), .B2(n_410), .B3(n_411), .Y(n_409) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_189), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_177), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_177), .A2(n_193), .B(n_201), .Y(n_192) );
INVx2_ASAP7_75t_L g217 ( .A(n_177), .Y(n_217) );
INVx2_ASAP7_75t_L g200 ( .A(n_180), .Y(n_200) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_182) );
INVx2_ASAP7_75t_L g185 ( .A(n_183), .Y(n_185) );
INVx4_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
INVx2_ASAP7_75t_L g462 ( .A(n_185), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_188), .A2(n_222), .B(n_223), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_188), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_188), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_191), .B(n_273), .Y(n_272) );
NOR3xp33_ASAP7_75t_L g332 ( .A(n_191), .B(n_333), .C(n_335), .Y(n_332) );
AND2x2_ASAP7_75t_L g358 ( .A(n_191), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_191), .B(n_365), .Y(n_368) );
AND2x2_ASAP7_75t_L g421 ( .A(n_191), .B(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g277 ( .A(n_192), .Y(n_277) );
OR2x2_ASAP7_75t_L g371 ( .A(n_192), .B(n_270), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .C(n_200), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_198), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_198), .A2(n_251), .B1(n_559), .B2(n_560), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_203), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_203), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_203), .A2(n_508), .B(n_514), .Y(n_507) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_230), .Y(n_204) );
AOI32xp33_ASAP7_75t_L g322 ( .A1(n_205), .A2(n_323), .A3(n_325), .B1(n_327), .B2(n_330), .Y(n_322) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_205), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g425 ( .A(n_205), .Y(n_425) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g357 ( .A(n_206), .B(n_341), .Y(n_357) );
AND2x2_ASAP7_75t_L g377 ( .A(n_206), .B(n_303), .Y(n_377) );
AND2x2_ASAP7_75t_L g445 ( .A(n_206), .B(n_363), .Y(n_445) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_220), .Y(n_206) );
INVx3_ASAP7_75t_L g266 ( .A(n_207), .Y(n_266) );
AND2x2_ASAP7_75t_L g280 ( .A(n_207), .B(n_264), .Y(n_280) );
OR2x2_ASAP7_75t_L g285 ( .A(n_207), .B(n_263), .Y(n_285) );
INVx1_ASAP7_75t_L g292 ( .A(n_207), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_207), .B(n_274), .Y(n_300) );
AND2x2_ASAP7_75t_L g302 ( .A(n_207), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_207), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g355 ( .A(n_207), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_207), .B(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_210), .B(n_217), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_214), .A2(n_225), .B(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_214), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_214), .A2(n_462), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
INVx1_ASAP7_75t_L g227 ( .A(n_217), .Y(n_227) );
INVx2_ASAP7_75t_L g264 ( .A(n_220), .Y(n_264) );
AND2x2_ASAP7_75t_L g310 ( .A(n_220), .B(n_231), .Y(n_310) );
AND2x2_ASAP7_75t_L g320 ( .A(n_220), .B(n_245), .Y(n_320) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_227), .B(n_228), .Y(n_220) );
INVx1_ASAP7_75t_L g553 ( .A(n_227), .Y(n_553) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_227), .A2(n_570), .B(n_571), .Y(n_569) );
INVx2_ASAP7_75t_L g440 ( .A(n_230), .Y(n_440) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_244), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_231), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
AND2x2_ASAP7_75t_L g325 ( .A(n_231), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g341 ( .A(n_231), .B(n_304), .Y(n_341) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g289 ( .A(n_232), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_232), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g354 ( .A(n_232), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_232), .B(n_264), .Y(n_386) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_242), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_233), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g562 ( .A(n_233), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_239), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g265 ( .A(n_244), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_244), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g363 ( .A(n_244), .Y(n_363) );
INVx1_ASAP7_75t_L g396 ( .A(n_244), .Y(n_396) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g274 ( .A(n_245), .B(n_264), .Y(n_274) );
INVx1_ASAP7_75t_L g304 ( .A(n_245), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_251), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_251), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_251), .B(n_522), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_261), .B1(n_267), .B2(n_274), .C(n_275), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_258), .B(n_278), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_258), .B(n_341), .Y(n_418) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_260), .B(n_308), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_260), .B(n_269), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_260), .B(n_283), .Y(n_412) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g334 ( .A(n_264), .Y(n_334) );
AND2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g387 ( .A(n_265), .Y(n_387) );
AND2x2_ASAP7_75t_L g319 ( .A(n_266), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_266), .B(n_289), .Y(n_335) );
AND2x2_ASAP7_75t_L g399 ( .A(n_266), .B(n_325), .Y(n_399) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g308 ( .A(n_270), .B(n_277), .Y(n_308) );
AND2x2_ASAP7_75t_L g404 ( .A(n_271), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_273), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_274), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_274), .B(n_281), .Y(n_369) );
AND2x2_ASAP7_75t_L g389 ( .A(n_274), .B(n_289), .Y(n_389) );
AND2x2_ASAP7_75t_L g410 ( .A(n_274), .B(n_354), .Y(n_410) );
OAI32xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .A3(n_281), .B1(n_282), .B2(n_285), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_SL g283 ( .A(n_277), .Y(n_283) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_277), .B(n_307), .Y(n_324) );
OR2x2_ASAP7_75t_L g328 ( .A(n_277), .B(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_277), .B(n_376), .Y(n_429) );
INVx1_ASAP7_75t_L g297 ( .A(n_278), .Y(n_297) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_279), .A2(n_370), .B1(n_416), .B2(n_419), .C(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g287 ( .A(n_280), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g330 ( .A(n_280), .B(n_303), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_280), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g408 ( .A(n_280), .B(n_341), .Y(n_408) );
INVxp67_ASAP7_75t_L g344 ( .A(n_281), .Y(n_344) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_L g414 ( .A(n_283), .B(n_401), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_283), .B(n_364), .Y(n_437) );
INVx1_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_285), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g430 ( .A(n_285), .B(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_290), .B(n_293), .Y(n_286) );
AND2x2_ASAP7_75t_L g299 ( .A(n_288), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g383 ( .A(n_292), .B(n_303), .Y(n_383) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g401 ( .A(n_294), .B(n_359), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_294), .B(n_358), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_295), .B(n_307), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_301), .C(n_311), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_332), .B1(n_336), .B2(n_339), .C(n_342), .Y(n_331) );
AOI31xp33_ASAP7_75t_L g426 ( .A1(n_297), .A2(n_427), .A3(n_428), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_307), .B2(n_309), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g427 ( .A(n_307), .Y(n_427) );
INVx1_ASAP7_75t_L g390 ( .A(n_308), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_310), .A2(n_434), .B(n_436), .C(n_438), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_315), .B2(n_319), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_318), .A2(n_352), .B1(n_371), .B2(n_407), .C(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g402 ( .A(n_319), .Y(n_402) );
INVx1_ASAP7_75t_L g356 ( .A(n_320), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g321 ( .A(n_322), .B(n_331), .C(n_346), .Y(n_321) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_323), .A2(n_373), .B(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_325), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g432 ( .A(n_326), .Y(n_432) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g370 ( .A(n_333), .B(n_353), .Y(n_370) );
INVx1_ASAP7_75t_L g345 ( .A(n_334), .Y(n_345) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g343 ( .A(n_337), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_337), .B(n_375), .Y(n_374) );
NOR4xp25_ASAP7_75t_L g342 ( .A(n_338), .B(n_343), .C(n_344), .D(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_351), .B1(n_357), .B2(n_358), .C1(n_360), .C2(n_364), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g444 ( .A(n_348), .Y(n_444) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_360), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_SL g420 ( .A1(n_365), .A2(n_421), .B(n_423), .Y(n_420) );
NOR4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_378), .C(n_391), .D(n_406), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_369), .B1(n_370), .B2(n_371), .C(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g447 ( .A(n_368), .Y(n_447) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_375), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OAI222xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_382), .B1(n_384), .B2(n_385), .C1(n_388), .C2(n_390), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_383), .A2(n_414), .B(n_415), .C(n_426), .Y(n_413) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
OAI222xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .B1(n_398), .B2(n_400), .C1(n_402), .C2(n_403), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_408), .A2(n_411), .B1(n_444), .B2(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_441), .B(n_443), .C(n_446), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_449), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_681), .Y(n_449) );
NOR4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_618), .C(n_652), .D(n_668), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_548), .C(n_582), .D(n_598), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_491), .B1(n_524), .B2(n_536), .C1(n_541), .C2(n_547), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI31xp33_ASAP7_75t_L g714 ( .A1(n_454), .A2(n_715), .A3(n_716), .B(n_718), .Y(n_714) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_467), .Y(n_454) );
AND2x2_ASAP7_75t_L g689 ( .A(n_455), .B(n_469), .Y(n_689) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g540 ( .A(n_456), .Y(n_540) );
AND2x2_ASAP7_75t_L g547 ( .A(n_456), .B(n_479), .Y(n_547) );
AND2x2_ASAP7_75t_L g603 ( .A(n_456), .B(n_470), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_467), .B(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_468), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_468), .B(n_551), .Y(n_593) );
AND2x2_ASAP7_75t_L g686 ( .A(n_468), .B(n_626), .Y(n_686) );
OAI321xp33_ASAP7_75t_L g720 ( .A1(n_468), .A2(n_540), .A3(n_693), .B1(n_721), .B2(n_723), .C(n_724), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_468), .B(n_527), .C(n_633), .D(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AND2x2_ASAP7_75t_L g588 ( .A(n_469), .B(n_538), .Y(n_588) );
AND2x2_ASAP7_75t_L g607 ( .A(n_469), .B(n_540), .Y(n_607) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g539 ( .A(n_470), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g563 ( .A(n_470), .B(n_479), .Y(n_563) );
AND2x2_ASAP7_75t_L g649 ( .A(n_470), .B(n_538), .Y(n_649) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_478), .Y(n_470) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_471), .A2(n_497), .B(n_503), .Y(n_496) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_471), .A2(n_517), .B(n_523), .Y(n_516) );
INVx3_ASAP7_75t_SL g538 ( .A(n_479), .Y(n_538) );
AND2x2_ASAP7_75t_L g581 ( .A(n_479), .B(n_568), .Y(n_581) );
OR2x2_ASAP7_75t_L g614 ( .A(n_479), .B(n_540), .Y(n_614) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_479), .Y(n_621) );
AND2x2_ASAP7_75t_L g650 ( .A(n_479), .B(n_539), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_479), .B(n_623), .Y(n_665) );
AND2x2_ASAP7_75t_L g697 ( .A(n_479), .B(n_689), .Y(n_697) );
AND2x2_ASAP7_75t_L g706 ( .A(n_479), .B(n_552), .Y(n_706) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_487), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
INVx1_ASAP7_75t_SL g674 ( .A(n_493), .Y(n_674) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g543 ( .A(n_494), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g526 ( .A(n_495), .B(n_506), .Y(n_526) );
AND2x2_ASAP7_75t_L g610 ( .A(n_495), .B(n_528), .Y(n_610) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g580 ( .A(n_496), .B(n_516), .Y(n_580) );
OR2x2_ASAP7_75t_L g591 ( .A(n_496), .B(n_528), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_496), .B(n_528), .Y(n_617) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_496), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_504), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_504), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g590 ( .A(n_505), .B(n_591), .Y(n_590) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_505), .A2(n_580), .A3(n_586), .B1(n_617), .B2(n_667), .C1(n_677), .C2(n_679), .Y(n_676) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_516), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_506), .B(n_527), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_506), .B(n_528), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_506), .B(n_544), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_506), .B(n_617), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_506), .Y(n_655) );
AND2x2_ASAP7_75t_L g667 ( .A(n_506), .B(n_516), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_506), .B(n_543), .Y(n_699) );
INVx4_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g564 ( .A(n_507), .B(n_516), .Y(n_564) );
BUFx3_ASAP7_75t_L g578 ( .A(n_507), .Y(n_578) );
AND3x2_ASAP7_75t_L g660 ( .A(n_507), .B(n_640), .C(n_661), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_516), .B(n_526), .C(n_527), .Y(n_525) );
INVx1_ASAP7_75t_SL g544 ( .A(n_516), .Y(n_544) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_516), .Y(n_645) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g639 ( .A(n_526), .B(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g646 ( .A(n_526), .Y(n_646) );
AND2x2_ASAP7_75t_L g684 ( .A(n_527), .B(n_662), .Y(n_684) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g565 ( .A(n_528), .Y(n_565) );
AND2x2_ASAP7_75t_L g640 ( .A(n_528), .B(n_544), .Y(n_640) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OR2x2_ASAP7_75t_L g584 ( .A(n_538), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g703 ( .A(n_538), .B(n_603), .Y(n_703) );
AND2x2_ASAP7_75t_L g717 ( .A(n_538), .B(n_540), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_539), .B(n_552), .Y(n_658) );
AND2x2_ASAP7_75t_L g705 ( .A(n_539), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g568 ( .A(n_540), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g585 ( .A(n_540), .B(n_552), .Y(n_585) );
INVx1_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
AND2x2_ASAP7_75t_L g626 ( .A(n_540), .B(n_552), .Y(n_626) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_542), .A2(n_669), .B1(n_673), .B2(n_675), .C(n_676), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g572 ( .A(n_543), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_546), .B(n_579), .Y(n_722) );
AOI322xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_564), .A3(n_565), .B1(n_566), .B2(n_572), .C1(n_574), .C2(n_581), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_563), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_551), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_551), .B(n_613), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_551), .A2(n_563), .B(n_637), .C(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_551), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_551), .B(n_607), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_551), .B(n_689), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_551), .B(n_717), .Y(n_716) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_552), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_552), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g678 ( .A(n_552), .B(n_565), .Y(n_678) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B(n_561), .Y(n_552) );
INVx1_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_561), .Y(n_571) );
INVx1_ASAP7_75t_L g653 ( .A(n_563), .Y(n_653) );
OAI31xp33_ASAP7_75t_L g663 ( .A1(n_563), .A2(n_588), .A3(n_664), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_563), .B(n_569), .Y(n_715) );
INVx1_ASAP7_75t_SL g576 ( .A(n_564), .Y(n_576) );
AND2x2_ASAP7_75t_L g609 ( .A(n_564), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g690 ( .A(n_564), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g600 ( .A(n_565), .Y(n_600) );
AND2x2_ASAP7_75t_L g627 ( .A(n_565), .B(n_580), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_565), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g719 ( .A(n_565), .B(n_667), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_567), .B(n_637), .Y(n_710) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g624 ( .A(n_569), .Y(n_624) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_575), .B(n_577), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_576), .A2(n_619), .B(n_625), .C(n_641), .Y(n_618) );
OR2x2_ASAP7_75t_L g693 ( .A(n_576), .B(n_674), .Y(n_693) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_578), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_578), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B(n_589), .C(n_592), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g633 ( .A(n_585), .Y(n_633) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_588), .B(n_626), .Y(n_631) );
INVx1_ASAP7_75t_L g637 ( .A(n_588), .Y(n_637) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g596 ( .A(n_591), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g629 ( .A(n_591), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g691 ( .A(n_591), .Y(n_691) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B(n_596), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_605), .B(n_608), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_604), .C(n_611), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_599), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_602), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g615 ( .A(n_603), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_605), .A2(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_610), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g635 ( .A(n_610), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_615), .B(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g666 ( .A(n_617), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_623), .B(n_649), .Y(n_675) );
AND2x2_ASAP7_75t_L g688 ( .A(n_623), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g702 ( .A(n_623), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g712 ( .A(n_623), .B(n_650), .Y(n_712) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_628), .C(n_636), .Y(n_625) );
INVx1_ASAP7_75t_L g672 ( .A(n_626), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_632), .B2(n_634), .Y(n_628) );
OR2x2_ASAP7_75t_L g634 ( .A(n_630), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_630), .B(n_691), .Y(n_713) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g707 ( .A(n_640), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_647), .B1(n_650), .B2(n_651), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g725 ( .A(n_645), .Y(n_725) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g671 ( .A(n_649), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_663), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_671), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR5xp2_ASAP7_75t_L g681 ( .A(n_682), .B(n_700), .C(n_708), .D(n_714), .E(n_720), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_687), .C(n_694), .Y(n_682) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_692), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_697), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_707), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g723 ( .A(n_703), .Y(n_723) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g752 ( .A(n_740), .Y(n_752) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_741) );
INVx1_ASAP7_75t_L g750 ( .A(n_742), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g759 ( .A(n_755), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule