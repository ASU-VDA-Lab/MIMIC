module real_jpeg_4523_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_279;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_1),
.A2(n_23),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_1),
.A2(n_23),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_164),
.B1(n_165),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_5),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_5),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_8),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_95),
.B(n_98),
.C(n_104),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_81),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_134),
.C(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_8),
.B(n_26),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_120),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_8),
.A2(n_65),
.B1(n_81),
.B2(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_56),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_11),
.A2(n_56),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_11),
.A2(n_56),
.B1(n_79),
.B2(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_203),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_201),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_139),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_15),
.B(n_139),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_93),
.C(n_108),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_16),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_58),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_17),
.B(n_59),
.C(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_22),
.Y(n_148)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_25),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_26),
.B(n_52),
.Y(n_196)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_38),
.Y(n_211)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_42),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_43),
.B(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_61),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_61),
.B(n_188),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_83),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_71),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_77),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_72),
.B(n_87),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_72),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_73),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_74),
.Y(n_226)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_91),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_81),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_81),
.A2(n_153),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_83),
.B(n_221),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_93),
.A2(n_108),
.B1(n_109),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_93),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_94),
.A2(n_105),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_94),
.Y(n_275)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_103),
.Y(n_233)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_123),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_112),
.A2(n_119),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_113),
.B(n_129),
.Y(n_215)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_120),
.B(n_124),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_120),
.B(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_123),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_129),
.B(n_230),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_137),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_174),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_162),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.A3(n_150),
.B1(n_152),
.B2(n_157),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_170),
.B(n_173),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_191),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_187),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_277),
.B(n_282),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_261),
.B(n_276),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_237),
.B(n_260),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_244),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_235),
.C(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_247),
.B(n_259),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_258),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_264),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_268),
.C(n_273),
.Y(n_281)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_281),
.Y(n_282)
);


endmodule