module fake_jpeg_13548_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_62),
.Y(n_69)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_1),
.B(n_4),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_50),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_49),
.B1(n_50),
.B2(n_48),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_78),
.B1(n_62),
.B2(n_61),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_39),
.B1(n_51),
.B2(n_43),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_75),
.B(n_5),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_55),
.B1(n_54),
.B2(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_7),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_46),
.B1(n_44),
.B2(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_44),
.B(n_6),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_92),
.C(n_18),
.Y(n_104)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_5),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_89),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_15),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_9),
.B(n_10),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.C(n_103),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_16),
.B(n_17),
.Y(n_96)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22x1_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_37),
.B1(n_20),
.B2(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_35),
.C(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_22),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_99),
.C(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_114),
.B1(n_96),
.B2(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_24),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_100),
.B1(n_115),
.B2(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_25),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_114),
.B1(n_113),
.B2(n_117),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_98),
.A3(n_118),
.B1(n_116),
.B2(n_121),
.C1(n_108),
.C2(n_112),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_30),
.C(n_31),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_32),
.Y(n_127)
);


endmodule