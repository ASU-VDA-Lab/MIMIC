module real_jpeg_26640_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_273, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_273;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_4),
.B1(n_25),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_3),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_20),
.B(n_22),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_29),
.B1(n_58),
.B2(n_59),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_29),
.B1(n_38),
.B2(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_19),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_5),
.B(n_38),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_55),
.B(n_59),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_37),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_4),
.A2(n_9),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_4),
.A2(n_8),
.B1(n_25),
.B2(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_4),
.A2(n_21),
.B(n_29),
.C(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_20),
.B1(n_23),
.B2(n_39),
.Y(n_42)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_20),
.B1(n_23),
.B2(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_38),
.B1(n_40),
.B2(n_47),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_9),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_9),
.A2(n_26),
.B1(n_38),
.B2(n_40),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_20),
.B1(n_23),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_10),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_207)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_11),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_77),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_76),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_16),
.B(n_62),
.Y(n_76)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_16),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_32),
.CI(n_43),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B(n_27),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_18),
.A2(n_27),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_19),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_19),
.B(n_30),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_20),
.A2(n_29),
.B(n_145),
.C(n_146),
.Y(n_144)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_28),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_29),
.A2(n_38),
.B(n_56),
.C(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_29),
.B(n_101),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_29),
.B(n_57),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_37),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_36),
.B(n_88),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_49),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_40),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.C(n_50),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_65),
.B1(n_85),
.B2(n_90),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_44),
.B(n_90),
.C(n_91),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_44),
.A2(n_65),
.B1(n_105),
.B2(n_128),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_44),
.B(n_128),
.C(n_223),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_50),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_50),
.A2(n_69),
.B1(n_72),
.B2(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_53),
.A2(n_57),
.B1(n_109),
.B2(n_115),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_57),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_58),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_98),
.Y(n_97)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_70),
.C(n_71),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_129),
.Y(n_263)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_105),
.C(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_70),
.A2(n_129),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_70),
.A2(n_129),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_71),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_72),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_87),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_254),
.A3(n_264),
.B1(n_269),
.B2(n_270),
.C(n_273),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_236),
.B(n_253),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_217),
.B(n_235),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_138),
.B(n_200),
.C(n_216),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_125),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_82),
.B(n_125),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_102),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_83),
.B(n_103),
.C(n_111),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_135),
.C(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_85),
.A2(n_90),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_85),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_85),
.B(n_242),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_95),
.A2(n_133),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_95),
.B(n_183),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_95),
.B(n_160),
.C(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_98),
.B(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_97),
.B(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_97),
.A2(n_101),
.B1(n_120),
.B2(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_110),
.B2(n_111),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_105),
.A2(n_112),
.B1(n_113),
.B2(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_112),
.A2(n_113),
.B1(n_167),
.B2(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_119),
.Y(n_210)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_128),
.C(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_113),
.B(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_134),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_126),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_129),
.B(n_210),
.C(n_212),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_134),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_135),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_199),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_193),
.B(n_198),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_163),
.B(n_192),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_151),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_151),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_150),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_160),
.C(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_162),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_162),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_206),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_187),
.B(n_191),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_174),
.B(n_186),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B(n_185),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.B(n_184),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_201),
.B(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_214),
.B2(n_215),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_209),
.C(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_234),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_226),
.C(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_231),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_231),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_245),
.B(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_237),
.B(n_238),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_251),
.B2(n_252),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_244),
.C(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_256),
.C(n_260),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_256),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_261),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);


endmodule