module real_jpeg_3516_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_1),
.B(n_64),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_1),
.B(n_30),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_34),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_3),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_30),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_3),
.B(n_53),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_3),
.B(n_28),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_48),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_4),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_53),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_5),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_5),
.B(n_53),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_5),
.B(n_55),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_64),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_8),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_8),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_8),
.B(n_38),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_8),
.B(n_53),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_30),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_8),
.B(n_28),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_8),
.B(n_48),
.Y(n_228)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_64),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_55),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_14),
.B(n_28),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_14),
.B(n_64),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_14),
.B(n_34),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_249),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_246),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_209),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_131),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_95),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_22),
.B(n_95),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.C(n_84),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_23),
.B(n_206),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_23),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_40),
.CI(n_44),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_40),
.C(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.C(n_37),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_25),
.A2(n_26),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_26),
.A2(n_77),
.B(n_149),
.C(n_228),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_27),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_27),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_27),
.A2(n_29),
.B1(n_77),
.B2(n_149),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_27),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_29),
.A2(n_74),
.B1(n_77),
.B2(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_31),
.B(n_130),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_33),
.B(n_37),
.Y(n_202)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g222 ( 
.A(n_38),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_43),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_43),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_52),
.C(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_46),
.B(n_75),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_46),
.B(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_47),
.B(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_51),
.A2(n_52),
.B1(n_265),
.B2(n_268),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_55),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_59),
.B(n_84),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_71),
.B2(n_83),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_72),
.C(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_68),
.C(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_65),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_76),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.C(n_82),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_93),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_85),
.B(n_89),
.CI(n_93),
.CON(n_196),
.SN(n_196)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_92),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_142),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_95),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_117),
.CI(n_118),
.CON(n_95),
.SN(n_95)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_96),
.B(n_117),
.C(n_118),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_97),
.B(n_100),
.C(n_107),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_101),
.B(n_103),
.C(n_105),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_116),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_112),
.B(n_113),
.C(n_115),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_120),
.B(n_121),
.C(n_123),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_128),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_125),
.B(n_127),
.C(n_129),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_204),
.B(n_208),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_192),
.B(n_203),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_164),
.B(n_191),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_155),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_139),
.CI(n_140),
.CON(n_156),
.SN(n_156)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_151),
.C(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.C(n_163),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_188),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_156),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_185),
.B(n_190),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_176),
.B(n_184),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_172),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B(n_183),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_199),
.C(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_207),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_245),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_245),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_214),
.C(n_230),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_229),
.B2(n_230),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_225),
.CI(n_226),
.CON(n_215),
.SN(n_215)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_225),
.C(n_226),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_221),
.C(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_235),
.C(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_243),
.B2(n_244),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_241),
.C(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_284),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_283),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_283),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_269),
.B2(n_282),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_281),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);


endmodule