module fake_jpeg_22997_n_65 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_18),
.B1(n_27),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_45),
.C(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_44),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_32),
.B(n_1),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_11),
.B(n_14),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_6),
.C(n_9),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_20),
.C(n_21),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_59),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_54),
.B(n_56),
.Y(n_61)
);

OA21x2_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_22),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_58),
.Y(n_65)
);


endmodule