module real_jpeg_11752_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_344, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_344;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_45),
.B1(n_47),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_167),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_167),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_167),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_44),
.B1(n_64),
.B2(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_5),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_260)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_7),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_45),
.B1(n_47),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_34),
.C(n_50),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g163 ( 
.A(n_8),
.B(n_83),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_118),
.B(n_171),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_8),
.A2(n_64),
.B(n_82),
.C(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_8),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_59),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_12),
.A2(n_45),
.B1(n_47),
.B2(n_127),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_127),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_13),
.A2(n_45),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_13),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_55),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_13),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_14),
.A2(n_45),
.B1(n_47),
.B2(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_85),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_15),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_15),
.A2(n_45),
.B1(n_47),
.B2(n_61),
.Y(n_249)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_16),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_20),
.B(n_341),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_17),
.B(n_342),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_18),
.A2(n_59),
.B1(n_60),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_18),
.A2(n_45),
.B1(n_47),
.B2(n_74),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_74),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_18),
.A2(n_64),
.B1(n_65),
.B2(n_74),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_336),
.B(n_339),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_328),
.B(n_332),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_315),
.B(n_327),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_143),
.B(n_312),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_130),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_105),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_26),
.B(n_105),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_75),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_27),
.B(n_76),
.C(n_91),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_28),
.A2(n_29),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_30),
.A2(n_31),
.B1(n_57),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_37),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_32),
.A2(n_37),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_32),
.B(n_172),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_32),
.A2(n_37),
.B1(n_117),
.B2(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_33),
.B(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_37),
.B(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_39),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B1(n_53),
.B2(n_56),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_43),
.A2(n_48),
.B1(n_56),
.B2(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_47),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_45),
.B(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_47),
.A2(n_81),
.B(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_56),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_48),
.B(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_48),
.A2(n_56),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_48),
.A2(n_56),
.B1(n_122),
.B2(n_249),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_54),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_52),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_52),
.B(n_155),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_52),
.A2(n_168),
.B(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_56),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_68),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_62),
.B1(n_70),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_71)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_60),
.A2(n_70),
.B(n_155),
.C(n_242),
.Y(n_241)
);

AOI32xp33_ASAP7_75t_L g255 ( 
.A1(n_60),
.A2(n_64),
.A3(n_67),
.B1(n_243),
.B2(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_73),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_62),
.A2(n_70),
.B1(n_103),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_62),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_62),
.A2(n_68),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_62),
.A2(n_70),
.B1(n_126),
.B2(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g256 ( 
.A(n_63),
.B(n_65),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_65),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_69),
.A2(n_223),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_69),
.A2(n_223),
.B1(n_322),
.B2(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_69),
.A2(n_223),
.B(n_330),
.Y(n_338)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_91),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_77),
.B(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_78),
.A2(n_86),
.B1(n_96),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_78),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_78),
.A2(n_86),
.B1(n_218),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_78),
.A2(n_204),
.B(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_83),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_79),
.B(n_205),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_79),
.A2(n_83),
.B(n_319),
.Y(n_318)
);

NOR2x1_ASAP7_75t_R g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_83),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_86),
.A2(n_218),
.B(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_86),
.A2(n_124),
.B(n_219),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_89),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_89),
.A2(n_156),
.B(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_93),
.B(n_98),
.C(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_98),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_98),
.B(n_135),
.C(n_139),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_102),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_102),
.B(n_134),
.C(n_141),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_111),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_112),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.C(n_125),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_113),
.A2(n_114),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_115),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_118),
.A2(n_119),
.B1(n_200),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_118),
.A2(n_119),
.B1(n_226),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_119),
.A2(n_177),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_119),
.A2(n_185),
.B(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_123),
.B(n_125),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_129),
.B(n_241),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_130),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_142),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_131),
.B(n_142),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_136),
.Y(n_321)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_140),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_306),
.B(n_311),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_294),
.B(n_305),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_262),
.A3(n_287),
.B1(n_292),
.B2(n_293),
.C(n_344),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_235),
.B(n_261),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_212),
.B(n_234),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_193),
.B(n_211),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_173),
.B(n_192),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_151),
.B(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_169),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_181),
.B(n_191),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_179),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_186),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_206),
.C(n_210),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_227),
.B2(n_228),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_230),
.C(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_221),
.C(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_251),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_252),
.C(n_253),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_244),
.B2(n_250),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_245),
.C(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_277),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_273),
.C(n_276),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_265),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_286),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_281),
.C(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_284),
.C(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_304),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.C(n_300),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_323),
.C(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_337),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_338),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);


endmodule