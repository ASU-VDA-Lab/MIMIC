module real_aes_15701_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_0), .Y(n_1462) );
OAI211xp5_ASAP7_75t_L g550 ( .A1(n_1), .A2(n_551), .B(n_553), .C(n_568), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_1), .B(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_2), .A2(n_124), .B1(n_930), .B2(n_932), .Y(n_1210) );
AOI22xp33_ASAP7_75t_SL g1226 ( .A1(n_2), .A2(n_132), .B1(n_1030), .B2(n_1031), .Y(n_1226) );
INVx1_ASAP7_75t_L g924 ( .A(n_3), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_4), .A2(n_153), .B1(n_418), .B2(n_1011), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1040 ( .A(n_4), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_5), .A2(n_69), .B1(n_595), .B2(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_5), .A2(n_52), .B1(n_827), .B2(n_828), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_6), .A2(n_228), .B1(n_830), .B2(n_903), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_6), .A2(n_264), .B1(n_611), .B2(n_790), .Y(n_994) );
INVx1_ASAP7_75t_L g651 ( .A(n_7), .Y(n_651) );
AO22x1_ASAP7_75t_L g677 ( .A1(n_7), .A2(n_150), .B1(n_563), .B2(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g297 ( .A(n_8), .Y(n_297) );
AND2x2_ASAP7_75t_L g349 ( .A(n_8), .B(n_241), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_8), .B(n_307), .Y(n_368) );
AND2x2_ASAP7_75t_L g382 ( .A(n_8), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g661 ( .A(n_9), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_9), .A2(n_98), .B1(n_522), .B2(n_558), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g1209 ( .A1(n_10), .A2(n_163), .B1(n_625), .B2(n_1011), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_10), .A2(n_14), .B1(n_908), .B2(n_1222), .C(n_1223), .Y(n_1221) );
INVx1_ASAP7_75t_L g867 ( .A(n_11), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_11), .A2(n_161), .B1(n_888), .B2(n_889), .C(n_890), .Y(n_887) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_12), .B(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_12), .B(n_102), .Y(n_1254) );
INVx2_ASAP7_75t_L g1258 ( .A(n_12), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_13), .A2(n_89), .B1(n_586), .B2(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g1213 ( .A1(n_14), .A2(n_29), .B1(n_750), .B2(n_803), .Y(n_1213) );
INVx1_ASAP7_75t_L g1461 ( .A(n_15), .Y(n_1461) );
INVx1_ASAP7_75t_L g1207 ( .A(n_16), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g1214 ( .A1(n_17), .A2(n_220), .B1(n_763), .B2(n_881), .Y(n_1214) );
INVx1_ASAP7_75t_L g1229 ( .A(n_17), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_18), .A2(n_47), .B1(n_875), .B2(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_18), .A2(n_280), .B1(n_827), .B2(n_945), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_19), .A2(n_181), .B1(n_1253), .B2(n_1259), .Y(n_1295) );
INVx1_ASAP7_75t_L g1169 ( .A(n_20), .Y(n_1169) );
OAI22xp33_ASAP7_75t_L g1185 ( .A1(n_20), .A2(n_179), .B1(n_763), .B2(n_1186), .Y(n_1185) );
OAI221xp5_ASAP7_75t_L g1175 ( .A1(n_21), .A2(n_55), .B1(n_851), .B2(n_949), .C(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1197 ( .A(n_21), .Y(n_1197) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_22), .A2(n_570), .B(n_572), .C(n_574), .Y(n_569) );
INVx1_ASAP7_75t_L g630 ( .A(n_22), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_23), .A2(n_160), .B1(n_1512), .B2(n_1514), .Y(n_1511) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_23), .A2(n_240), .B1(n_905), .B2(n_1223), .C(n_1486), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1502 ( .A1(n_24), .A2(n_1503), .B1(n_1504), .B2(n_1534), .Y(n_1502) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_24), .Y(n_1503) );
INVx1_ASAP7_75t_L g922 ( .A(n_25), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_25), .A2(n_145), .B1(n_889), .B2(n_949), .C(n_950), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_26), .A2(n_206), .B1(n_1249), .B2(n_1256), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_27), .A2(n_172), .B1(n_750), .B2(n_930), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_27), .A2(n_148), .B1(n_903), .B2(n_1031), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_28), .A2(n_270), .B1(n_1108), .B2(n_1112), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1146 ( .A1(n_28), .A2(n_270), .B1(n_1147), .B2(n_1150), .Y(n_1146) );
A2O1A1Ixp33_ASAP7_75t_L g1230 ( .A1(n_29), .A2(n_850), .B(n_1231), .C(n_1237), .Y(n_1230) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_30), .A2(n_280), .B1(n_929), .B2(n_930), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_30), .A2(n_47), .B1(n_558), .B2(n_560), .C(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_31), .A2(n_85), .B1(n_416), .B2(n_750), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_31), .A2(n_168), .B1(n_823), .B2(n_905), .C(n_908), .Y(n_904) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_32), .B(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_32), .A2(n_164), .B1(n_416), .B2(n_759), .Y(n_758) );
XNOR2xp5_ASAP7_75t_L g962 ( .A(n_33), .B(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_34), .A2(n_164), .B1(n_555), .B2(n_678), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_34), .A2(n_256), .B1(n_416), .B2(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g1524 ( .A(n_35), .Y(n_1524) );
INVx1_ASAP7_75t_L g1466 ( .A(n_36), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_37), .A2(n_57), .B1(n_586), .B2(n_805), .Y(n_1217) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_37), .A2(n_1023), .B(n_1220), .C(n_1227), .Y(n_1219) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_38), .A2(n_111), .B1(n_1249), .B2(n_1256), .Y(n_1269) );
AOI22xp5_ASAP7_75t_L g1276 ( .A1(n_39), .A2(n_215), .B1(n_1249), .B2(n_1259), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_40), .A2(n_171), .B1(n_830), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_40), .A2(n_125), .B1(n_439), .B2(n_811), .Y(n_996) );
INVx1_ASAP7_75t_L g483 ( .A(n_41), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g1294 ( .A1(n_42), .A2(n_94), .B1(n_1249), .B2(n_1256), .Y(n_1294) );
XNOR2x2_ASAP7_75t_L g1201 ( .A(n_43), .B(n_1202), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_44), .A2(n_240), .B1(n_875), .B2(n_1512), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_44), .A2(n_160), .B1(n_1030), .B2(n_1031), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_45), .A2(n_63), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_45), .A2(n_275), .B1(n_418), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_46), .A2(n_137), .B1(n_800), .B2(n_801), .Y(n_799) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_46), .Y(n_848) );
INVx1_ASAP7_75t_L g406 ( .A(n_48), .Y(n_406) );
INVx1_ASAP7_75t_L g414 ( .A(n_48), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_49), .A2(n_131), .B1(n_416), .B2(n_418), .Y(n_1516) );
AOI221xp5_ASAP7_75t_L g1526 ( .A1(n_49), .A2(n_68), .B1(n_727), .B2(n_908), .C(n_1028), .Y(n_1526) );
INVx1_ASAP7_75t_L g709 ( .A(n_50), .Y(n_709) );
INVxp67_ASAP7_75t_SL g1160 ( .A(n_51), .Y(n_1160) );
AND4x1_ASAP7_75t_L g1200 ( .A(n_51), .B(n_1162), .C(n_1165), .D(n_1183), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_52), .A2(n_143), .B1(n_595), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_53), .A2(n_132), .B1(n_930), .B2(n_1069), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_53), .A2(n_124), .B1(n_1044), .B2(n_1233), .C(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g925 ( .A(n_54), .Y(n_925) );
INVx1_ASAP7_75t_L g1199 ( .A(n_55), .Y(n_1199) );
INVx1_ASAP7_75t_L g290 ( .A(n_56), .Y(n_290) );
INVx2_ASAP7_75t_L g426 ( .A(n_58), .Y(n_426) );
INVx1_ASAP7_75t_L g697 ( .A(n_59), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_60), .A2(n_80), .B1(n_1256), .B2(n_1264), .Y(n_1277) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_61), .Y(n_917) );
INVx1_ASAP7_75t_L g807 ( .A(n_62), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_63), .A2(n_97), .B1(n_418), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_64), .A2(n_65), .B1(n_418), .B2(n_803), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_64), .A2(n_153), .B1(n_825), .B2(n_1026), .C(n_1028), .Y(n_1025) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_65), .Y(n_1042) );
INVx1_ASAP7_75t_L g761 ( .A(n_66), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_67), .A2(n_193), .B1(n_796), .B2(n_873), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_67), .A2(n_138), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1510 ( .A1(n_68), .A2(n_239), .B1(n_418), .B2(n_803), .Y(n_1510) );
INVx1_ASAP7_75t_L g843 ( .A(n_69), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_70), .A2(n_130), .B1(n_1249), .B2(n_1256), .Y(n_1283) );
INVx1_ASAP7_75t_L g512 ( .A(n_71), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_71), .A2(n_133), .B1(n_521), .B2(n_524), .C(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_72), .A2(n_222), .B1(n_694), .B2(n_805), .Y(n_918) );
OAI211xp5_ASAP7_75t_L g937 ( .A1(n_72), .A2(n_900), .B(n_938), .C(n_946), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_73), .A2(n_268), .B1(n_763), .B2(n_881), .Y(n_1017) );
INVx1_ASAP7_75t_L g1035 ( .A(n_73), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_74), .A2(n_182), .B1(n_432), .B2(n_875), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_74), .A2(n_83), .B1(n_828), .B2(n_903), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_75), .A2(n_217), .B1(n_694), .B2(n_805), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1166 ( .A1(n_75), .A2(n_1023), .B(n_1167), .C(n_1170), .Y(n_1166) );
OAI222xp33_ASAP7_75t_L g667 ( .A1(n_76), .A2(n_214), .B1(n_455), .B2(n_459), .C1(n_668), .C2(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g681 ( .A(n_76), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_77), .Y(n_1064) );
INVx1_ASAP7_75t_L g782 ( .A(n_78), .Y(n_782) );
OAI222xp33_ASAP7_75t_L g834 ( .A1(n_78), .A2(n_127), .B1(n_835), .B2(n_838), .C1(n_844), .C2(n_851), .Y(n_834) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_79), .A2(n_100), .B1(n_720), .B2(n_721), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g735 ( .A1(n_79), .A2(n_614), .B(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g1468 ( .A1(n_81), .A2(n_88), .B1(n_428), .B2(n_932), .Y(n_1468) );
AOI221xp5_ASAP7_75t_L g1481 ( .A1(n_81), .A2(n_126), .B1(n_727), .B2(n_908), .C(n_1028), .Y(n_1481) );
INVx1_ASAP7_75t_L g1506 ( .A(n_82), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_83), .A2(n_107), .B1(n_873), .B2(n_875), .Y(n_872) );
INVx1_ASAP7_75t_L g968 ( .A(n_84), .Y(n_968) );
INVxp67_ASAP7_75t_SL g892 ( .A(n_85), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_86), .A2(n_129), .B1(n_1249), .B2(n_1256), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_87), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g1485 ( .A1(n_88), .A2(n_216), .B1(n_521), .B2(n_1223), .C(n_1486), .Y(n_1485) );
OAI211xp5_ASAP7_75t_L g973 ( .A1(n_89), .A2(n_900), .B(n_974), .C(n_982), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_90), .A2(n_273), .B1(n_563), .B2(n_945), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_90), .A2(n_113), .B1(n_875), .B2(n_1191), .Y(n_1192) );
AOI22xp5_ASAP7_75t_SL g1273 ( .A1(n_91), .A2(n_265), .B1(n_1259), .B2(n_1264), .Y(n_1273) );
INVx1_ASAP7_75t_L g365 ( .A(n_92), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_92), .A2(n_227), .B1(n_428), .B2(n_430), .C(n_433), .Y(n_427) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_93), .Y(n_292) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_93), .B(n_290), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_95), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g1489 ( .A1(n_96), .A2(n_805), .B(n_1490), .Y(n_1489) );
AOI221xp5_ASAP7_75t_SL g565 ( .A1(n_97), .A2(n_275), .B1(n_522), .B2(n_566), .C(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g657 ( .A(n_98), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_99), .A2(n_714), .B(n_715), .C(n_716), .Y(n_713) );
INVxp33_ASAP7_75t_SL g737 ( .A(n_99), .Y(n_737) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_100), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_101), .Y(n_774) );
INVx1_ASAP7_75t_L g1252 ( .A(n_102), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_102), .B(n_1258), .Y(n_1260) );
AOI22xp33_ASAP7_75t_SL g1268 ( .A1(n_103), .A2(n_112), .B1(n_1253), .B2(n_1259), .Y(n_1268) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_104), .A2(n_244), .B1(n_468), .B2(n_471), .Y(n_467) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_104), .Y(n_477) );
INVxp67_ASAP7_75t_SL g1179 ( .A(n_105), .Y(n_1179) );
AOI22xp33_ASAP7_75t_SL g1194 ( .A1(n_105), .A2(n_218), .B1(n_437), .B2(n_1195), .Y(n_1194) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_106), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_107), .A2(n_182), .B1(n_894), .B2(n_895), .C(n_898), .Y(n_893) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_108), .A2(n_174), .B1(n_880), .B2(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g911 ( .A(n_108), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_109), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_110), .A2(n_276), .B1(n_1249), .B2(n_1253), .Y(n_1248) );
XNOR2xp5_ASAP7_75t_L g1457 ( .A(n_110), .B(n_1458), .Y(n_1457) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_110), .A2(n_1498), .B1(n_1501), .B2(n_1535), .Y(n_1497) );
AOI221xp5_ASAP7_75t_L g1180 ( .A1(n_113), .A2(n_230), .B1(n_558), .B2(n_898), .C(n_1181), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_114), .Y(n_1077) );
INVx1_ASAP7_75t_L g424 ( .A(n_115), .Y(n_424) );
INVx2_ASAP7_75t_L g435 ( .A(n_115), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_115), .B(n_426), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_116), .A2(n_158), .B1(n_410), .B2(n_438), .Y(n_517) );
INVx1_ASAP7_75t_L g532 ( .A(n_116), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g971 ( .A1(n_117), .A2(n_560), .B(n_824), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_117), .A2(n_171), .B1(n_439), .B2(n_616), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_118), .A2(n_183), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g1125 ( .A1(n_118), .A2(n_183), .B1(n_1126), .B2(n_1129), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g1265 ( .A1(n_119), .A2(n_248), .B1(n_1249), .B2(n_1256), .Y(n_1265) );
INVx1_ASAP7_75t_L g387 ( .A(n_120), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_121), .A2(n_154), .B1(n_319), .B2(n_326), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_121), .A2(n_213), .B1(n_437), .B2(n_439), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_122), .A2(n_144), .B1(n_570), .B2(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g609 ( .A(n_122), .Y(n_609) );
INVx1_ASAP7_75t_L g665 ( .A(n_123), .Y(n_665) );
NAND2xp33_ASAP7_75t_SL g690 ( .A(n_123), .B(n_522), .Y(n_690) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_125), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_126), .A2(n_148), .B1(n_428), .B2(n_1472), .C(n_1473), .Y(n_1471) );
INVx1_ASAP7_75t_L g780 ( .A(n_127), .Y(n_780) );
INVx1_ASAP7_75t_L g986 ( .A(n_128), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_131), .A2(n_239), .B1(n_1031), .B2(n_1530), .Y(n_1529) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_133), .A2(n_254), .B1(n_417), .B2(n_506), .C(n_507), .Y(n_505) );
XNOR2xp5_ASAP7_75t_L g484 ( .A(n_134), .B(n_485), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_135), .Y(n_1066) );
XOR2x2_ASAP7_75t_L g861 ( .A(n_136), .B(n_862), .Y(n_861) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_137), .A2(n_271), .B1(n_820), .B2(n_823), .C(n_825), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_138), .A2(n_250), .B1(n_796), .B2(n_873), .Y(n_1013) );
OAI211xp5_ASAP7_75t_SL g1095 ( .A1(n_139), .A2(n_1090), .B(n_1096), .C(n_1099), .Y(n_1095) );
INVx1_ASAP7_75t_L g1145 ( .A(n_139), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_140), .A2(n_155), .B1(n_803), .B2(n_935), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_140), .A2(n_188), .B1(n_825), .B2(n_940), .C(n_942), .Y(n_939) );
INVx1_ASAP7_75t_L g984 ( .A(n_141), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_141), .A2(n_189), .B1(n_614), .B2(n_880), .Y(n_999) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_142), .Y(n_1073) );
INVx1_ASAP7_75t_L g839 ( .A(n_143), .Y(n_839) );
INVx1_ASAP7_75t_L g627 ( .A(n_144), .Y(n_627) );
INVx1_ASAP7_75t_L g921 ( .A(n_145), .Y(n_921) );
CKINVDCx16_ASAP7_75t_R g669 ( .A(n_146), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_147), .A2(n_272), .B1(n_468), .B2(n_471), .Y(n_492) );
INVxp33_ASAP7_75t_SL g542 ( .A(n_147), .Y(n_542) );
NAND5xp2_ASAP7_75t_L g548 ( .A(n_149), .B(n_549), .C(n_588), .D(n_612), .E(n_621), .Y(n_548) );
INVx1_ASAP7_75t_L g634 ( .A(n_149), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g1281 ( .A1(n_149), .A2(n_259), .B1(n_1259), .B2(n_1282), .Y(n_1281) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_150), .A2(n_423), .B(n_438), .Y(n_666) );
INVx1_ASAP7_75t_L g692 ( .A(n_151), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_152), .A2(n_178), .B1(n_694), .B2(n_805), .Y(n_1020) );
OAI211xp5_ASAP7_75t_SL g1022 ( .A1(n_152), .A2(n_1023), .B(n_1024), .C(n_1032), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_154), .A2(n_262), .B1(n_402), .B2(n_409), .Y(n_401) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_155), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_156), .Y(n_1076) );
BUFx3_ASAP7_75t_L g408 ( .A(n_157), .Y(n_408) );
INVx1_ASAP7_75t_L g526 ( .A(n_158), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_159), .Y(n_495) );
INVx1_ASAP7_75t_L g866 ( .A(n_161), .Y(n_866) );
INVx1_ASAP7_75t_L g499 ( .A(n_162), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_162), .A2(n_205), .B1(n_521), .B2(n_524), .C(n_525), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_163), .B(n_1236), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_165), .A2(n_264), .B1(n_825), .B2(n_976), .C(n_978), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_165), .A2(n_228), .B1(n_800), .B2(n_803), .Y(n_998) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_166), .A2(n_805), .B(n_806), .Y(n_804) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_167), .Y(n_304) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_168), .A2(n_247), .B1(n_803), .B2(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g487 ( .A(n_169), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_170), .A2(n_212), .B1(n_556), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_170), .A2(n_204), .B1(n_439), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g1482 ( .A1(n_172), .A2(n_267), .B1(n_1030), .B2(n_1031), .Y(n_1482) );
CKINVDCx20_ASAP7_75t_R g1518 ( .A(n_173), .Y(n_1518) );
INVx1_ASAP7_75t_L g910 ( .A(n_174), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_175), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_176), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_177), .A2(n_213), .B1(n_326), .B2(n_361), .C(n_363), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_177), .A2(n_219), .B1(n_416), .B2(n_418), .C(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g1168 ( .A(n_179), .Y(n_1168) );
AOI22xp33_ASAP7_75t_SL g927 ( .A1(n_180), .A2(n_188), .B1(n_418), .B2(n_801), .Y(n_927) );
INVx1_ASAP7_75t_L g951 ( .A(n_180), .Y(n_951) );
INVx1_ASAP7_75t_L g510 ( .A(n_184), .Y(n_510) );
INVx1_ASAP7_75t_L g809 ( .A(n_185), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_186), .Y(n_1061) );
INVx1_ASAP7_75t_L g644 ( .A(n_187), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_187), .B(n_468), .Y(n_646) );
INVx1_ASAP7_75t_L g983 ( .A(n_189), .Y(n_983) );
XOR2xp5_ASAP7_75t_L g1002 ( .A(n_190), .B(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g785 ( .A(n_191), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_192), .A2(n_279), .B1(n_1259), .B2(n_1264), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_193), .A2(n_250), .B1(n_820), .B2(n_823), .C(n_1044), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_194), .A2(n_197), .B1(n_1253), .B2(n_1259), .Y(n_1343) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_195), .A2(n_524), .B(n_560), .Y(n_732) );
INVx1_ASAP7_75t_L g746 ( .A(n_195), .Y(n_746) );
INVx1_ASAP7_75t_L g1104 ( .A(n_196), .Y(n_1104) );
OAI211xp5_ASAP7_75t_L g1132 ( .A1(n_196), .A2(n_1133), .B(n_1135), .C(n_1137), .Y(n_1132) );
XOR2x2_ASAP7_75t_L g1052 ( .A(n_197), .B(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g620 ( .A(n_198), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_199), .Y(n_1507) );
INVxp67_ASAP7_75t_SL g1177 ( .A(n_200), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_200), .A2(n_229), .B1(n_750), .B2(n_1189), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_201), .Y(n_884) );
INVx1_ASAP7_75t_L g1523 ( .A(n_202), .Y(n_1523) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_203), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_204), .A2(n_253), .B1(n_522), .B2(n_558), .C(n_560), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_205), .A2(n_432), .B(n_433), .Y(n_516) );
XOR2x2_ASAP7_75t_L g704 ( .A(n_207), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1519 ( .A(n_208), .Y(n_1519) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_209), .A2(n_263), .B1(n_678), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g748 ( .A(n_209), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_210), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_211), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_212), .A2(n_253), .B1(n_439), .B2(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_R g683 ( .A(n_214), .B(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g1474 ( .A1(n_216), .A2(n_267), .B1(n_796), .B2(n_932), .Y(n_1474) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_218), .A2(n_229), .B1(n_825), .B2(n_940), .C(n_1172), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_219), .A2(n_227), .B1(n_330), .B2(n_334), .C(n_338), .Y(n_329) );
INVx1_ASAP7_75t_L g1228 ( .A(n_220), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_221), .A2(n_242), .B1(n_694), .B2(n_805), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_223), .Y(n_1059) );
INVx1_ASAP7_75t_L g639 ( .A(n_224), .Y(n_639) );
INVx1_ASAP7_75t_L g1206 ( .A(n_225), .Y(n_1206) );
INVx1_ASAP7_75t_L g1007 ( .A(n_226), .Y(n_1007) );
OAI221xp5_ASAP7_75t_SL g1038 ( .A1(n_226), .A2(n_277), .B1(n_851), .B2(n_949), .C(n_1039), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_230), .A2(n_273), .B1(n_875), .B2(n_1191), .Y(n_1190) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_231), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_231), .A2(n_236), .B1(n_455), .B2(n_459), .C(n_462), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_232), .A2(n_271), .B1(n_428), .B2(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_232), .Y(n_845) );
INVx1_ASAP7_75t_L g1465 ( .A(n_233), .Y(n_1465) );
OAI211xp5_ASAP7_75t_SL g493 ( .A1(n_234), .A2(n_449), .B(n_462), .C(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g537 ( .A(n_234), .Y(n_537) );
INVx1_ASAP7_75t_L g1478 ( .A(n_235), .Y(n_1478) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_236), .A2(n_246), .B1(n_345), .B2(n_353), .C(n_358), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_237), .Y(n_718) );
OAI211xp5_ASAP7_75t_L g965 ( .A1(n_238), .A2(n_949), .B(n_966), .C(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g992 ( .A(n_238), .Y(n_992) );
BUFx3_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
INVx1_ASAP7_75t_L g383 ( .A(n_241), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g899 ( .A1(n_242), .A2(n_900), .B(n_901), .C(n_909), .Y(n_899) );
XOR2x2_ASAP7_75t_L g914 ( .A(n_243), .B(n_915), .Y(n_914) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_244), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_245), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_246), .A2(n_249), .B1(n_441), .B2(n_445), .Y(n_440) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_247), .Y(n_891) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_249), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g1070 ( .A(n_251), .Y(n_1070) );
INVx1_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
INVx2_ASAP7_75t_L g348 ( .A(n_252), .Y(n_348) );
INVx1_ASAP7_75t_L g373 ( .A(n_252), .Y(n_373) );
INVx1_ASAP7_75t_L g527 ( .A(n_254), .Y(n_527) );
INVx1_ASAP7_75t_L g654 ( .A(n_255), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_255), .A2(n_281), .B1(n_556), .B2(n_563), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_256), .B(n_524), .Y(n_723) );
INVx1_ASAP7_75t_L g1479 ( .A(n_257), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_258), .A2(n_260), .B1(n_1256), .B2(n_1259), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1532 ( .A1(n_261), .A2(n_805), .B(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g364 ( .A(n_262), .Y(n_364) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_263), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_266), .Y(n_504) );
INVx1_ASAP7_75t_L g1033 ( .A(n_268), .Y(n_1033) );
INVx1_ASAP7_75t_L g857 ( .A(n_269), .Y(n_857) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_272), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_274), .Y(n_717) );
INVx1_ASAP7_75t_L g1008 ( .A(n_277), .Y(n_1008) );
INVx1_ASAP7_75t_L g729 ( .A(n_278), .Y(n_729) );
INVx1_ASAP7_75t_L g663 ( .A(n_281), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_308), .B(n_1241), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx4f_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_287), .B(n_296), .Y(n_1496) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1500 ( .A(n_289), .B(n_292), .Y(n_1500) );
INVx1_ASAP7_75t_L g1538 ( .A(n_289), .Y(n_1538) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g1540 ( .A(n_292), .B(n_1538), .Y(n_1540) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_296), .B(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g340 ( .A(n_297), .B(n_307), .Y(n_340) );
AND2x4_ASAP7_75t_L g561 ( .A(n_297), .B(n_306), .Y(n_561) );
INVx1_ASAP7_75t_L g1118 ( .A(n_298), .Y(n_1118) );
AND2x4_ASAP7_75t_SL g1495 ( .A(n_298), .B(n_1496), .Y(n_1495) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
OR2x6_ASAP7_75t_L g1110 ( .A(n_300), .B(n_1111), .Y(n_1110) );
INVxp67_ASAP7_75t_L g1236 ( .A(n_300), .Y(n_1236) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_301), .Y(n_571) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx2_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
NAND2x1_ASAP7_75t_L g337 ( .A(n_303), .B(n_304), .Y(n_337) );
INVx1_ASAP7_75t_L g356 ( .A(n_303), .Y(n_356) );
AND2x2_ASAP7_75t_L g481 ( .A(n_303), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g523 ( .A(n_303), .B(n_304), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_304), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g332 ( .A(n_304), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
INVx1_ASAP7_75t_L g377 ( .A(n_304), .Y(n_377) );
AND2x2_ASAP7_75t_L g386 ( .A(n_304), .B(n_325), .Y(n_386) );
INVx2_ASAP7_75t_L g482 ( .A(n_304), .Y(n_482) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g1098 ( .A(n_306), .Y(n_1098) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_307), .Y(n_1102) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_307), .B(n_355), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_958), .B1(n_1239), .B2(n_1240), .Y(n_308) );
INVx1_ASAP7_75t_L g1239 ( .A(n_309), .Y(n_1239) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_860), .B1(n_956), .B2(n_957), .Y(n_309) );
XOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_544), .Y(n_310) );
XNOR2x1_ASAP7_75t_L g957 ( .A(n_311), .B(n_544), .Y(n_957) );
BUFx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
XNOR2x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_484), .Y(n_313) );
XNOR2x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_483), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_399), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_369), .C(n_392), .Y(n_316) );
AOI211xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_329), .B(n_344), .C(n_360), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_320), .A2(n_327), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_950) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_320), .Y(n_1178) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g528 ( .A(n_322), .Y(n_528) );
INVx4_ASAP7_75t_L g721 ( .A(n_322), .Y(n_721) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_322), .Y(n_850) );
INVx1_ASAP7_75t_L g1041 ( .A(n_322), .Y(n_1041) );
INVx8_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g362 ( .A(n_323), .Y(n_362) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_323), .B(n_1102), .Y(n_1116) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_328), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_525) );
OAI22x1_ASAP7_75t_SL g531 ( .A1(n_328), .A2(n_504), .B1(n_528), .B2(n_532), .Y(n_531) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_328), .Y(n_1089) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_331), .A2(n_335), .B1(n_364), .B2(n_365), .C(n_366), .Y(n_363) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g688 ( .A(n_332), .Y(n_688) );
BUFx2_ASAP7_75t_L g720 ( .A(n_332), .Y(n_720) );
BUFx2_ASAP7_75t_L g842 ( .A(n_332), .Y(n_842) );
AND2x2_ASAP7_75t_L g376 ( .A(n_333), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_333), .Y(n_578) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_335), .A2(n_561), .B1(n_839), .B2(n_840), .C(n_843), .Y(n_838) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x6_ASAP7_75t_L g358 ( .A(n_336), .B(n_359), .Y(n_358) );
INVx4_ASAP7_75t_L g573 ( .A(n_336), .Y(n_573) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_336), .Y(n_584) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g390 ( .A(n_337), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_338), .A2(n_358), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_SL g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x4_ASAP7_75t_L g533 ( .A(n_340), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g567 ( .A(n_340), .Y(n_567) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_340), .B(n_723), .C(n_724), .D(n_726), .Y(n_722) );
INVx1_ASAP7_75t_SL g825 ( .A(n_340), .Y(n_825) );
INVx4_ASAP7_75t_L g908 ( .A(n_340), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_340), .B(n_534), .Y(n_1093) );
INVx1_ASAP7_75t_L g535 ( .A(n_341), .Y(n_535) );
OR2x2_ASAP7_75t_L g618 ( .A(n_341), .B(n_444), .Y(n_618) );
OR2x2_ASAP7_75t_L g744 ( .A(n_341), .B(n_434), .Y(n_744) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_341), .Y(n_1157) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g357 ( .A(n_342), .Y(n_357) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g538 ( .A(n_345), .Y(n_538) );
INVx2_ASAP7_75t_SL g682 ( .A(n_345), .Y(n_682) );
NAND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
INVx1_ASAP7_75t_L g359 ( .A(n_346), .Y(n_359) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
BUFx2_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
INVx2_ASAP7_75t_L g475 ( .A(n_348), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_349), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_349), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g581 ( .A(n_349), .Y(n_581) );
AND2x6_ASAP7_75t_L g831 ( .A(n_349), .B(n_522), .Y(n_831) );
AND2x2_ASAP7_75t_L g967 ( .A(n_349), .B(n_575), .Y(n_967) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g575 ( .A(n_352), .Y(n_575) );
INVx1_ASAP7_75t_L g854 ( .A(n_352), .Y(n_854) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_352), .B(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_SL g680 ( .A(n_353), .Y(n_680) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
OR2x2_ASAP7_75t_L g540 ( .A(n_354), .B(n_357), .Y(n_540) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
INVxp67_ASAP7_75t_L g587 ( .A(n_357), .Y(n_587) );
INVx1_ASAP7_75t_L g1123 ( .A(n_357), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_358), .Y(n_543) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_366), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_366), .B(n_676), .Y(n_675) );
INVx4_ASAP7_75t_L g1079 ( .A(n_366), .Y(n_1079) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OR2x6_ASAP7_75t_L g602 ( .A(n_367), .B(n_423), .Y(n_602) );
INVx1_ASAP7_75t_L g701 ( .A(n_367), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_378), .B1(n_379), .B2(n_387), .C1(n_388), .C2(n_391), .Y(n_369) );
AOI21xp33_ASAP7_75t_SL g541 ( .A1(n_370), .A2(n_542), .B(n_543), .Y(n_541) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g605 ( .A(n_372), .B(n_452), .Y(n_605) );
OR2x2_ASAP7_75t_L g699 ( .A(n_372), .B(n_375), .Y(n_699) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_373), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g754 ( .A(n_373), .Y(n_754) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g398 ( .A(n_376), .B(n_382), .Y(n_398) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_376), .Y(n_555) );
INVx3_ASAP7_75t_L g564 ( .A(n_376), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g536 ( .A1(n_379), .A2(n_495), .B1(n_510), .B2(n_537), .C1(n_538), .C2(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g695 ( .A(n_379), .Y(n_695) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_384), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g389 ( .A(n_381), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g684 ( .A(n_381), .B(n_390), .Y(n_684) );
AND2x2_ASAP7_75t_L g479 ( .A(n_382), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g552 ( .A(n_382), .B(n_384), .Y(n_552) );
BUFx2_ASAP7_75t_L g582 ( .A(n_382), .Y(n_582) );
AND2x4_ASAP7_75t_SL g711 ( .A(n_382), .B(n_522), .Y(n_711) );
AND2x4_ASAP7_75t_L g817 ( .A(n_382), .B(n_480), .Y(n_817) );
AND2x4_ASAP7_75t_L g833 ( .A(n_382), .B(n_678), .Y(n_833) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_383), .Y(n_1111) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g945 ( .A(n_385), .Y(n_945) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g556 ( .A(n_386), .Y(n_556) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_386), .Y(n_678) );
BUFx3_ASAP7_75t_L g830 ( .A(n_386), .Y(n_830) );
AOI211xp5_ASAP7_75t_L g447 ( .A1(n_387), .A2(n_448), .B(n_454), .C(n_467), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g519 ( .A1(n_388), .A2(n_496), .B1(n_520), .B2(n_529), .C1(n_530), .C2(n_533), .Y(n_519) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g731 ( .A(n_390), .Y(n_731) );
BUFx2_ASAP7_75t_SL g1090 ( .A(n_390), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_395), .B(n_763), .Y(n_762) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_396), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_396), .A2(n_478), .B1(n_643), .B2(n_644), .Y(n_642) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x4_ASAP7_75t_L g478 ( .A(n_397), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g816 ( .A(n_398), .Y(n_816) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_398), .Y(n_947) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_447), .B(n_473), .C(n_476), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_415), .B1(n_427), .B2(n_436), .C(n_440), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x6_ASAP7_75t_SL g468 ( .A(n_403), .B(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g616 ( .A(n_403), .Y(n_616) );
BUFx2_ASAP7_75t_L g874 ( .A(n_403), .Y(n_874) );
BUFx2_ASAP7_75t_L g933 ( .A(n_403), .Y(n_933) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_404), .Y(n_432) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_404), .Y(n_596) );
BUFx8_ASAP7_75t_L g811 ( .A(n_404), .Y(n_811) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
AND2x4_ASAP7_75t_L g420 ( .A(n_407), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_408), .Y(n_411) );
AND2x4_ASAP7_75t_L g417 ( .A(n_408), .B(n_413), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_408), .B(n_414), .Y(n_503) );
OR2x2_ASAP7_75t_L g650 ( .A(n_408), .B(n_422), .Y(n_650) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx12f_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
AND2x4_ASAP7_75t_L g472 ( .A(n_410), .B(n_470), .Y(n_472) );
INVx5_ASAP7_75t_L g794 ( .A(n_410), .Y(n_794) );
BUFx3_ASAP7_75t_L g875 ( .A(n_410), .Y(n_875) );
BUFx3_ASAP7_75t_L g930 ( .A(n_410), .Y(n_930) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx2_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_411), .B(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g1141 ( .A(n_411), .Y(n_1141) );
INVx1_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g465 ( .A(n_414), .Y(n_465) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g429 ( .A(n_417), .Y(n_429) );
AND2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_443), .Y(n_446) );
BUFx2_ASAP7_75t_L g593 ( .A(n_417), .Y(n_593) );
BUFx2_ASAP7_75t_L g611 ( .A(n_417), .Y(n_611) );
BUFx2_ASAP7_75t_L g803 ( .A(n_417), .Y(n_803) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_417), .B(n_425), .Y(n_1136) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_417), .Y(n_1189) );
INVx8_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_419), .Y(n_506) );
INVx2_ASAP7_75t_L g625 ( .A(n_419), .Y(n_625) );
INVx3_ASAP7_75t_L g800 ( .A(n_419), .Y(n_800) );
INVx2_ASAP7_75t_L g1472 ( .A(n_419), .Y(n_1472) );
INVx8_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AND2x2_ASAP7_75t_L g442 ( .A(n_420), .B(n_443), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_420), .B(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g750 ( .A(n_420), .Y(n_750) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_420), .Y(n_759) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g508 ( .A(n_423), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND3x1_ASAP7_75t_L g753 ( .A(n_424), .B(n_425), .C(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_L g452 ( .A(n_425), .B(n_453), .Y(n_452) );
OR2x4_ASAP7_75t_L g1128 ( .A(n_425), .B(n_650), .Y(n_1128) );
INVx1_ASAP7_75t_L g1131 ( .A(n_425), .Y(n_1131) );
OR2x6_ASAP7_75t_L g1151 ( .A(n_425), .B(n_1152), .Y(n_1151) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp33_ASAP7_75t_SL g434 ( .A(n_426), .B(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g591 ( .A(n_426), .Y(n_591) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g600 ( .A(n_429), .Y(n_600) );
INVx1_ASAP7_75t_L g1195 ( .A(n_429), .Y(n_1195) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_431), .A2(n_499), .B1(n_500), .B2(n_504), .C(n_505), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_431), .A2(n_463), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_655) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g660 ( .A(n_432), .Y(n_660) );
INVx5_ASAP7_75t_L g756 ( .A(n_432), .Y(n_756) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g453 ( .A(n_435), .Y(n_453) );
AND3x4_ASAP7_75t_L g590 ( .A(n_435), .B(n_475), .C(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g658 ( .A(n_435), .B(n_591), .Y(n_658) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_435), .Y(n_1155) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g796 ( .A(n_439), .Y(n_796) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_442), .A2(n_446), .B1(n_487), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g586 ( .A(n_451), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g694 ( .A(n_451), .B(n_587), .Y(n_694) );
AND2x6_ASAP7_75t_L g456 ( .A(n_452), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g460 ( .A(n_452), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g466 ( .A(n_452), .Y(n_466) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_456), .A2(n_460), .B1(n_495), .B2(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_457), .B(n_605), .Y(n_604) );
NAND2x1_ASAP7_75t_L g740 ( .A(n_457), .B(n_605), .Y(n_740) );
AND2x2_ASAP7_75t_L g781 ( .A(n_457), .B(n_605), .Y(n_781) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_457), .B(n_605), .Y(n_1198) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g608 ( .A(n_461), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_462), .A2(n_648), .B1(n_655), .B2(n_659), .C(n_664), .Y(n_647) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_464), .Y(n_515) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_464), .Y(n_1072) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_465), .Y(n_1144) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_470), .Y(n_671) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_472), .B(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_473), .Y(n_734) );
INVx1_ASAP7_75t_L g1046 ( .A(n_473), .Y(n_1046) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21x1_ASAP7_75t_L g549 ( .A1(n_474), .A2(n_550), .B(n_585), .Y(n_549) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_474), .Y(n_955) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI31xp33_ASAP7_75t_SL g491 ( .A1(n_475), .A2(n_492), .A3(n_493), .B(n_497), .Y(n_491) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_475), .A2(n_646), .A3(n_647), .B(n_667), .Y(n_645) );
INVx2_ASAP7_75t_SL g913 ( .A(n_475), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_478), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g619 ( .A(n_478), .Y(n_619) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_480), .Y(n_824) );
INVx2_ASAP7_75t_L g897 ( .A(n_480), .Y(n_897) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
INVx2_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
AND2x4_ASAP7_75t_L g1120 ( .A(n_481), .B(n_1111), .Y(n_1120) );
AOI211x1_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_488), .C(n_518), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_509), .C(n_511), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_500), .A2(n_729), .B1(n_756), .B2(n_757), .C(n_758), .Y(n_755) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g629 ( .A(n_501), .B(n_618), .Y(n_629) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_502), .Y(n_653) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g1152 ( .A(n_503), .Y(n_1152) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI211xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_516), .C(n_517), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_513), .A2(n_665), .B(n_666), .Y(n_664) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g1062 ( .A(n_514), .Y(n_1062) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g623 ( .A(n_515), .B(n_618), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_536), .C(n_541), .Y(n_518) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx3_ASAP7_75t_L g727 ( .A(n_522), .Y(n_727) );
BUFx3_ASAP7_75t_L g894 ( .A(n_522), .Y(n_894) );
INVx1_ASAP7_75t_L g941 ( .A(n_522), .Y(n_941) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_522), .Y(n_978) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_522), .B(n_1098), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g822 ( .A(n_523), .Y(n_822) );
INVx1_ASAP7_75t_L g977 ( .A(n_524), .Y(n_977) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_524), .Y(n_1028) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g805 ( .A(n_540), .B(n_623), .Y(n_805) );
AND2x4_ASAP7_75t_L g988 ( .A(n_540), .B(n_623), .Y(n_988) );
AO22x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_771), .B1(n_858), .B2(n_859), .Y(n_544) );
INVx1_ASAP7_75t_L g858 ( .A(n_545), .Y(n_858) );
XNOR2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_704), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_638), .B1(n_702), .B2(n_703), .Y(n_546) );
INVx1_ASAP7_75t_L g703 ( .A(n_547), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_631), .C(n_635), .Y(n_547) );
INVx1_ASAP7_75t_L g632 ( .A(n_549), .Y(n_632) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .B1(n_562), .B2(n_565), .Y(n_553) );
INVx3_ASAP7_75t_L g981 ( .A(n_555), .Y(n_981) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g566 ( .A(n_559), .Y(n_566) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g898 ( .A(n_561), .Y(n_898) );
INVx2_ASAP7_75t_L g1044 ( .A(n_561), .Y(n_1044) );
INVx1_ASAP7_75t_L g1486 ( .A(n_561), .Y(n_1486) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g725 ( .A(n_564), .Y(n_725) );
INVx2_ASAP7_75t_L g827 ( .A(n_564), .Y(n_827) );
INVx1_ASAP7_75t_L g903 ( .A(n_564), .Y(n_903) );
INVx2_ASAP7_75t_L g1030 ( .A(n_564), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1530 ( .A(n_564), .Y(n_1530) );
INVx2_ASAP7_75t_L g943 ( .A(n_566), .Y(n_943) );
INVx1_ASAP7_75t_L g1173 ( .A(n_566), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_566), .Y(n_1234) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_580), .B1(n_582), .B2(n_583), .Y(n_568) );
INVx2_ASAP7_75t_SL g1082 ( .A(n_570), .Y(n_1082) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g714 ( .A(n_571), .Y(n_714) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_571), .Y(n_847) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g715 ( .A(n_573), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_577), .B2(n_579), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_575), .A2(n_577), .B1(n_717), .B2(n_718), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_576), .A2(n_604), .B1(n_606), .B2(n_609), .C(n_610), .Y(n_603) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_579), .A2(n_622), .B1(n_624), .B2(n_627), .C1(n_628), .C2(n_630), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_580), .A2(n_582), .B1(n_713), .B2(n_719), .Y(n_712) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2x1_ASAP7_75t_L g853 ( .A(n_581), .B(n_854), .Y(n_853) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_584), .A2(n_970), .B(n_971), .C(n_972), .Y(n_969) );
INVx5_ASAP7_75t_L g769 ( .A(n_586), .Y(n_769) );
INVx3_ASAP7_75t_L g1460 ( .A(n_586), .Y(n_1460) );
INVx1_ASAP7_75t_L g633 ( .A(n_588), .Y(n_633) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_603), .Y(n_588) );
AOI33xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .A3(n_594), .B1(n_597), .B2(n_599), .B3(n_601), .Y(n_589) );
BUFx3_ASAP7_75t_L g788 ( .A(n_590), .Y(n_788) );
AOI33xp33_ASAP7_75t_L g868 ( .A1(n_590), .A2(n_869), .A3(n_872), .B1(n_876), .B2(n_877), .B3(n_878), .Y(n_868) );
AOI33xp33_ASAP7_75t_L g993 ( .A1(n_590), .A2(n_994), .A3(n_995), .B1(n_996), .B2(n_997), .B3(n_998), .Y(n_993) );
AOI33xp33_ASAP7_75t_L g1187 ( .A1(n_590), .A2(n_1188), .A3(n_1190), .B1(n_1192), .B2(n_1193), .B3(n_1194), .Y(n_1187) );
INVx3_ASAP7_75t_L g1140 ( .A(n_591), .Y(n_1140) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_596), .Y(n_598) );
INVx2_ASAP7_75t_L g1065 ( .A(n_596), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_596), .B(n_1131), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_600), .A2(n_625), .B1(n_643), .B2(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g997 ( .A(n_602), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_604), .A2(n_606), .B1(n_968), .B2(n_992), .Y(n_991) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_605), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g610 ( .A(n_605), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g741 ( .A(n_605), .B(n_607), .Y(n_741) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx3_ASAP7_75t_L g770 ( .A(n_610), .Y(n_770) );
INVx3_ASAP7_75t_L g786 ( .A(n_610), .Y(n_786) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_610), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_611), .Y(n_1011) );
INVx1_ASAP7_75t_L g637 ( .A(n_612), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_620), .Y(n_612) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_619), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVxp67_ASAP7_75t_L g766 ( .A(n_617), .Y(n_766) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g626 ( .A(n_618), .Y(n_626) );
INVx1_ASAP7_75t_L g636 ( .A(n_621), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_622), .A2(n_628), .B1(n_718), .B2(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_624), .A2(n_810), .B1(n_924), .B2(n_925), .Y(n_923) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x4_ASAP7_75t_L g808 ( .A(n_625), .B(n_626), .Y(n_808) );
AND2x4_ASAP7_75t_L g810 ( .A(n_626), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g776 ( .A(n_629), .B(n_699), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_634), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_634), .A2(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g702 ( .A(n_638), .Y(n_702) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_672), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_652), .B2(n_654), .Y(n_648) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_649), .Y(n_1060) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g765 ( .A(n_650), .Y(n_765) );
OR2x4_ASAP7_75t_L g1149 ( .A(n_650), .B(n_1131), .Y(n_1149) );
OAI22xp33_ASAP7_75t_L g1075 ( .A1(n_652), .A2(n_1060), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g662 ( .A(n_653), .Y(n_662) );
INVx3_ASAP7_75t_L g747 ( .A(n_653), .Y(n_747) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_656), .A2(n_687), .B(n_689), .C(n_690), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_660), .A2(n_746), .B1(n_747), .B2(n_748), .C(n_749), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_662), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_669), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_691), .C(n_696), .Y(n_672) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_683), .C(n_685), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_677), .B(n_679), .Y(n_674) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
BUFx2_ASAP7_75t_L g856 ( .A(n_701), .Y(n_856) );
INVx1_ASAP7_75t_L g1182 ( .A(n_701), .Y(n_1182) );
AND5x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_738), .C(n_760), .D(n_767), .E(n_770), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_734), .B(n_735), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .C(n_722), .D(n_728), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AOI221x1_ASAP7_75t_L g738 ( .A1(n_709), .A2(n_717), .B1(n_739), .B2(n_741), .C(n_742), .Y(n_738) );
AOI222xp33_ASAP7_75t_L g1483 ( .A1(n_710), .A2(n_1465), .B1(n_1466), .B2(n_1484), .C1(n_1485), .C2(n_1487), .Y(n_1483) );
AOI222xp33_ASAP7_75t_L g1528 ( .A1(n_710), .A2(n_1487), .B1(n_1518), .B2(n_1519), .C1(n_1529), .C2(n_1531), .Y(n_1528) );
BUFx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g837 ( .A(n_711), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_720), .A2(n_730), .B1(n_1064), .B2(n_1070), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_720), .A2(n_1061), .B1(n_1077), .B2(n_1083), .Y(n_1086) );
INVx2_ASAP7_75t_L g1084 ( .A(n_721), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B(n_732), .C(n_733), .Y(n_728) );
INVx5_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_739), .A2(n_741), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_739), .A2(n_741), .B1(n_921), .B2(n_922), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_739), .A2(n_741), .B1(n_1518), .B2(n_1519), .Y(n_1517) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AO22x1_ASAP7_75t_L g779 ( .A1(n_741), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_741), .A2(n_781), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_741), .A2(n_1197), .B1(n_1198), .B2(n_1199), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_741), .A2(n_781), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_741), .A2(n_781), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_745), .B1(n_751), .B2(n_755), .Y(n_742) );
BUFx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx4f_ASAP7_75t_L g1057 ( .A(n_744), .Y(n_1057) );
INVx2_ASAP7_75t_SL g791 ( .A(n_750), .Y(n_791) );
INVx1_ASAP7_75t_L g871 ( .A(n_750), .Y(n_871) );
BUFx3_ASAP7_75t_L g935 ( .A(n_750), .Y(n_935) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_752), .Y(n_1015) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g798 ( .A(n_753), .Y(n_798) );
INVx8_ASAP7_75t_L g1069 ( .A(n_756), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
OR2x6_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
OR2x2_ASAP7_75t_L g880 ( .A(n_764), .B(n_766), .Y(n_880) );
INVx2_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_769), .B(n_785), .Y(n_784) );
INVx2_ASAP7_75t_SL g882 ( .A(n_770), .Y(n_882) );
NAND4xp75_ASAP7_75t_L g915 ( .A(n_770), .B(n_916), .C(n_919), .D(n_936), .Y(n_915) );
AND4x1_ASAP7_75t_L g1183 ( .A(n_770), .B(n_1184), .C(n_1187), .D(n_1196), .Y(n_1183) );
NAND3xp33_ASAP7_75t_SL g1463 ( .A(n_770), .B(n_1464), .C(n_1467), .Y(n_1463) );
NAND3xp33_ASAP7_75t_SL g1508 ( .A(n_770), .B(n_1509), .C(n_1517), .Y(n_1508) );
INVx2_ASAP7_75t_L g859 ( .A(n_771), .Y(n_859) );
XOR2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_857), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_773), .B(n_812), .Y(n_772) );
AOI211x1_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B(n_777), .C(n_804), .Y(n_773) );
AOI21xp33_ASAP7_75t_SL g883 ( .A1(n_775), .A2(n_884), .B(n_885), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_775), .A2(n_917), .B(n_918), .Y(n_916) );
AOI21xp33_ASAP7_75t_L g985 ( .A1(n_775), .A2(n_986), .B(n_987), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_775), .A2(n_1019), .B(n_1020), .Y(n_1018) );
AOI21xp33_ASAP7_75t_L g1162 ( .A1(n_775), .A2(n_1163), .B(n_1164), .Y(n_1162) );
AOI21xp5_ASAP7_75t_L g1215 ( .A1(n_775), .A2(n_1216), .B(n_1217), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_775), .A2(n_1460), .B1(n_1461), .B2(n_1462), .C(n_1463), .Y(n_1459) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_775), .A2(n_1460), .B1(n_1506), .B2(n_1507), .C(n_1508), .Y(n_1505) );
INVx8_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_787), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_783), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_784), .B(n_786), .Y(n_783) );
NAND2xp5_ASAP7_75t_R g832 ( .A(n_785), .B(n_833), .Y(n_832) );
AOI33xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .A3(n_792), .B1(n_795), .B2(n_797), .B3(n_799), .Y(n_787) );
AOI33xp33_ASAP7_75t_L g926 ( .A1(n_788), .A2(n_877), .A3(n_927), .B1(n_928), .B2(n_931), .B3(n_934), .Y(n_926) );
AOI33xp33_ASAP7_75t_L g1009 ( .A1(n_788), .A2(n_1010), .A3(n_1012), .B1(n_1013), .B2(n_1014), .B3(n_1016), .Y(n_1009) );
AOI33xp33_ASAP7_75t_L g1208 ( .A1(n_788), .A2(n_1209), .A3(n_1210), .B1(n_1211), .B2(n_1212), .B3(n_1213), .Y(n_1208) );
INVx1_ASAP7_75t_L g1473 ( .A(n_788), .Y(n_1473) );
AOI33xp33_ASAP7_75t_L g1509 ( .A1(n_788), .A2(n_1014), .A3(n_1510), .B1(n_1511), .B2(n_1515), .B3(n_1516), .Y(n_1509) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g1514 ( .A(n_794), .Y(n_1514) );
BUFx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g877 ( .A(n_798), .Y(n_877) );
BUFx2_ASAP7_75t_L g1193 ( .A(n_798), .Y(n_1193) );
BUFx2_ASAP7_75t_L g1212 ( .A(n_798), .Y(n_1212) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_807), .A2(n_809), .B1(n_815), .B2(n_817), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_808), .A2(n_810), .B1(n_1478), .B2(n_1479), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_808), .A2(n_810), .B1(n_1523), .B2(n_1524), .Y(n_1533) );
INVx2_ASAP7_75t_L g881 ( .A(n_810), .Y(n_881) );
INVx2_ASAP7_75t_L g1186 ( .A(n_810), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_811), .Y(n_929) );
INVx2_ASAP7_75t_SL g1513 ( .A(n_811), .Y(n_1513) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_834), .B(n_855), .Y(n_812) );
NAND3xp33_ASAP7_75t_SL g813 ( .A(n_814), .B(n_818), .C(n_832), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_815), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_815), .A2(n_1036), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_817), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_817), .A2(n_924), .B1(n_925), .B2(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1037 ( .A(n_817), .Y(n_1037) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_826), .B(n_831), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g1233 ( .A(n_821), .Y(n_1233) );
BUFx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g907 ( .A(n_822), .Y(n_907) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_830), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_831), .A2(n_902), .B(n_904), .Y(n_901) );
AOI21xp5_ASAP7_75t_SL g938 ( .A1(n_831), .A2(n_939), .B(n_944), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g974 ( .A1(n_831), .A2(n_975), .B(n_979), .Y(n_974) );
AOI21xp5_ASAP7_75t_L g1024 ( .A1(n_831), .A2(n_1025), .B(n_1029), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g1170 ( .A1(n_831), .A2(n_1171), .B(n_1174), .Y(n_1170) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_831), .A2(n_1221), .B(n_1226), .Y(n_1220) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_831), .A2(n_833), .B1(n_1461), .B2(n_1481), .C(n_1482), .Y(n_1480) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_831), .A2(n_833), .B1(n_1506), .B2(n_1526), .C(n_1527), .Y(n_1525) );
INVx2_ASAP7_75t_SL g900 ( .A(n_833), .Y(n_900) );
INVx3_ASAP7_75t_L g1023 ( .A(n_833), .Y(n_1023) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g888 ( .A(n_836), .Y(n_888) );
INVx2_ASAP7_75t_L g949 ( .A(n_836), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_836), .A2(n_853), .B1(n_1206), .B2(n_1207), .Y(n_1237) );
INVx4_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx4_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_848), .B2(n_849), .Y(n_844) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_846), .A2(n_849), .B1(n_891), .B2(n_892), .C(n_893), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g1039 ( .A1(n_846), .A2(n_1040), .B1(n_1041), .B2(n_1042), .C(n_1043), .Y(n_1039) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx5_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g889 ( .A(n_853), .Y(n_889) );
OAI21xp5_ASAP7_75t_SL g964 ( .A1(n_855), .A2(n_965), .B(n_973), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g1475 ( .A1(n_855), .A2(n_1476), .B(n_1489), .Y(n_1475) );
AOI21xp5_ASAP7_75t_L g1520 ( .A1(n_855), .A2(n_1521), .B(n_1532), .Y(n_1520) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g956 ( .A(n_860), .Y(n_956) );
XNOR2x1_ASAP7_75t_L g860 ( .A(n_861), .B(n_914), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_883), .C(n_886), .Y(n_862) );
NOR3xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_879), .C(n_882), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g1074 ( .A(n_877), .Y(n_1074) );
NOR3xp33_ASAP7_75t_L g1004 ( .A(n_882), .B(n_1005), .C(n_1017), .Y(n_1004) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_899), .B(n_913), .Y(n_886) );
BUFx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g1225 ( .A(n_897), .Y(n_1225) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_912), .A2(n_947), .B1(n_983), .B2(n_984), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_912), .A2(n_947), .B1(n_1168), .B2(n_1169), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_912), .A2(n_1034), .B1(n_1478), .B2(n_1479), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_912), .A2(n_1034), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
AND3x1_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .C(n_926), .Y(n_919) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
OAI21xp5_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_948), .B(n_955), .Y(n_936) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g954 ( .A(n_941), .Y(n_954) );
INVx1_ASAP7_75t_L g1181 ( .A(n_941), .Y(n_1181) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_947), .Y(n_1034) );
INVxp67_ASAP7_75t_SL g1240 ( .A(n_958), .Y(n_1240) );
XOR2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_1048), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_1001), .B2(n_1047), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_985), .C(n_989), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g1488 ( .A(n_967), .Y(n_1488) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g1027 ( .A(n_978), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_978), .Y(n_1222) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_999), .C(n_1000), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_993), .Y(n_990) );
NOR3xp33_ASAP7_75t_L g1203 ( .A(n_1000), .B(n_1204), .C(n_1214), .Y(n_1203) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1001), .Y(n_1047) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_1002), .Y(n_1001) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1018), .C(n_1021), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1009), .Y(n_1005) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1038), .B(n_1045), .Y(n_1021) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1032) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
OAI21xp5_ASAP7_75t_L g1218 ( .A1(n_1045), .A2(n_1219), .B(n_1230), .Y(n_1218) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1050), .B1(n_1201), .B2(n_1238), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OA22x2_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1052), .B1(n_1158), .B2(n_1159), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NAND3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1094), .C(n_1124), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1078), .Y(n_1054) );
OAI33xp33_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1058), .A3(n_1063), .B1(n_1067), .B2(n_1074), .B3(n_1075), .Y(n_1055) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1060), .B1(n_1061), .B2(n_1062), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_1059), .A2(n_1076), .B1(n_1081), .B2(n_1083), .Y(n_1080) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1065), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_1066), .A2(n_1073), .B1(n_1088), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1070), .B1(n_1071), .B2(n_1073), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1072), .Y(n_1134) );
OAI33xp33_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1080), .A3(n_1085), .B1(n_1086), .B2(n_1087), .B3(n_1091), .Y(n_1078) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
OAI221xp5_ASAP7_75t_L g1176 ( .A1(n_1088), .A2(n_1177), .B1(n_1178), .B2(n_1179), .C(n_1180), .Y(n_1176) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OAI31xp33_ASAP7_75t_SL g1094 ( .A1(n_1095), .A2(n_1107), .A3(n_1117), .B(n_1121), .Y(n_1094) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1103), .B1(n_1104), .B2(n_1105), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_1103), .A2(n_1138), .B1(n_1142), .B2(n_1145), .Y(n_1137) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx3_ASAP7_75t_SL g1119 ( .A(n_1120), .Y(n_1119) );
BUFx3_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
OAI31xp33_ASAP7_75t_SL g1124 ( .A1(n_1125), .A2(n_1132), .A3(n_1146), .B(n_1153), .Y(n_1124) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
CKINVDCx8_ASAP7_75t_R g1135 ( .A(n_1136), .Y(n_1135) );
BUFx3_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_1140), .B(n_1144), .Y(n_1143) );
BUFx6f_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx2_ASAP7_75t_SL g1148 ( .A(n_1149), .Y(n_1148) );
BUFx3_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1156), .Y(n_1153) );
INVx1_ASAP7_75t_SL g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
AO21x2_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B(n_1200), .Y(n_1159) );
NAND3xp33_ASAP7_75t_SL g1161 ( .A(n_1162), .B(n_1165), .C(n_1183), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1175), .B(n_1182), .Y(n_1165) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1193), .B(n_1470), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_1201), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1215), .C(n_1218), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1208), .Y(n_1204) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .Y(n_1231) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1451), .B1(n_1454), .B2(n_1491), .C(n_1497), .Y(n_1241) );
NOR3xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1389), .C(n_1431), .Y(n_1242) );
A2O1A1Ixp33_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1323), .B(n_1341), .C(n_1345), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1270), .B1(n_1278), .B2(n_1289), .C(n_1296), .Y(n_1244) );
AOI221xp5_ASAP7_75t_SL g1390 ( .A1(n_1245), .A2(n_1329), .B1(n_1391), .B2(n_1393), .C(n_1395), .Y(n_1390) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1261), .Y(n_1246) );
INVx3_ASAP7_75t_L g1322 ( .A(n_1247), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1331 ( .A(n_1247), .B(n_1312), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1247), .B(n_1262), .Y(n_1333) );
INVx3_ASAP7_75t_L g1347 ( .A(n_1247), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1247), .B(n_1355), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1247), .B(n_1303), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1247), .B(n_1262), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1247), .B(n_1310), .Y(n_1450) );
AND2x4_ASAP7_75t_SL g1247 ( .A(n_1248), .B(n_1255), .Y(n_1247) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1249), .Y(n_1453) );
AND2x6_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1251), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1250), .B(n_1254), .Y(n_1253) );
AND2x4_ASAP7_75t_L g1256 ( .A(n_1250), .B(n_1257), .Y(n_1256) );
AND2x6_ASAP7_75t_L g1259 ( .A(n_1250), .B(n_1260), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1250), .B(n_1254), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1250), .B(n_1254), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g1537 ( .A(n_1251), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1252), .B(n_1258), .Y(n_1257) );
INVx2_ASAP7_75t_SL g1382 ( .A(n_1261), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1266), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1262), .B(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_SL g1297 ( .A(n_1262), .B(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1262), .B(n_1267), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1262), .B(n_1322), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1380 ( .A(n_1262), .B(n_1267), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1430 ( .A(n_1262), .B(n_1342), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1265), .Y(n_1262) );
AND2x4_ASAP7_75t_L g1351 ( .A(n_1263), .B(n_1265), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1266), .B(n_1351), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1266), .B(n_1318), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_1266), .B(n_1293), .Y(n_1423) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1267), .Y(n_1303) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1267), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1269), .Y(n_1267) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1270), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1270), .B(n_1340), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1270), .B(n_1306), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1270), .B(n_1358), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1275), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1271), .B(n_1288), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1271), .B(n_1275), .Y(n_1330) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1271), .Y(n_1372) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1272), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1272), .B(n_1275), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1274), .Y(n_1272) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1275), .Y(n_1288) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1275), .Y(n_1320) );
NOR2xp33_ASAP7_75t_L g1434 ( .A(n_1275), .B(n_1301), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1285), .Y(n_1278) );
OAI22xp33_ASAP7_75t_L g1448 ( .A1(n_1279), .A2(n_1353), .B1(n_1415), .B2(n_1449), .Y(n_1448) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1284), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1280), .B(n_1287), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1280), .B(n_1339), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1283), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1281), .B(n_1283), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1284), .B(n_1309), .Y(n_1308) );
A2O1A1Ixp33_ASAP7_75t_L g1374 ( .A1(n_1285), .A2(n_1375), .B(n_1377), .C(n_1381), .Y(n_1374) );
OAI221xp5_ASAP7_75t_L g1414 ( .A1(n_1285), .A2(n_1415), .B1(n_1416), .B2(n_1417), .C(n_1418), .Y(n_1414) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1286), .B(n_1318), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1287), .B(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1287), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1287), .B(n_1309), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1288), .B(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1354 ( .A(n_1291), .B(n_1319), .Y(n_1354) );
AOI32xp33_ASAP7_75t_L g1363 ( .A1(n_1291), .A2(n_1364), .A3(n_1368), .B1(n_1369), .B2(n_1373), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1291), .B(n_1406), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1291), .B(n_1327), .Y(n_1416) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1292), .B(n_1326), .Y(n_1325) );
NAND2xp5_ASAP7_75t_SL g1349 ( .A(n_1292), .B(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1292), .B(n_1379), .Y(n_1378) );
NAND2xp5_ASAP7_75t_SL g1440 ( .A(n_1292), .B(n_1329), .Y(n_1440) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1293), .B(n_1303), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1293), .B(n_1301), .Y(n_1306) );
INVx3_ASAP7_75t_L g1318 ( .A(n_1293), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1293), .B(n_1301), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1293), .B(n_1322), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1295), .Y(n_1293) );
NAND3xp33_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1304), .C(n_1311), .Y(n_1296) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1302), .Y(n_1298) );
CKINVDCx14_ASAP7_75t_R g1299 ( .A(n_1300), .Y(n_1299) );
AOI32xp33_ASAP7_75t_L g1381 ( .A1(n_1300), .A2(n_1382), .A3(n_1383), .B1(n_1384), .B2(n_1388), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g1309 ( .A(n_1301), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1301), .B(n_1316), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1301), .B(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1301), .B(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1301), .B(n_1372), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1301), .B(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1303), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1303), .B(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1303), .Y(n_1386) );
OAI322xp33_ASAP7_75t_L g1395 ( .A1(n_1303), .A2(n_1352), .A3(n_1355), .B1(n_1396), .B2(n_1397), .C1(n_1400), .C2(n_1401), .Y(n_1395) );
O2A1O1Ixp33_ASAP7_75t_L g1424 ( .A1(n_1303), .A2(n_1425), .B(n_1426), .C(n_1429), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_1303), .A2(n_1307), .B1(n_1436), .B2(n_1438), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1303), .B(n_1437), .Y(n_1436) );
OAI21xp5_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1307), .B(n_1310), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1306), .B(n_1329), .Y(n_1388) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1309), .B(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1309), .B(n_1365), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1309), .B(n_1372), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_1309), .B(n_1440), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1309), .B(n_1327), .Y(n_1447) );
AOI222xp33_ASAP7_75t_L g1432 ( .A1(n_1310), .A2(n_1326), .B1(n_1350), .B2(n_1358), .C1(n_1382), .C2(n_1433), .Y(n_1432) );
A2O1A1Ixp33_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1314), .B(n_1317), .C(n_1321), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1312), .B(n_1321), .Y(n_1373) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1313), .B(n_1326), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1313), .B(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1316), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1318), .Y(n_1340) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1320), .Y(n_1394) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1321), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1322), .B(n_1379), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1322), .B(n_1380), .Y(n_1415) );
NOR3xp33_ASAP7_75t_L g1422 ( .A(n_1322), .B(n_1366), .C(n_1423), .Y(n_1422) );
NOR2xp33_ASAP7_75t_L g1443 ( .A(n_1322), .B(n_1444), .Y(n_1443) );
O2A1O1Ixp33_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1328), .B(n_1331), .C(n_1332), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1327), .B(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1327), .Y(n_1367) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1328), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1329), .B(n_1358), .Y(n_1437) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
OAI21xp5_ASAP7_75t_L g1332 ( .A1(n_1333), .A2(n_1334), .B(n_1335), .Y(n_1332) );
A2O1A1Ixp33_ASAP7_75t_L g1384 ( .A1(n_1333), .A2(n_1385), .B(n_1386), .C(n_1387), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1337), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1336), .B(n_1340), .Y(n_1421) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1340), .B(n_1371), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1340), .B(n_1434), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1341), .B(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1341), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_1341), .A2(n_1411), .B1(n_1412), .B2(n_1414), .C(n_1424), .Y(n_1410) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
OAI221xp5_ASAP7_75t_L g1389 ( .A1(n_1342), .A2(n_1385), .B1(n_1390), .B2(n_1402), .C(n_1410), .Y(n_1389) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1342), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1344), .Y(n_1342) );
AOI211xp5_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1348), .B(n_1359), .C(n_1374), .Y(n_1345) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1347), .Y(n_1400) );
OAI221xp5_ASAP7_75t_L g1348 ( .A1(n_1349), .A2(n_1352), .B1(n_1353), .B2(n_1355), .C(n_1356), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1350), .B(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1350), .Y(n_1404) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1351), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1351), .B(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
OAI21xp33_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1361), .B(n_1363), .Y(n_1359) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1362), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1367), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1398 ( .A(n_1366), .B(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1368), .Y(n_1417) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1383), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1385), .B(n_1400), .Y(n_1441) );
NOR2xp33_ASAP7_75t_L g1407 ( .A(n_1386), .B(n_1408), .Y(n_1407) );
INVxp67_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
AOI31xp33_ASAP7_75t_SL g1418 ( .A1(n_1394), .A2(n_1419), .A3(n_1421), .B(n_1422), .Y(n_1418) );
INVxp67_ASAP7_75t_SL g1397 ( .A(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1399), .Y(n_1446) );
NOR2xp33_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1407), .Y(n_1402) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1405), .Y(n_1403) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
AOI211xp5_ASAP7_75t_L g1442 ( .A1(n_1409), .A2(n_1430), .B(n_1443), .C(n_1448), .Y(n_1442) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
A2O1A1Ixp33_ASAP7_75t_L g1431 ( .A1(n_1432), .A2(n_1435), .B(n_1441), .C(n_1442), .Y(n_1431) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVxp67_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
CKINVDCx20_ASAP7_75t_R g1451 ( .A(n_1452), .Y(n_1451) );
CKINVDCx20_ASAP7_75t_R g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NAND2xp67_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1475), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_1468), .A2(n_1469), .B1(n_1471), .B2(n_1474), .Y(n_1467) );
NAND3xp33_ASAP7_75t_SL g1476 ( .A(n_1477), .B(n_1480), .C(n_1483), .Y(n_1476) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
CKINVDCx20_ASAP7_75t_R g1491 ( .A(n_1492), .Y(n_1491) );
CKINVDCx20_ASAP7_75t_R g1492 ( .A(n_1493), .Y(n_1492) );
INVx3_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
BUFx3_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
HB1xp67_ASAP7_75t_SL g1498 ( .A(n_1499), .Y(n_1498) );
BUFx3_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVxp33_ASAP7_75t_SL g1501 ( .A(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1504), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1520), .Y(n_1504) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
NAND3xp33_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1525), .C(n_1528), .Y(n_1521) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
OAI21xp5_ASAP7_75t_L g1536 ( .A1(n_1537), .A2(n_1538), .B(n_1539), .Y(n_1536) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
endmodule