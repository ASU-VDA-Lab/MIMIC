module fake_jpeg_6562_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_46),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_19),
.C(n_28),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_44),
.B(n_26),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_19),
.B(n_25),
.C(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_25),
.B1(n_38),
.B2(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_15),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_33),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_74),
.B1(n_77),
.B2(n_44),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_21),
.A3(n_20),
.B1(n_39),
.B2(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_25),
.B1(n_37),
.B2(n_29),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_56),
.B1(n_53),
.B2(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_26),
.B1(n_20),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_16),
.A3(n_41),
.B1(n_23),
.B2(n_27),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_45),
.Y(n_83)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_48),
.B(n_42),
.C(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_47),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_103),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_102),
.B1(n_94),
.B2(n_107),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_71),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_43),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_55),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_74),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_45),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_59),
.C(n_52),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_62),
.B1(n_54),
.B2(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_66),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_82),
.B1(n_65),
.B2(n_73),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_133),
.B1(n_78),
.B2(n_51),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_82),
.B(n_59),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_93),
.B(n_49),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_122),
.B(n_93),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_127),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_86),
.B1(n_24),
.B2(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_67),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_100),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_66),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_138),
.B(n_143),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_86),
.B1(n_72),
.B2(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_145),
.B1(n_150),
.B2(n_91),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_154),
.C(n_156),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_108),
.B1(n_78),
.B2(n_75),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_75),
.B1(n_91),
.B2(n_63),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_41),
.C(n_49),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_144),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_63),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_16),
.B(n_23),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_114),
.B(n_118),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_160),
.B(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_164),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_125),
.B1(n_122),
.B2(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_113),
.B1(n_110),
.B2(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_122),
.B1(n_115),
.B2(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_127),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_151),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_156),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_191),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_152),
.C(n_121),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_187),
.C(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_115),
.C(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_181),
.C(n_167),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_148),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_163),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_114),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_197),
.C(n_200),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_158),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_112),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_165),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_110),
.C(n_139),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_112),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_184),
.B1(n_175),
.B2(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_205),
.Y(n_214)
);

XNOR2x2_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_146),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_178),
.B1(n_173),
.B2(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_139),
.C(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_168),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_200),
.B(n_117),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_172),
.B1(n_180),
.B2(n_163),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_168),
.B1(n_132),
.B2(n_91),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_221),
.A2(n_225),
.B(n_226),
.Y(n_229)
);

NOR2x1_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_185),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_164),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_75),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_206),
.B(n_196),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_237),
.B(n_239),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_187),
.B1(n_188),
.B2(n_201),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_191),
.B1(n_195),
.B2(n_186),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_202),
.C(n_197),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_238),
.C(n_233),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_151),
.C(n_134),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_244),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_117),
.B(n_96),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_243),
.B(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_217),
.B1(n_213),
.B2(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_245),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_96),
.B(n_69),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_51),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_1),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_211),
.B(n_242),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_224),
.B(n_210),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_252),
.A2(n_260),
.B(n_261),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_210),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_234),
.B(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_216),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_250),
.Y(n_266)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_252),
.C(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_244),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_271),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_255),
.B(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_268),
.C(n_269),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_216),
.B(n_96),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_216),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_11),
.B(n_14),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_69),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_11),
.C(n_14),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_8),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_11),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_8),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_282),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_16),
.Y(n_279)
);

NOR3xp33_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_280),
.C(n_16),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_16),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_10),
.B(n_14),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_284),
.A3(n_8),
.B1(n_13),
.B2(n_12),
.C1(n_5),
.C2(n_6),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_272),
.B1(n_12),
.B2(n_13),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_290),
.A3(n_291),
.B1(n_2),
.B2(n_3),
.C1(n_23),
.C2(n_27),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_7),
.A3(n_6),
.B1(n_12),
.B2(n_27),
.C1(n_23),
.C2(n_1),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_7),
.A3(n_6),
.B1(n_3),
.B2(n_2),
.C1(n_1),
.C2(n_23),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_277),
.C(n_3),
.Y(n_292)
);

AOI31xp33_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_295),
.A3(n_296),
.B(n_27),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_2),
.B(n_3),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.C(n_27),
.Y(n_299)
);

OAI31xp33_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_27),
.A3(n_41),
.B(n_294),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_27),
.Y(n_300)
);


endmodule