module fake_jpeg_16672_n_395 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_45),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_55),
.Y(n_99)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_23),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_5),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_34),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_94),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_39),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_85),
.B1(n_91),
.B2(n_93),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_98),
.B1(n_26),
.B2(n_33),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_30),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_44),
.A2(n_24),
.B1(n_36),
.B2(n_23),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_36),
.B1(n_60),
.B2(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_34),
.B1(n_31),
.B2(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_111),
.B1(n_14),
.B2(n_33),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_31),
.B1(n_28),
.B2(n_34),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_21),
.Y(n_132)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_42),
.A2(n_33),
.B1(n_26),
.B2(n_14),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_55),
.B1(n_51),
.B2(n_47),
.Y(n_121)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_43),
.A2(n_33),
.B1(n_26),
.B2(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_27),
.Y(n_131)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_41),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_164)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_121),
.A2(n_110),
.B1(n_108),
.B2(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_128),
.Y(n_170)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_127),
.A2(n_149),
.B(n_0),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_79),
.B(n_49),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_13),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_130),
.A2(n_146),
.B1(n_29),
.B2(n_4),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_132),
.B(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_27),
.Y(n_135)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_136),
.A2(n_169),
.B1(n_16),
.B2(n_29),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_26),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_148),
.B1(n_153),
.B2(n_161),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_87),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_27),
.Y(n_142)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_12),
.Y(n_145)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_5),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_92),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_73),
.A2(n_61),
.B(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_46),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_76),
.B(n_21),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_10),
.Y(n_154)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_87),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_158),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_84),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_76),
.B(n_19),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_86),
.B(n_10),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_165),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_96),
.B(n_46),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_16),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_72),
.A2(n_117),
.B1(n_83),
.B2(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_171),
.B(n_123),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_126),
.B1(n_122),
.B2(n_150),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_172),
.A2(n_192),
.B1(n_163),
.B2(n_162),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_72),
.B1(n_97),
.B2(n_114),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_147),
.B1(n_159),
.B2(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_157),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_181),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_118),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_179),
.B(n_188),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_184),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_128),
.B(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_145),
.C(n_152),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_83),
.B1(n_108),
.B2(n_101),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_186),
.A2(n_189),
.B1(n_155),
.B2(n_167),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_77),
.B1(n_101),
.B2(n_19),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_141),
.B1(n_155),
.B2(n_167),
.Y(n_234)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_77),
.B1(n_74),
.B2(n_19),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_199),
.B(n_200),
.Y(n_224)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_205),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_0),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_0),
.B(n_3),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_0),
.B(n_3),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_210),
.B(n_70),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_202),
.B(n_213),
.Y(n_246)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_67),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_67),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_R g210 ( 
.A1(n_130),
.A2(n_29),
.B1(n_70),
.B2(n_4),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_4),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_124),
.C(n_135),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_218),
.B(n_233),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_219),
.A2(n_246),
.B1(n_240),
.B2(n_236),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_172),
.A2(n_193),
.B1(n_182),
.B2(n_170),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_222),
.A2(n_256),
.B1(n_207),
.B2(n_173),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_124),
.A3(n_153),
.B1(n_131),
.B2(n_154),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_226),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_119),
.B(n_120),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_228),
.A2(n_237),
.B(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_146),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_231),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_146),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_165),
.B(n_144),
.C(n_129),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_204),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_138),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g285 ( 
.A1(n_234),
.A2(n_257),
.B(n_256),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_158),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_235),
.B(n_236),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_248),
.B1(n_175),
.B2(n_205),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_144),
.Y(n_242)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_156),
.A3(n_157),
.B1(n_143),
.B2(n_125),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_171),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_185),
.B(n_147),
.C(n_123),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_222),
.C(n_244),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_208),
.B(n_123),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_199),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_203),
.A2(n_147),
.B1(n_159),
.B2(n_195),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_259),
.C(n_269),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_221),
.C(n_226),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_249),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_266),
.B(n_272),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_267),
.B1(n_279),
.B2(n_283),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_203),
.B(n_176),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_189),
.B1(n_173),
.B2(n_212),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_268),
.A2(n_285),
.B1(n_230),
.B2(n_217),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_221),
.B(n_214),
.C(n_192),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_199),
.B(n_214),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_179),
.B(n_174),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_287),
.B(n_241),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_290),
.B1(n_219),
.B2(n_253),
.Y(n_292)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_196),
.B1(n_197),
.B2(n_174),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_177),
.B1(n_183),
.B2(n_186),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_228),
.A2(n_177),
.B1(n_211),
.B2(n_198),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_284),
.A2(n_278),
.B1(n_269),
.B2(n_290),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_235),
.B(n_237),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_231),
.C(n_229),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_309),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_242),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_300),
.C(n_303),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_266),
.A2(n_238),
.B(n_232),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_304),
.B(n_308),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_243),
.B1(n_234),
.B2(n_220),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_297),
.A2(n_312),
.B1(n_316),
.B2(n_265),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_227),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_217),
.Y(n_301)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_R g302 ( 
.A1(n_289),
.A2(n_274),
.B1(n_271),
.B2(n_264),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_313),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_250),
.Y(n_303)
);

NAND2x1p5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_247),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_273),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_310),
.B(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_230),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_282),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_265),
.C(n_272),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_277),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_260),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_264),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_328),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_334),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_333),
.A2(n_299),
.B1(n_304),
.B2(n_307),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_303),
.B(n_262),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_312),
.A2(n_260),
.B1(n_281),
.B2(n_284),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_304),
.B1(n_309),
.B2(n_308),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_341),
.C(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_267),
.C(n_283),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_279),
.C(n_318),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_343),
.B(n_360),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_301),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_SL g372 ( 
.A(n_345),
.B(n_346),
.C(n_352),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_293),
.C(n_323),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_316),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_328),
.C(n_339),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_313),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_350),
.B(n_322),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_355),
.B1(n_331),
.B2(n_336),
.Y(n_365)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_356),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_315),
.B1(n_296),
.B2(n_299),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_317),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_332),
.A2(n_307),
.B(n_293),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_359),
.A2(n_351),
.B(n_350),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_321),
.A2(n_311),
.B1(n_341),
.B2(n_324),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_360),
.A2(n_321),
.B1(n_342),
.B2(n_340),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_363),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_362),
.A2(n_369),
.B(n_370),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_352),
.A2(n_327),
.B1(n_336),
.B2(n_330),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_365),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_367),
.C(n_371),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_311),
.B1(n_339),
.B2(n_359),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_345),
.B(n_349),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_353),
.B1(n_359),
.B2(n_347),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_348),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_376),
.C(n_378),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_354),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_344),
.C(n_354),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_372),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_379),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_368),
.B1(n_372),
.B2(n_369),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_375),
.B1(n_377),
.B2(n_368),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_377),
.A2(n_367),
.B(n_371),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_381),
.C(n_384),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_379),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_390),
.Y(n_391)
);

OAI321xp33_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_389),
.A3(n_362),
.B1(n_386),
.B2(n_387),
.C(n_364),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_346),
.B(n_378),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_SL g394 ( 
.A1(n_393),
.A2(n_363),
.B(n_344),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_348),
.Y(n_395)
);


endmodule