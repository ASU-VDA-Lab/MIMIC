module real_aes_7480_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_0), .A2(n_247), .B1(n_673), .B2(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_1), .A2(n_272), .B1(n_344), .B2(n_349), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_2), .A2(n_108), .B1(n_548), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_3), .A2(n_260), .B1(n_446), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_4), .A2(n_261), .B1(n_508), .B2(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_5), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_6), .B(n_342), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_7), .B(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_8), .A2(n_176), .B1(n_666), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_9), .A2(n_99), .B1(n_354), .B2(n_448), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_10), .A2(n_25), .B1(n_318), .B2(n_329), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_11), .A2(n_165), .B1(n_398), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_12), .A2(n_282), .B1(n_568), .B2(n_765), .Y(n_764) );
XOR2x2_ASAP7_75t_L g624 ( .A(n_13), .B(n_625), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_14), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_15), .A2(n_137), .B1(n_394), .B2(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_16), .A2(n_184), .B1(n_354), .B2(n_606), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_17), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_18), .A2(n_118), .B1(n_398), .B2(n_399), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_19), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_20), .A2(n_226), .B1(n_362), .B2(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_21), .A2(n_139), .B1(n_393), .B2(n_402), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_22), .A2(n_110), .B1(n_133), .B2(n_366), .C1(n_369), .C2(n_374), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_23), .A2(n_191), .B1(n_393), .B2(n_394), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_24), .Y(n_609) );
INVx1_ASAP7_75t_L g573 ( .A(n_26), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_27), .A2(n_277), .B1(n_507), .B2(n_508), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_28), .A2(n_34), .B1(n_329), .B2(n_496), .Y(n_495) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_29), .A2(n_83), .B1(n_308), .B2(n_313), .Y(n_317) );
INVx1_ASAP7_75t_L g821 ( .A(n_29), .Y(n_821) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_30), .A2(n_45), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_31), .A2(n_36), .B1(n_371), .B2(n_374), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_32), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_33), .A2(n_43), .B1(n_485), .B2(n_600), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_35), .A2(n_156), .B1(n_360), .B2(n_362), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_37), .A2(n_173), .B1(n_429), .B2(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_38), .A2(n_270), .B1(n_398), .B2(n_633), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_39), .A2(n_58), .B1(n_369), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_276), .B1(n_350), .B2(n_513), .Y(n_512) );
AOI222xp33_ASAP7_75t_L g748 ( .A1(n_41), .A2(n_126), .B1(n_202), .B2(n_366), .C1(n_369), .C2(n_593), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_42), .A2(n_244), .B1(n_487), .B2(n_489), .Y(n_486) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_44), .A2(n_86), .B1(n_308), .B2(n_309), .Y(n_315) );
INVx1_ASAP7_75t_L g822 ( .A(n_44), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_46), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_47), .A2(n_193), .B1(n_455), .B2(n_457), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_48), .A2(n_100), .B1(n_450), .B2(n_452), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_49), .A2(n_206), .B1(n_375), .B2(n_570), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_50), .A2(n_161), .B1(n_324), .B2(n_329), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_51), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_52), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_53), .A2(n_285), .B1(n_324), .B2(n_489), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_54), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_55), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_56), .Y(n_595) );
XOR2xp5_ASAP7_75t_L g300 ( .A(n_57), .B(n_301), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_59), .A2(n_248), .B1(n_611), .B2(n_746), .Y(n_745) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_60), .B(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_61), .A2(n_141), .B1(n_350), .B2(n_508), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_62), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_63), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_64), .A2(n_251), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_65), .A2(n_203), .B1(n_303), .B2(n_700), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_66), .A2(n_192), .B1(n_360), .B2(n_394), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_67), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g639 ( .A(n_68), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_69), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_70), .A2(n_130), .B1(n_393), .B2(n_448), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_71), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_72), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_73), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_74), .A2(n_157), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_75), .A2(n_265), .B1(n_372), .B2(n_389), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_76), .A2(n_84), .B1(n_336), .B2(n_341), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_77), .A2(n_246), .B1(n_666), .B2(n_668), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_78), .A2(n_220), .B1(n_446), .B2(n_457), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_79), .A2(n_148), .B1(n_702), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_80), .A2(n_214), .B1(n_349), .B2(n_375), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_81), .A2(n_125), .B1(n_489), .B2(n_496), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_82), .A2(n_146), .B1(n_318), .B2(n_746), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_85), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_87), .A2(n_182), .B1(n_446), .B2(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g293 ( .A(n_88), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_89), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_90), .A2(n_127), .B1(n_455), .B2(n_492), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_91), .A2(n_111), .B1(n_354), .B2(n_356), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_92), .A2(n_199), .B1(n_344), .B2(n_371), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_93), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_94), .A2(n_190), .B1(n_401), .B2(n_402), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_95), .A2(n_113), .B1(n_356), .B2(n_601), .Y(n_737) );
INVx1_ASAP7_75t_L g290 ( .A(n_96), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_97), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_98), .A2(n_232), .B1(n_389), .B2(n_796), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_101), .A2(n_242), .B1(n_318), .B2(n_629), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_102), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_103), .A2(n_235), .B1(n_354), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_104), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_105), .A2(n_218), .B1(n_606), .B2(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_106), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_107), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_109), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_112), .A2(n_134), .B1(n_350), .B2(n_389), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_114), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_115), .A2(n_219), .B1(n_600), .B2(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_116), .A2(n_240), .B1(n_401), .B2(n_632), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_117), .A2(n_778), .B1(n_805), .B2(n_806), .Y(n_777) );
INVx1_ASAP7_75t_L g805 ( .A(n_117), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_119), .A2(n_163), .B1(n_393), .B2(n_487), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_120), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_121), .A2(n_222), .B1(n_304), .B2(n_451), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_122), .B(n_834), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_123), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_124), .A2(n_267), .B1(n_372), .B2(n_374), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_128), .A2(n_159), .B1(n_459), .B2(n_705), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_129), .A2(n_208), .B1(n_432), .B2(n_654), .Y(n_653) );
XOR2x2_ASAP7_75t_L g411 ( .A(n_131), .B(n_412), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_132), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_135), .A2(n_223), .B1(n_457), .B2(n_707), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_136), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_138), .Y(n_555) );
INVx2_ASAP7_75t_L g294 ( .A(n_140), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_142), .A2(n_179), .B1(n_601), .B2(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_143), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_144), .A2(n_151), .B1(n_611), .B2(n_629), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_145), .A2(n_221), .B1(n_448), .B2(n_496), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_147), .A2(n_236), .B1(n_633), .B2(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g404 ( .A(n_149), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_150), .B(n_342), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_152), .B(n_336), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_153), .A2(n_278), .B1(n_329), .B2(n_450), .Y(n_602) );
AND2x6_ASAP7_75t_L g289 ( .A(n_154), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_154), .Y(n_815) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_155), .A2(n_231), .B1(n_308), .B2(n_309), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_158), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_160), .A2(n_262), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_162), .A2(n_169), .B1(n_700), .B2(n_879), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_164), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_166), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_167), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_168), .A2(n_258), .B1(n_570), .B2(n_572), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_170), .B(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_171), .A2(n_217), .B1(n_345), .B2(n_350), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_172), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_174), .A2(n_255), .B1(n_330), .B2(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_175), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_177), .B(n_386), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_178), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_180), .A2(n_284), .B1(n_336), .B2(n_341), .Y(n_636) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_181), .A2(n_250), .B1(n_308), .B2(n_313), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_183), .A2(n_281), .B1(n_318), .B2(n_360), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_185), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_186), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_187), .A2(n_227), .B1(n_360), .B2(n_362), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_188), .A2(n_211), .B1(n_432), .B2(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_189), .A2(n_263), .B1(n_494), .B2(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_SL g711 ( .A1(n_194), .A2(n_712), .B1(n_732), .B2(n_733), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_194), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_195), .Y(n_740) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_196), .B(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_197), .A2(n_210), .B1(n_428), .B2(n_478), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_198), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_200), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_201), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_204), .A2(n_273), .B1(n_318), .B2(n_702), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_205), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_207), .A2(n_280), .B1(n_398), .B2(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_209), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_212), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_213), .B(n_386), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_215), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_216), .B(n_342), .Y(n_511) );
OA22x2_ASAP7_75t_L g754 ( .A1(n_224), .A2(n_755), .B1(n_756), .B2(n_774), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_224), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_225), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_228), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_229), .A2(n_825), .B1(n_843), .B2(n_844), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_229), .Y(n_843) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_230), .A2(n_287), .B(n_295), .C(n_823), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_231), .B(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_233), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_234), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_237), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_238), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_239), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_241), .A2(n_245), .B1(n_393), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_243), .A2(n_283), .B1(n_364), .B2(n_460), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_249), .Y(n_531) );
INVx1_ASAP7_75t_L g818 ( .A(n_250), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_252), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_253), .B(n_432), .Y(n_431) );
OA22x2_ASAP7_75t_L g578 ( .A1(n_254), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_254), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_256), .B(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_257), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_259), .Y(n_683) );
INVx1_ASAP7_75t_L g852 ( .A(n_264), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_264), .A2(n_852), .B1(n_854), .B2(n_882), .Y(n_853) );
INVx1_ASAP7_75t_L g308 ( .A(n_266), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_268), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_269), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_271), .A2(n_275), .B1(n_303), .B2(n_318), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_274), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_279), .B(n_429), .Y(n_865) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_290), .Y(n_814) );
OA21x2_ASAP7_75t_L g850 ( .A1(n_291), .A2(n_813), .B(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_675), .B1(n_808), .B2(n_809), .C(n_810), .Y(n_295) );
INVx1_ASAP7_75t_L g808 ( .A(n_296), .Y(n_808) );
AOI22xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_619), .B1(n_620), .B2(n_674), .Y(n_296) );
INVx1_ASAP7_75t_L g674 ( .A(n_297), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_407), .B2(n_618), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_377), .B1(n_405), .B2(n_406), .Y(n_299) );
INVx1_ASAP7_75t_L g405 ( .A(n_300), .Y(n_405) );
NAND5xp2_ASAP7_75t_SL g301 ( .A(n_302), .B(n_323), .C(n_334), .D(n_352), .E(n_365), .Y(n_301) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
INVx6_ASAP7_75t_L g493 ( .A(n_304), .Y(n_493) );
BUFx3_ASAP7_75t_L g673 ( .A(n_304), .Y(n_673) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_314), .Y(n_304) );
AND2x2_ASAP7_75t_L g361 ( .A(n_305), .B(n_326), .Y(n_361) );
AND2x6_ASAP7_75t_L g364 ( .A(n_305), .B(n_339), .Y(n_364) );
AND2x6_ASAP7_75t_L g367 ( .A(n_305), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_311), .Y(n_305) );
AND2x2_ASAP7_75t_L g328 ( .A(n_306), .B(n_312), .Y(n_328) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g321 ( .A(n_307), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_307), .B(n_312), .Y(n_333) );
AND2x2_ASAP7_75t_L g348 ( .A(n_307), .B(n_317), .Y(n_348) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_310), .Y(n_313) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g322 ( .A(n_312), .Y(n_322) );
INVx1_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
AND2x2_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
AND2x6_ASAP7_75t_L g342 ( .A(n_314), .B(n_328), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_314), .B(n_328), .Y(n_424) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
INVx1_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
OR2x2_ASAP7_75t_L g340 ( .A(n_315), .B(n_316), .Y(n_340) );
AND2x2_ASAP7_75t_L g368 ( .A(n_315), .B(n_317), .Y(n_368) );
AND2x2_ASAP7_75t_L g326 ( .A(n_316), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx5_ASAP7_75t_L g399 ( .A(n_319), .Y(n_399) );
INVx4_ASAP7_75t_L g451 ( .A(n_319), .Y(n_451) );
INVx2_ASAP7_75t_L g494 ( .A(n_319), .Y(n_494) );
BUFx3_ASAP7_75t_L g667 ( .A(n_319), .Y(n_667) );
INVx8_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g355 ( .A(n_321), .B(n_326), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_321), .B(n_326), .Y(n_558) );
INVx1_ASAP7_75t_L g376 ( .A(n_322), .Y(n_376) );
BUFx2_ASAP7_75t_L g457 ( .A(n_324), .Y(n_457) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_325), .Y(n_401) );
BUFx3_ASAP7_75t_L g496 ( .A(n_325), .Y(n_496) );
BUFx3_ASAP7_75t_L g611 ( .A(n_325), .Y(n_611) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x4_ASAP7_75t_L g357 ( .A(n_326), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g346 ( .A(n_327), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g403 ( .A(n_327), .Y(n_403) );
AND2x4_ASAP7_75t_L g338 ( .A(n_328), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g419 ( .A(n_328), .Y(n_419) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g629 ( .A(n_330), .Y(n_629) );
BUFx2_ASAP7_75t_L g881 ( .A(n_330), .Y(n_881) );
INVx6_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g452 ( .A(n_331), .Y(n_452) );
INVx1_ASAP7_75t_SL g668 ( .A(n_331), .Y(n_668) );
INVx1_ASAP7_75t_SL g702 ( .A(n_331), .Y(n_702) );
OR2x6_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g351 ( .A(n_332), .Y(n_351) );
INVx1_ASAP7_75t_L g358 ( .A(n_333), .Y(n_358) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_335), .B(n_343), .Y(n_334) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g386 ( .A(n_337), .Y(n_386) );
INVx5_ASAP7_75t_L g535 ( .A(n_337), .Y(n_535) );
INVx2_ASAP7_75t_L g568 ( .A(n_337), .Y(n_568) );
INVx4_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g418 ( .A(n_340), .B(n_419), .Y(n_418) );
BUFx4f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g566 ( .A(n_342), .Y(n_566) );
INVx1_ASAP7_75t_SL g766 ( .A(n_342), .Y(n_766) );
BUFx2_ASAP7_75t_L g834 ( .A(n_342), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_344), .Y(n_798) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_345), .Y(n_432) );
BUFx2_ASAP7_75t_L g478 ( .A(n_345), .Y(n_478) );
BUFx4f_ASAP7_75t_SL g513 ( .A(n_345), .Y(n_513) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
AND2x4_ASAP7_75t_L g350 ( .A(n_348), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g372 ( .A(n_348), .B(n_373), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_348), .B(n_403), .Y(n_436) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g571 ( .A(n_350), .Y(n_571) );
BUFx2_ASAP7_75t_L g796 ( .A(n_350), .Y(n_796) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_359), .Y(n_352) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
BUFx3_ASAP7_75t_L g460 ( .A(n_355), .Y(n_460) );
BUFx3_ASAP7_75t_L g875 ( .A(n_355), .Y(n_875) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_357), .Y(n_448) );
BUFx3_ASAP7_75t_L g489 ( .A(n_357), .Y(n_489) );
INVx1_ASAP7_75t_L g613 ( .A(n_357), .Y(n_613) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_357), .Y(n_705) );
AND2x2_ASAP7_75t_L g402 ( .A(n_358), .B(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g447 ( .A(n_360), .Y(n_447) );
BUFx3_ASAP7_75t_L g700 ( .A(n_360), .Y(n_700) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g488 ( .A(n_361), .Y(n_488) );
BUFx2_ASAP7_75t_SL g632 ( .A(n_361), .Y(n_632) );
INVx5_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g485 ( .A(n_363), .Y(n_485) );
INVx2_ASAP7_75t_SL g516 ( .A(n_363), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_363), .A2(n_493), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g601 ( .A(n_363), .Y(n_601) );
INVx11_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx11_ASAP7_75t_L g456 ( .A(n_364), .Y(n_456) );
INVx2_ASAP7_75t_SL g800 ( .A(n_366), .Y(n_800) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g382 ( .A(n_367), .Y(n_382) );
BUFx3_ASAP7_75t_L g473 ( .A(n_367), .Y(n_473) );
INVx4_ASAP7_75t_L g505 ( .A(n_367), .Y(n_505) );
INVx2_ASAP7_75t_SL g689 ( .A(n_367), .Y(n_689) );
INVx2_ASAP7_75t_L g759 ( .A(n_367), .Y(n_759) );
AND2x4_ASAP7_75t_L g375 ( .A(n_368), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g441 ( .A(n_368), .Y(n_441) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx4f_ASAP7_75t_SL g563 ( .A(n_371), .Y(n_563) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_372), .Y(n_507) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_375), .Y(n_508) );
BUFx2_ASAP7_75t_SL g572 ( .A(n_375), .Y(n_572) );
BUFx2_ASAP7_75t_SL g830 ( .A(n_375), .Y(n_830) );
INVx1_ASAP7_75t_L g442 ( .A(n_376), .Y(n_442) );
INVx2_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
XOR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_404), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_379), .B(n_390), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_384), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_382), .A2(n_426), .B1(n_427), .B2(n_430), .C(n_431), .Y(n_425) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_382), .A2(n_652), .B(n_653), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .C(n_388), .Y(n_384) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_389), .Y(n_687) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_396), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx4_ASAP7_75t_L g664 ( .A(n_401), .Y(n_664) );
INVx3_ASAP7_75t_L g643 ( .A(n_406), .Y(n_643) );
INVx1_ASAP7_75t_L g618 ( .A(n_407), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_521), .B1(n_615), .B2(n_617), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g616 ( .A(n_410), .Y(n_616) );
OA22x2_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_461), .B1(n_519), .B2(n_520), .Y(n_410) );
INVx2_ASAP7_75t_L g519 ( .A(n_411), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_443), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_425), .C(n_433), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_420), .B2(n_421), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_418), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_418), .Y(n_586) );
BUFx3_ASAP7_75t_L g649 ( .A(n_418), .Y(n_649) );
OAI221xp5_ASAP7_75t_SL g792 ( .A1(n_421), .A2(n_586), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g588 ( .A(n_423), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g682 ( .A1(n_423), .A2(n_586), .B1(n_683), .B2(n_684), .Y(n_682) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g803 ( .A(n_429), .Y(n_803) );
BUFx2_ASAP7_75t_L g593 ( .A(n_432), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_433) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx4_ASAP7_75t_L g481 ( .A(n_436), .Y(n_481) );
OAI22xp33_ASAP7_75t_SL g594 ( .A1(n_436), .A2(n_438), .B1(n_595), .B2(n_596), .Y(n_594) );
BUFx3_ASAP7_75t_L g694 ( .A(n_436), .Y(n_694) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_438), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g659 ( .A(n_439), .Y(n_659) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_440), .A2(n_657), .B1(n_722), .B2(n_723), .Y(n_721) );
BUFx2_ASAP7_75t_L g869 ( .A(n_440), .Y(n_869) );
OR2x6_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_449), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_447), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_553) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g549 ( .A(n_451), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_458), .Y(n_453) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g633 ( .A(n_456), .Y(n_633) );
INVx3_ASAP7_75t_L g728 ( .A(n_456), .Y(n_728) );
BUFx4f_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g708 ( .A(n_460), .Y(n_708) );
INVx2_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_497), .Y(n_461) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_482), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_470), .C(n_475), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g717 ( .A(n_469), .Y(n_717) );
INVx1_ASAP7_75t_SL g859 ( .A(n_469), .Y(n_859) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_474), .Y(n_470) );
OAI21xp33_ASAP7_75t_SL g590 ( .A1(n_472), .A2(n_591), .B(n_592), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_472), .A2(n_639), .B(n_640), .Y(n_638) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_SL g657 ( .A(n_481), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_490), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g600 ( .A(n_488), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
INVx3_ASAP7_75t_L g746 ( .A(n_493), .Y(n_746) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_494), .Y(n_786) );
BUFx2_ASAP7_75t_L g789 ( .A(n_496), .Y(n_789) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_518), .Y(n_497) );
NAND3x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .C(n_514), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_506), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_505), .A2(n_531), .B(n_532), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_505), .A2(n_561), .B(n_562), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g827 ( .A1(n_505), .A2(n_828), .B(n_829), .Y(n_827) );
BUFx2_ASAP7_75t_L g861 ( .A(n_505), .Y(n_861) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_507), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .C(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g863 ( .A(n_513), .Y(n_863) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_575), .B1(n_576), .B2(n_614), .Y(n_521) );
INVx1_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
OA22x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B1(n_542), .B2(n_574), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_523), .A2(n_524), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
XOR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_541), .Y(n_524) );
NAND3x1_ASAP7_75t_SL g525 ( .A(n_526), .B(n_529), .C(n_538), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_533), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .C(n_537), .Y(n_533) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_535), .Y(n_742) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g574 ( .A(n_542), .Y(n_574) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_573), .Y(n_542) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_544), .B(n_559), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .C(n_553), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_556), .A2(n_604), .B1(n_605), .B2(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g781 ( .A(n_557), .Y(n_781) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .C(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_597), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .C(n_594), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_586), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_586), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_588), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .C(n_608), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_611), .Y(n_879) );
INVx1_ASAP7_75t_L g671 ( .A(n_613), .Y(n_671) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AO22x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_641), .B2(n_642), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NOR4xp75_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .C(n_635), .D(n_638), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_631), .B(n_634), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
XNOR2x1_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_660), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .C(n_655), .Y(n_646) );
INVx1_ASAP7_75t_L g691 ( .A(n_654), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_657), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_669), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx4_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g809 ( .A(n_675), .Y(n_809) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_753), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_709), .B1(n_710), .B2(n_752), .Y(n_677) );
INVx2_ASAP7_75t_L g752 ( .A(n_678), .Y(n_752) );
XNOR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_697), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .C(n_693), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_689), .B2(n_690), .C1(n_691), .C2(n_692), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_689), .A2(n_719), .B(n_720), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_703), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g783 ( .A(n_705), .Y(n_783) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AO22x1_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_734), .B1(n_750), .B2(n_751), .Y(n_710) );
INVx1_ASAP7_75t_L g750 ( .A(n_711), .Y(n_750) );
INVx2_ASAP7_75t_L g732 ( .A(n_712), .Y(n_732) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_724), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .C(n_721), .Y(n_713) );
OA211x2_ASAP7_75t_L g739 ( .A1(n_717), .A2(n_740), .B(n_741), .C(n_743), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_729), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g751 ( .A(n_734), .Y(n_751) );
XOR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_749), .Y(n_734) );
NAND4xp75_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .C(n_744), .D(n_748), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_775), .B1(n_776), .B2(n_807), .Y(n_753) );
INVx1_ASAP7_75t_L g807 ( .A(n_754), .Y(n_807) );
INVx2_ASAP7_75t_L g774 ( .A(n_756), .Y(n_774) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_767), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_762), .Y(n_757) );
OAI21xp5_ASAP7_75t_SL g758 ( .A1(n_759), .A2(n_760), .B(n_761), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g806 ( .A(n_778), .Y(n_806) );
AND2x2_ASAP7_75t_SL g778 ( .A(n_779), .B(n_791), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_787), .Y(n_779) );
OAI221xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_782), .B1(n_783), .B2(n_784), .C(n_785), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
NOR2xp33_ASAP7_75t_SL g791 ( .A(n_792), .B(n_797), .Y(n_791) );
OAI222xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_800), .B2(n_801), .C1(n_802), .C2(n_804), .Y(n_797) );
INVxp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
NOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_816), .Y(n_811) );
OR2x2_ASAP7_75t_SL g885 ( .A(n_812), .B(n_817), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_813), .Y(n_846) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_814), .B(n_849), .Y(n_851) );
CKINVDCx16_ASAP7_75t_R g849 ( .A(n_815), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
OAI322xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_845), .A3(n_847), .B1(n_850), .B2(n_852), .C1(n_853), .C2(n_883), .Y(n_823) );
INVx1_ASAP7_75t_L g844 ( .A(n_825), .Y(n_844) );
AND2x4_ASAP7_75t_L g825 ( .A(n_826), .B(n_836), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .Y(n_826) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .C(n_835), .Y(n_831) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_840), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g882 ( .A(n_854), .Y(n_882) );
AND2x2_ASAP7_75t_SL g854 ( .A(n_855), .B(n_870), .Y(n_854) );
NOR3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .C(n_866), .Y(n_855) );
OAI221xp5_ASAP7_75t_SL g860 ( .A1(n_861), .A2(n_862), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_877), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_876), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_885), .Y(n_884) );
endmodule