module fake_netlist_1_10068_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
XNOR2xp5_ASAP7_75t_L g13 ( .A(n_0), .B(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
NOR2xp33_ASAP7_75t_SL g15 ( .A(n_1), .B(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_11), .Y(n_16) );
NOR2xp67_ASAP7_75t_L g17 ( .A(n_2), .B(n_10), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_5), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_14), .B(n_3), .C(n_4), .Y(n_20) );
BUFx4f_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B1(n_13), .B2(n_18), .Y(n_22) );
NOR2xp33_ASAP7_75t_R g23 ( .A(n_22), .B(n_21), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OAI221xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_13), .B1(n_18), .B2(n_15), .C(n_17), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_15), .B1(n_16), .B2(n_17), .C(n_7), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI22xp33_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_25), .B1(n_5), .B2(n_6), .Y(n_28) );
AOI222xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_4), .B1(n_6), .B2(n_8), .C1(n_9), .C2(n_12), .Y(n_29) );
endmodule