module fake_jpeg_24717_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_21),
.B1(n_35),
.B2(n_45),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_20),
.B1(n_30),
.B2(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_35),
.B1(n_22),
.B2(n_19),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_32),
.B1(n_33),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_71),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_29),
.B1(n_22),
.B2(n_32),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_44),
.B1(n_31),
.B2(n_19),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_29),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_45),
.B1(n_38),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_93),
.B1(n_107),
.B2(n_52),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_45),
.B1(n_19),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_79),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_32),
.B1(n_44),
.B2(n_39),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_44),
.B(n_32),
.C(n_42),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_34),
.B1(n_17),
.B2(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_100),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_24),
.B1(n_33),
.B2(n_20),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_20),
.B1(n_30),
.B2(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_18),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_1),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_18),
.B1(n_28),
.B2(n_26),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_0),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_63),
.B1(n_69),
.B2(n_62),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_117),
.B(n_102),
.Y(n_145)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_116),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_1),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_105),
.B1(n_103),
.B2(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_52),
.B1(n_18),
.B2(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_94),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_26),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_77),
.Y(n_140)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_26),
.B1(n_55),
.B2(n_47),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_55),
.B1(n_47),
.B2(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_142),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_153),
.B1(n_165),
.B2(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_78),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_74),
.B(n_84),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_150),
.B(n_152),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_156),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_170),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_105),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_87),
.B1(n_73),
.B2(n_90),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_90),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_157),
.B(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_13),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_95),
.B(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_118),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_96),
.B1(n_79),
.B2(n_104),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_10),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_76),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_3),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_3),
.B(n_4),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_3),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_184),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_119),
.B(n_127),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_183),
.B(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_181),
.B1(n_196),
.B2(n_183),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_127),
.C(n_128),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_189),
.C(n_145),
.Y(n_209)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_113),
.B1(n_121),
.B2(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_114),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_113),
.B(n_128),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_114),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_135),
.C(n_109),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_138),
.B(n_109),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_200),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_139),
.A2(n_109),
.B1(n_121),
.B2(n_76),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_199),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_150),
.B(n_3),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_140),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_211),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_151),
.B(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_213),
.B(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_153),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_152),
.B(n_143),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_141),
.B1(n_163),
.B2(n_159),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_218),
.B1(n_181),
.B2(n_180),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_177),
.B(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_198),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_226),
.Y(n_230)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_144),
.C(n_164),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_221),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_171),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_144),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_167),
.B(n_162),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_139),
.B(n_160),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_191),
.B(n_179),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_231),
.A2(n_241),
.B1(n_249),
.B2(n_211),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_233),
.A2(n_227),
.B(n_220),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_199),
.B1(n_185),
.B2(n_180),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_240),
.B1(n_242),
.B2(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_185),
.B1(n_175),
.B2(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_175),
.B1(n_193),
.B2(n_177),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_205),
.B1(n_211),
.B2(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_172),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_204),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_194),
.B1(n_187),
.B2(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_224),
.A2(n_190),
.B1(n_189),
.B2(n_160),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_258),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_229),
.B(n_222),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_255),
.B1(n_266),
.B2(n_237),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_262),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_231),
.B1(n_243),
.B2(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_209),
.C(n_217),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_238),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_228),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_226),
.C(n_213),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_206),
.C(n_208),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_227),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_244),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_220),
.B(n_190),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_233),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_242),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_275),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_281),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_274),
.B(n_277),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_254),
.C(n_230),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_280),
.B1(n_253),
.B2(n_261),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_234),
.B1(n_239),
.B2(n_250),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_279),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_262),
.B(n_250),
.Y(n_284)
);

AOI21x1_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_288),
.B(n_9),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_273),
.B1(n_280),
.B2(n_271),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_268),
.B1(n_247),
.B2(n_259),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_256),
.B(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_293),
.C(n_14),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_195),
.C(n_76),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_12),
.B(n_15),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_9),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_12),
.B(n_15),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_284),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_281),
.B1(n_276),
.B2(n_13),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_8),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_16),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_304),
.B(n_285),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_302),
.CI(n_296),
.CON(n_311),
.SN(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_310),
.A3(n_14),
.B1(n_16),
.B2(n_6),
.C1(n_4),
.C2(n_5),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_304),
.B(n_293),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_4),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_290),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_312),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_306),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.C(n_313),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_6),
.Y(n_320)
);


endmodule