module fake_netlist_6_2370_n_2459 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2459);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2459;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_383;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_437;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_2127;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_374;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_330;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_1456;
wire n_394;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_115),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_68),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_96),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_162),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_118),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_132),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_102),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_59),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_160),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_230),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_127),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_129),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_107),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_215),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_24),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_54),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_130),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_15),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_49),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_163),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_173),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_222),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_176),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_186),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_117),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_226),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_44),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_17),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_63),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_72),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_90),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_97),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_90),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_111),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_94),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_58),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_192),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_139),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_71),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_82),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_185),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_73),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_102),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_193),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_142),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_131),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_201),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_7),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_60),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_124),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_146),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_190),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_145),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_33),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_198),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_137),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_39),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_61),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_197),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_134),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_184),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_189),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_24),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_140),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_19),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_88),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_34),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_107),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_108),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_76),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_151),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_88),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_39),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_85),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_205),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_208),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_180),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_156),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_174),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_56),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_29),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_65),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_18),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_200),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_191),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_20),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_52),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_25),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_113),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_85),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_42),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_65),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_152),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_161),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_30),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_43),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_77),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_19),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_168),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_170),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_188),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_49),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_12),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_70),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_48),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_128),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_68),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_23),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_78),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_159),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_64),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_164),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_175),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_126),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_116),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_71),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_8),
.Y(n_384)
);

BUFx2_ASAP7_75t_SL g385 ( 
.A(n_29),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_91),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_155),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_12),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_228),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_50),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_112),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_147),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_3),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_109),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_224),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_27),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_54),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_231),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_41),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_16),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_4),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_76),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_227),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_42),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_26),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_70),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_86),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_167),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_135),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_218),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_21),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_80),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_179),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_121),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_53),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_86),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_7),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_105),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_45),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_22),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_63),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_77),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_223),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_84),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_84),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_27),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_51),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_183),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_136),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_110),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_199),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_149),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_58),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_6),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_105),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_10),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_67),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_80),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_9),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_92),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_141),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_69),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_100),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_5),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_55),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_104),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_203),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_207),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_98),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_37),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_15),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_178),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_119),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_57),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_96),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_270),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_351),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_246),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_270),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_270),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_241),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_236),
.Y(n_464)
);

BUFx2_ASAP7_75t_SL g465 ( 
.A(n_415),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_270),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_270),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_270),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_439),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_363),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_259),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_243),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_245),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_247),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_275),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_350),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_252),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_442),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_448),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_347),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_270),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_270),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_316),
.B(n_415),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_270),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_369),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_253),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_255),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_240),
.B(n_0),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_260),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_314),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_314),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_314),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_314),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_408),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_261),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_262),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_314),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_269),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_314),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_314),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_272),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_274),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_314),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_276),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_277),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_314),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_316),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_338),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_345),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_338),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_338),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_279),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_338),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_233),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_369),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_289),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_347),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_295),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_237),
.B(n_0),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_234),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_302),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_338),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_338),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_309),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_345),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_310),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_353),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_353),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_353),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_353),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_311),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_320),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_321),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_353),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_353),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_372),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_323),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_372),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_328),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_386),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_372),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_234),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_372),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_334),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_340),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_372),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_344),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_372),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_322),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_344),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_390),
.B(n_2),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_344),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_384),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_324),
.B(n_2),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_384),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_384),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_386),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_341),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_342),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_343),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_388),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_355),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_234),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_384),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_390),
.B(n_5),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_359),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_384),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_360),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_324),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_365),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_324),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_248),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_366),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_449),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_367),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_464),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_462),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_520),
.B(n_264),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_550),
.B(n_322),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_463),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_472),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_473),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_477),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_486),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_510),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_550),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_483),
.B(n_368),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_470),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_510),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_543),
.B(n_264),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_487),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_480),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_511),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_511),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_373),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_550),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_460),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_459),
.B(n_377),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_460),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_489),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_548),
.A2(n_553),
.B(n_551),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_495),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_513),
.B(n_264),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_474),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_523),
.B(n_326),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_523),
.B(n_326),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_524),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_528),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_475),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_461),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_496),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_498),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_461),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_485),
.A2(n_266),
.B1(n_286),
.B2(n_239),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_528),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_491),
.B(n_322),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_501),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_326),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_469),
.B(n_280),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_531),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_491),
.A2(n_466),
.B(n_457),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_531),
.B(n_370),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_465),
.B(n_379),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_535),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_457),
.A2(n_449),
.B(n_244),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_502),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_535),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_469),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_504),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_476),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_466),
.A2(n_244),
.B(n_237),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_536),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_536),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_548),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_R g657 ( 
.A(n_505),
.B(n_380),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_478),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_539),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_542),
.B(n_370),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_512),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_479),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_515),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_544),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_465),
.B(n_381),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_516),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_548),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_544),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_547),
.Y(n_670)
);

NAND2x1_ASAP7_75t_L g671 ( 
.A(n_547),
.B(n_322),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_527),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_549),
.B(n_258),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_549),
.B(n_370),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_532),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_551),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_554),
.B(n_387),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_638),
.B(n_257),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_641),
.B(n_573),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_640),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_514),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_322),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_642),
.B(n_533),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_588),
.B(n_485),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_641),
.B(n_573),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_584),
.B(n_322),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_640),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_641),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_R g690 ( 
.A(n_664),
.B(n_494),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_613),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_613),
.Y(n_692)
);

INVx6_ASAP7_75t_L g693 ( 
.A(n_619),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_605),
.B(n_534),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_657),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_650),
.B(n_281),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_666),
.B(n_538),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_660),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_588),
.B(n_558),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_605),
.B(n_540),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_596),
.B(n_545),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_666),
.B(n_546),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_660),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_596),
.B(n_577),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_660),
.B(n_575),
.Y(n_706)
);

BUFx4f_ASAP7_75t_L g707 ( 
.A(n_673),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_613),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_585),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_613),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_619),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_674),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_584),
.B(n_599),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_677),
.B(n_563),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_599),
.B(n_507),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_673),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_607),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_581),
.B(n_578),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_608),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_677),
.B(n_580),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_599),
.B(n_554),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_597),
.B(n_558),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_589),
.B(n_518),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_674),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_590),
.B(n_521),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_609),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_674),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_591),
.B(n_522),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_609),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_619),
.B(n_575),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_607),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_657),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_619),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_619),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_607),
.Y(n_737)
);

INVx4_ASAP7_75t_SL g738 ( 
.A(n_632),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_583),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_582),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_673),
.B(n_577),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_615),
.B(n_576),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_583),
.Y(n_743)
);

AND2x6_ASAP7_75t_L g744 ( 
.A(n_673),
.B(n_258),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_587),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_609),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_629),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_629),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_638),
.B(n_471),
.C(n_458),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_592),
.B(n_525),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_594),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_609),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_615),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_629),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_627),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_609),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_615),
.A2(n_519),
.B1(n_555),
.B2(n_552),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_608),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_618),
.B(n_637),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_618),
.B(n_556),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_609),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_618),
.B(n_556),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_594),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_598),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_610),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_637),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_664),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_637),
.B(n_576),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_650),
.A2(n_555),
.B1(n_569),
.B2(n_552),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_644),
.B(n_268),
.Y(n_773)
);

CKINVDCx8_ASAP7_75t_R g774 ( 
.A(n_647),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_627),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_627),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_627),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_598),
.B(n_557),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_610),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_602),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_646),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_597),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_610),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_610),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_646),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_602),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_603),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_601),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_600),
.B(n_559),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_611),
.B(n_268),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_603),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_616),
.B(n_620),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_616),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_610),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_620),
.B(n_557),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_647),
.B(n_541),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_610),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_614),
.B(n_625),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_644),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_626),
.B(n_278),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_636),
.A2(n_561),
.B1(n_570),
.B2(n_565),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_610),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_645),
.B(n_572),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_621),
.B(n_622),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_622),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_644),
.B(n_650),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_624),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_560),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_631),
.B(n_560),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_648),
.B(n_574),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_633),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_662),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_624),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_624),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_278),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_667),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_612),
.B(n_257),
.Y(n_821)
);

INVxp33_ASAP7_75t_L g822 ( 
.A(n_628),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_624),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_634),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_634),
.B(n_567),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_632),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_671),
.B(n_305),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_624),
.B(n_293),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_612),
.B(n_385),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_624),
.B(n_293),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_635),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_651),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_617),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_635),
.B(n_567),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_639),
.B(n_571),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_639),
.B(n_304),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_623),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_649),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_651),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_761),
.B(n_304),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_691),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_681),
.B(n_672),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_691),
.B(n_585),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_761),
.B(n_675),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_761),
.B(n_630),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_755),
.B(n_630),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_720),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_690),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_702),
.B(n_562),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_770),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_683),
.B(n_564),
.Y(n_851)
);

AND2x2_ASAP7_75t_SL g852 ( 
.A(n_772),
.B(n_315),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_691),
.B(n_708),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_630),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_769),
.B(n_630),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_769),
.B(n_630),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_698),
.B(n_630),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_703),
.B(n_471),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_714),
.B(n_630),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_716),
.B(n_396),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_SL g861 ( 
.A(n_822),
.B(n_298),
.C(n_291),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_716),
.B(n_404),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_714),
.B(n_643),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_770),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_712),
.B(n_315),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_694),
.B(n_658),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_735),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_736),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_720),
.B(n_410),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_820),
.Y(n_870)
);

BUFx8_ASAP7_75t_L g871 ( 
.A(n_805),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_773),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_732),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_760),
.B(n_411),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_773),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_685),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_709),
.B(n_710),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_760),
.B(n_414),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_691),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_696),
.B(n_429),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_689),
.B(n_509),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_692),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_714),
.B(n_652),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_734),
.B(n_432),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_714),
.A2(n_389),
.B1(n_399),
.B2(n_382),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_691),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_SL g887 ( 
.A(n_678),
.B(n_280),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_701),
.B(n_280),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_708),
.B(n_653),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_732),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_692),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_699),
.A2(n_628),
.B1(n_569),
.B2(n_331),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_695),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_695),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_712),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_715),
.B(n_663),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_708),
.B(n_653),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_L g898 ( 
.A(n_759),
.B(n_389),
.C(n_382),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_708),
.B(n_654),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_708),
.B(n_654),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_732),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_693),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_833),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_721),
.B(n_655),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_697),
.B(n_585),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_680),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_722),
.B(n_655),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_711),
.B(n_659),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_684),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_688),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_705),
.B(n_280),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_711),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_697),
.B(n_585),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_711),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_693),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_693),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_742),
.B(n_659),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_693),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_773),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_742),
.B(n_661),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_742),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_704),
.A2(n_713),
.B1(n_729),
.B2(n_726),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_771),
.B(n_661),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_833),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_705),
.B(n_306),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_771),
.A2(n_399),
.B1(n_424),
.B2(n_409),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_665),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_679),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_679),
.B(n_509),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_808),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_709),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_679),
.B(n_665),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_686),
.B(n_669),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_686),
.B(n_669),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_686),
.B(n_706),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_790),
.B(n_801),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_706),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_741),
.A2(n_488),
.B(n_444),
.C(n_571),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_706),
.B(n_670),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_819),
.B(n_836),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_820),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_718),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_739),
.B(n_670),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_781),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_743),
.B(n_586),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_819),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_744),
.A2(n_409),
.B1(n_430),
.B2(n_424),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_745),
.B(n_586),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_750),
.B(n_586),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_753),
.B(n_586),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_819),
.B(n_430),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_685),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_678),
.A2(n_332),
.B1(n_398),
.B2(n_333),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_678),
.A2(n_418),
.B1(n_446),
.B2(n_433),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_719),
.B(n_283),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_766),
.B(n_606),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_836),
.B(n_678),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_767),
.B(n_606),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_744),
.A2(n_433),
.B1(n_454),
.B2(n_453),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_718),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_808),
.A2(n_671),
.B(n_553),
.C(n_568),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_836),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_781),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_805),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_780),
.B(n_606),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_790),
.B(n_306),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_801),
.B(n_306),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_733),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_786),
.B(n_606),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_787),
.B(n_791),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_796),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_838),
.Y(n_972)
);

OAI221xp5_ASAP7_75t_L g973 ( 
.A1(n_751),
.A2(n_488),
.B1(n_444),
.B2(n_319),
.C(n_301),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_758),
.A2(n_794),
.B(n_717),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_839),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_741),
.B(n_306),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_733),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_793),
.B(n_798),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_SL g979 ( 
.A1(n_762),
.A2(n_454),
.B1(n_453),
.B2(n_256),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_815),
.B(n_312),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_737),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_744),
.A2(n_385),
.B1(n_632),
.B2(n_468),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_807),
.B(n_593),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_814),
.B(n_593),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_824),
.B(n_593),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_707),
.A2(n_723),
.B(n_717),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_831),
.B(n_595),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_737),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_764),
.B(n_595),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_792),
.B(n_595),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_806),
.B(n_604),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_800),
.B(n_526),
.Y(n_993)
);

BUFx6f_ASAP7_75t_SL g994 ( 
.A(n_820),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_782),
.B(n_376),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_815),
.B(n_312),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_700),
.B(n_235),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_682),
.B(n_604),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_682),
.B(n_604),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_682),
.B(n_632),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_839),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_682),
.B(n_632),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_707),
.A2(n_468),
.B1(n_481),
.B2(n_467),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_707),
.B(n_312),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_682),
.B(n_632),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_700),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_747),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_682),
.B(n_632),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_687),
.A2(n_744),
.B1(n_808),
.B2(n_822),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_785),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_687),
.B(n_632),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_957),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_870),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_882),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_993),
.B(n_821),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_858),
.B(n_799),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_882),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_903),
.B(n_838),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_SL g1019 ( 
.A(n_955),
.B(n_796),
.C(n_774),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_964),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_904),
.B(n_993),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_861),
.B(n_972),
.C(n_924),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_852),
.B(n_687),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_852),
.B(n_687),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_881),
.B(n_821),
.Y(n_1025)
);

AND3x1_ASAP7_75t_SL g1026 ( 
.A(n_973),
.B(n_256),
.C(n_240),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_995),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_941),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_919),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_891),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_879),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_L g1032 ( 
.A(n_844),
.B(n_799),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_919),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_903),
.B(n_924),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_879),
.Y(n_1035)
);

OR2x6_ASAP7_75t_SL g1036 ( 
.A(n_847),
.B(n_802),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_891),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_879),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_851),
.B(n_725),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_849),
.B(n_727),
.Y(n_1040)
);

CKINVDCx8_ASAP7_75t_R g1041 ( 
.A(n_847),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_941),
.B(n_730),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_944),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_886),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_971),
.B(n_724),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_852),
.B(n_687),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_842),
.B(n_752),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_893),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_944),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_963),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_886),
.B(n_789),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_963),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_893),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_871),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_848),
.B(n_804),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_894),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_898),
.A2(n_744),
.B1(n_687),
.B2(n_723),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_871),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_894),
.B(n_841),
.Y(n_1059)
);

BUFx4f_ASAP7_75t_L g1060 ( 
.A(n_957),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_850),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_972),
.Y(n_1062)
);

AND2x6_ASAP7_75t_SL g1063 ( 
.A(n_896),
.B(n_813),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_886),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_871),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_914),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_870),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_912),
.B(n_940),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_SL g1069 ( 
.A(n_929),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_898),
.A2(n_744),
.B1(n_717),
.B2(n_723),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_881),
.B(n_821),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_1006),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_895),
.B(n_821),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_887),
.B(n_774),
.Y(n_1074)
);

INVx3_ASAP7_75t_SL g1075 ( 
.A(n_1004),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_975),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_887),
.B(n_724),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_895),
.B(n_829),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_921),
.B(n_829),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_864),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_975),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_870),
.B(n_837),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_936),
.A2(n_829),
.B1(n_788),
.B2(n_827),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_914),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_876),
.B(n_740),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_871),
.Y(n_1086)
);

INVx6_ASAP7_75t_L g1087 ( 
.A(n_930),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_872),
.A2(n_827),
.B1(n_826),
.B2(n_829),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_942),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_853),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_940),
.B(n_728),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_952),
.B(n_526),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_994),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_997),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_929),
.B(n_738),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_946),
.B(n_728),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_873),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_853),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1001),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_946),
.B(n_728),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_962),
.B(n_748),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_840),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1001),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_930),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_942),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1010),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_921),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_931),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_960),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_962),
.B(n_826),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_928),
.B(n_738),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_872),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1010),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_960),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_930),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_994),
.B(n_866),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_867),
.B(n_748),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_867),
.B(n_748),
.Y(n_1118)
);

OAI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_954),
.A2(n_826),
.B1(n_428),
.B2(n_440),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_875),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_937),
.B(n_738),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_968),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_840),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_875),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_968),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_994),
.B(n_754),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_868),
.B(n_754),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_868),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_979),
.A2(n_795),
.B(n_811),
.C(n_778),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_937),
.B(n_738),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_930),
.B(n_797),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_977),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_977),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_930),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_935),
.B(n_754),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_930),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_902),
.B(n_763),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_860),
.Y(n_1138)
);

INVx8_ASAP7_75t_L g1139 ( 
.A(n_840),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_902),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_922),
.B(n_763),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_873),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_981),
.Y(n_1143)
);

INVxp33_ASAP7_75t_SL g1144 ( 
.A(n_953),
.Y(n_1144)
);

CKINVDCx16_ASAP7_75t_R g1145 ( 
.A(n_953),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_889),
.A2(n_803),
.B(n_763),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_859),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_981),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_988),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_922),
.B(n_803),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_988),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_991),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_890),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_991),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_862),
.B(n_427),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_954),
.B(n_709),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_869),
.B(n_797),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_R g1158 ( 
.A(n_890),
.B(n_803),
.Y(n_1158)
);

AND3x1_ASAP7_75t_L g1159 ( 
.A(n_892),
.B(n_273),
.C(n_267),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_970),
.B(n_810),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_840),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1007),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1007),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_978),
.B(n_810),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_915),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_885),
.A2(n_951),
.B1(n_865),
.B2(n_901),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_910),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_880),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_SL g1169 ( 
.A(n_966),
.B(n_242),
.C(n_238),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_901),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_874),
.B(n_812),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_865),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_967),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_906),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_910),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_906),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_865),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_878),
.B(n_825),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_884),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_909),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_SL g1181 ( 
.A1(n_892),
.A2(n_249),
.B1(n_251),
.B2(n_250),
.Y(n_1181)
);

CKINVDCx6p67_ASAP7_75t_R g1182 ( 
.A(n_980),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_931),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_996),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_888),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1009),
.B(n_709),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1009),
.A2(n_428),
.B1(n_440),
.B2(n_427),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_865),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_915),
.A2(n_810),
.B1(n_823),
.B2(n_818),
.Y(n_1189)
);

INVx8_ASAP7_75t_L g1190 ( 
.A(n_951),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_931),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_909),
.Y(n_1192)
);

AOI221xp5_ASAP7_75t_SL g1193 ( 
.A1(n_979),
.A2(n_337),
.B1(n_431),
.B2(n_267),
.C(n_273),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_897),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_911),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_857),
.A2(n_823),
.B1(n_818),
.B2(n_816),
.Y(n_1196)
);

INVx3_ASAP7_75t_SL g1197 ( 
.A(n_976),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_917),
.B(n_920),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_845),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_986),
.A2(n_823),
.B1(n_818),
.B2(n_816),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_951),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_R g1202 ( 
.A(n_916),
.B(n_254),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_916),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_923),
.B(n_710),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_899),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_900),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1045),
.B(n_925),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1014),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1021),
.B(n_907),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1147),
.B(n_918),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1146),
.A2(n_961),
.B(n_974),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1080),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1020),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_SL g1214 ( 
.A1(n_1023),
.A2(n_1046),
.B(n_1024),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1108),
.A2(n_843),
.B(n_877),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1069),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1039),
.B(n_951),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1128),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1054),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1128),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1199),
.A2(n_883),
.B(n_863),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1040),
.A2(n_938),
.B(n_926),
.C(n_932),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1196),
.A2(n_854),
.B(n_846),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1041),
.B(n_312),
.Y(n_1224)
);

BUFx2_ASAP7_75t_SL g1225 ( 
.A(n_1041),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1027),
.B(n_927),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1094),
.B(n_933),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1029),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1200),
.A2(n_856),
.B(n_855),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1064),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1117),
.A2(n_908),
.B(n_989),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1194),
.B(n_934),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_843),
.B(n_877),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1064),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1118),
.A2(n_984),
.B(n_983),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1194),
.A2(n_939),
.B(n_990),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1108),
.A2(n_913),
.B(n_905),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1193),
.A2(n_987),
.B(n_985),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1205),
.B(n_943),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1141),
.A2(n_1003),
.A3(n_992),
.B(n_948),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1029),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1166),
.A2(n_918),
.B1(n_959),
.B2(n_947),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1033),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1064),
.Y(n_1245)
);

AO32x2_ASAP7_75t_L g1246 ( 
.A1(n_1088),
.A2(n_816),
.A3(n_913),
.B1(n_905),
.B2(n_998),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1016),
.B(n_945),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1031),
.A2(n_982),
.B1(n_950),
.B2(n_956),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1206),
.B(n_949),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1031),
.A2(n_965),
.B1(n_969),
.B2(n_958),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1127),
.A2(n_999),
.B(n_1000),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1111),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1055),
.B(n_749),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1108),
.A2(n_746),
.B(n_731),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1150),
.A2(n_553),
.A3(n_568),
.B(n_551),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1108),
.A2(n_1035),
.B(n_1031),
.Y(n_1256)
);

O2A1O1Ixp5_ASAP7_75t_L g1257 ( 
.A1(n_1051),
.A2(n_1005),
.B(n_1008),
.C(n_1002),
.Y(n_1257)
);

BUFx5_ASAP7_75t_L g1258 ( 
.A(n_1201),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1174),
.A2(n_1011),
.B(n_809),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1033),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1167),
.A2(n_1175),
.A3(n_1176),
.B(n_1174),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1047),
.A2(n_830),
.B1(n_828),
.B2(n_746),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1167),
.A2(n_428),
.B(n_440),
.C(n_427),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1068),
.B(n_1142),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1035),
.A2(n_746),
.B1(n_768),
.B2(n_731),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1035),
.A2(n_746),
.B(n_731),
.Y(n_1266)
);

OAI22x1_ASAP7_75t_L g1267 ( 
.A1(n_1184),
.A2(n_263),
.B1(n_271),
.B2(n_265),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1176),
.A2(n_809),
.B(n_785),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1198),
.A2(n_835),
.B(n_834),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1054),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1175),
.A2(n_287),
.B(n_292),
.C(n_284),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1080),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1038),
.A2(n_1044),
.B(n_1059),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1043),
.A2(n_832),
.B(n_756),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1170),
.B(n_756),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1180),
.A2(n_832),
.B(n_765),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1034),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1043),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1144),
.B(n_282),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1186),
.A2(n_765),
.B(n_757),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1045),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1049),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1049),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1028),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1067),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1147),
.B(n_731),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1170),
.B(n_757),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1025),
.B(n_248),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1050),
.Y(n_1289)
);

AOI221x1_ASAP7_75t_L g1290 ( 
.A1(n_1019),
.A2(n_284),
.B1(n_287),
.B2(n_421),
.C(n_431),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1032),
.B(n_775),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1052),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1107),
.B(n_775),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1052),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1076),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1144),
.B(n_285),
.Y(n_1296)
);

AOI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1076),
.A2(n_777),
.B(n_776),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1069),
.B(n_288),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1038),
.A2(n_746),
.B1(n_768),
.B2(n_731),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1119),
.A2(n_297),
.B(n_292),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1081),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1014),
.Y(n_1302)
);

INVxp67_ASAP7_75t_SL g1303 ( 
.A(n_1038),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1018),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1092),
.B(n_290),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1180),
.A2(n_777),
.B(n_776),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1099),
.A2(n_579),
.A3(n_568),
.B(n_301),
.Y(n_1307)
);

OAI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1092),
.A2(n_296),
.B(n_294),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1135),
.A2(n_830),
.B(n_828),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1131),
.A2(n_579),
.B(n_651),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1147),
.B(n_768),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1025),
.B(n_248),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1131),
.A2(n_579),
.B(n_484),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1147),
.B(n_768),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1061),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1067),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1107),
.B(n_768),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1099),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1044),
.A2(n_783),
.B(n_779),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1044),
.A2(n_783),
.B(n_779),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1131),
.A2(n_484),
.B(n_482),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1145),
.B(n_300),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1066),
.A2(n_492),
.B(n_490),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1066),
.A2(n_492),
.B(n_490),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1104),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1084),
.A2(n_497),
.B(n_493),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1103),
.A2(n_392),
.A3(n_308),
.B(n_319),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1015),
.B(n_779),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1072),
.B(n_1085),
.Y(n_1329)
);

BUFx4_ASAP7_75t_SL g1330 ( 
.A(n_1065),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1062),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1084),
.A2(n_497),
.B(n_493),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1183),
.A2(n_783),
.B(n_779),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1172),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1093),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1015),
.B(n_779),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1017),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1103),
.A2(n_500),
.B(n_499),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1129),
.A2(n_830),
.B(n_828),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1098),
.A2(n_500),
.B(n_499),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1098),
.A2(n_506),
.B(n_503),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1071),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1104),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1097),
.B(n_783),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1172),
.B(n_783),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1106),
.A2(n_506),
.B(n_503),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1098),
.A2(n_1110),
.B(n_1165),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_SL g1348 ( 
.A1(n_1097),
.A2(n_308),
.B(n_297),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1104),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1062),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1071),
.Y(n_1351)
);

OAI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1083),
.A2(n_1155),
.B(n_1077),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1183),
.A2(n_817),
.B(n_784),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1104),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1172),
.B(n_784),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1017),
.Y(n_1356)
);

NOR2x1_ASAP7_75t_L g1357 ( 
.A(n_1042),
.B(n_1028),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1030),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1165),
.A2(n_329),
.B(n_325),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1153),
.B(n_784),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1172),
.B(n_784),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1165),
.A2(n_329),
.B(n_325),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1145),
.B(n_303),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1138),
.B(n_307),
.Y(n_1364)
);

BUFx4f_ASAP7_75t_L g1365 ( 
.A(n_1075),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1073),
.B(n_248),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1063),
.B(n_1184),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1030),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1096),
.A2(n_336),
.B(n_335),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1100),
.A2(n_336),
.B(n_335),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1209),
.B(n_1226),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1268),
.A2(n_1101),
.B(n_1106),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1252),
.B(n_1342),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1218),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1220),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1278),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1268),
.A2(n_1113),
.B(n_1160),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1238),
.A2(n_1070),
.B(n_1183),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1227),
.B(n_1217),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1369),
.A2(n_1164),
.B(n_1113),
.Y(n_1381)
);

AOI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_1279),
.A2(n_1159),
.B1(n_1181),
.B2(n_1185),
.C(n_1074),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1261),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1210),
.B(n_1147),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1212),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1261),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1259),
.A2(n_1105),
.B(n_1089),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1222),
.A2(n_1091),
.B(n_1157),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1315),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1259),
.A2(n_1105),
.B(n_1089),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1276),
.A2(n_1114),
.B(n_1109),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1276),
.A2(n_1114),
.B(n_1109),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1313),
.A2(n_1125),
.B(n_1122),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1270),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1331),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1219),
.B(n_1139),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1313),
.A2(n_1125),
.B(n_1122),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1347),
.A2(n_1214),
.B(n_1310),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1282),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1210),
.B(n_1104),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1279),
.A2(n_1296),
.B(n_1329),
.C(n_1352),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1264),
.A2(n_1060),
.B1(n_1012),
.B2(n_1188),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1240),
.B(n_1168),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1232),
.B(n_1102),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1300),
.A2(n_1153),
.B(n_1189),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1237),
.B(n_1123),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1252),
.B(n_1172),
.Y(n_1407)
);

CKINVDCx6p67_ASAP7_75t_R g1408 ( 
.A(n_1285),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1347),
.A2(n_1154),
.B(n_1148),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1310),
.A2(n_1154),
.B(n_1148),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1222),
.A2(n_1178),
.B(n_1171),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1272),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1247),
.A2(n_1173),
.B(n_1060),
.C(n_1012),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1261),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1306),
.A2(n_1163),
.B(n_1162),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1263),
.A2(n_1133),
.A3(n_1143),
.B(n_1132),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1296),
.A2(n_1197),
.B(n_1075),
.C(n_1195),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1369),
.A2(n_1133),
.B(n_1132),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1283),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1329),
.B(n_1179),
.Y(n_1420)
);

OAI222xp33_ASAP7_75t_L g1421 ( 
.A1(n_1363),
.A2(n_1185),
.B1(n_1187),
.B2(n_1086),
.C1(n_1065),
.C2(n_1155),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1351),
.B(n_1161),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1306),
.A2(n_1163),
.B(n_1162),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1370),
.A2(n_1149),
.B(n_1143),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1339),
.A2(n_1204),
.B(n_1158),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1221),
.A2(n_1057),
.B(n_1156),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1230),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1274),
.A2(n_1151),
.B(n_1149),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1297),
.A2(n_1152),
.B(n_1151),
.Y(n_1430)
);

NAND2x1_ASAP7_75t_L g1431 ( 
.A(n_1230),
.B(n_1234),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1288),
.B(n_1095),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1289),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1323),
.A2(n_1326),
.B(n_1324),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1292),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1323),
.A2(n_1152),
.B(n_1136),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1213),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1208),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1177),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1363),
.A2(n_1060),
.B1(n_1012),
.B2(n_1079),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1324),
.A2(n_1136),
.B(n_1120),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1208),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1365),
.B(n_1116),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1230),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1294),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1207),
.A2(n_1079),
.B1(n_1073),
.B2(n_1078),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1326),
.A2(n_1136),
.B(n_1120),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1332),
.A2(n_1120),
.B(n_1112),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1332),
.A2(n_1124),
.B(n_1112),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1312),
.B(n_1095),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1247),
.B(n_1073),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1295),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1229),
.A2(n_1124),
.B(n_1112),
.Y(n_1453)
);

AO32x2_ASAP7_75t_L g1454 ( 
.A1(n_1243),
.A2(n_1248),
.A3(n_1250),
.B1(n_1246),
.B2(n_1265),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1302),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1322),
.B(n_1036),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1301),
.Y(n_1457)
);

AND2x6_ASAP7_75t_L g1458 ( 
.A(n_1230),
.B(n_1090),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1229),
.A2(n_1048),
.B(n_1037),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1223),
.A2(n_1202),
.B(n_1169),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1234),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1318),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1340),
.A2(n_1048),
.B(n_1037),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1286),
.B(n_1115),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1340),
.A2(n_1056),
.B(n_1053),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1228),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1341),
.A2(n_1056),
.B(n_1053),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1216),
.B(n_1177),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1234),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1284),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1242),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1364),
.A2(n_1197),
.B(n_1075),
.C(n_1271),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1244),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1257),
.A2(n_1137),
.B(n_1079),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1260),
.A2(n_1303),
.B1(n_1177),
.B2(n_1317),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1370),
.A2(n_1022),
.B(n_346),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1236),
.B(n_1177),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1341),
.A2(n_1130),
.B(n_1121),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1253),
.B(n_1249),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1302),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1223),
.A2(n_1130),
.B(n_1121),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1211),
.A2(n_1192),
.B(n_346),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1263),
.A2(n_337),
.A3(n_441),
.B(n_356),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1359),
.A2(n_358),
.B(n_356),
.Y(n_1484)
);

NOR2xp67_ASAP7_75t_L g1485 ( 
.A(n_1277),
.B(n_1093),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1331),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1359),
.A2(n_374),
.B(n_358),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1362),
.A2(n_392),
.B(n_374),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1362),
.A2(n_402),
.B(n_400),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1337),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1211),
.A2(n_1126),
.B(n_1137),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1337),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1317),
.A2(n_1177),
.B1(n_1078),
.B2(n_1140),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1256),
.A2(n_1191),
.B(n_1090),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1364),
.A2(n_1197),
.B(n_1271),
.C(n_1224),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1321),
.A2(n_1192),
.B(n_402),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1231),
.A2(n_412),
.B(n_400),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1321),
.A2(n_1192),
.B(n_421),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1277),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1330),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1365),
.B(n_1078),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1328),
.A2(n_1190),
.B(n_1139),
.C(n_1137),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1348),
.A2(n_1273),
.B(n_1338),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1309),
.A2(n_1111),
.B(n_441),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1284),
.Y(n_1505)
);

NOR2xp67_ASAP7_75t_L g1506 ( 
.A(n_1298),
.B(n_1058),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_L g1507 ( 
.A(n_1298),
.B(n_1058),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1356),
.Y(n_1508)
);

AO31x2_ASAP7_75t_L g1509 ( 
.A1(n_1290),
.A2(n_412),
.A3(n_1026),
.B(n_1086),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1356),
.B(n_1111),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1231),
.A2(n_1192),
.B(n_1190),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_R g1512 ( 
.A(n_1270),
.B(n_1225),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1308),
.A2(n_423),
.B1(n_317),
.B2(n_318),
.C(n_327),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1251),
.A2(n_1192),
.B(n_1190),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1235),
.A2(n_1346),
.B(n_1251),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1350),
.A2(n_1182),
.B1(n_1013),
.B2(n_1190),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1358),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_SL g1518 ( 
.A1(n_1286),
.A2(n_1201),
.B(n_1139),
.C(n_1036),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1358),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1336),
.A2(n_1139),
.B(n_1203),
.C(n_1140),
.Y(n_1520)
);

NOR3xp33_ASAP7_75t_SL g1521 ( 
.A(n_1367),
.B(n_1013),
.C(n_339),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_SL g1522 ( 
.A1(n_1291),
.A2(n_1201),
.B(n_1203),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1235),
.A2(n_348),
.B(n_313),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1215),
.A2(n_1090),
.B(n_1203),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1367),
.A2(n_1304),
.B1(n_1366),
.B2(n_1305),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1368),
.B(n_1203),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1262),
.A2(n_1203),
.B(n_1140),
.C(n_1134),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1233),
.A2(n_1134),
.B(n_1115),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1368),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1269),
.A2(n_352),
.B(n_349),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1266),
.A2(n_1134),
.B(n_1115),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1319),
.A2(n_1134),
.B(n_1115),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1275),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1311),
.B(n_1115),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1345),
.B(n_1140),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1307),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1287),
.B(n_1219),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1320),
.A2(n_1353),
.B(n_1333),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1254),
.A2(n_1134),
.B(n_1087),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1219),
.B(n_1140),
.Y(n_1540)
);

BUFx8_ASAP7_75t_SL g1541 ( 
.A(n_1285),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1280),
.A2(n_1087),
.B(n_830),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1311),
.B(n_784),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1327),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1314),
.A2(n_357),
.B(n_354),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1267),
.A2(n_391),
.B1(n_393),
.B2(n_1082),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1293),
.B(n_1087),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1314),
.A2(n_1087),
.B(n_830),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1299),
.A2(n_830),
.B(n_828),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1307),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1317),
.B(n_361),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1422),
.B(n_1327),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1486),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1438),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1371),
.B(n_1357),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1385),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1234),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1541),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1438),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1403),
.B(n_1327),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1419),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1380),
.B(n_1361),
.Y(n_1562)
);

CKINVDCx16_ASAP7_75t_R g1563 ( 
.A(n_1486),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1401),
.A2(n_1245),
.B1(n_1361),
.B2(n_1355),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1500),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1456),
.A2(n_1316),
.B1(n_1335),
.B2(n_330),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1382),
.A2(n_330),
.B1(n_437),
.B2(n_393),
.Y(n_1567)
);

CKINVDCx14_ASAP7_75t_R g1568 ( 
.A(n_1500),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1419),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1533),
.B(n_1361),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1422),
.B(n_1327),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1420),
.B(n_1307),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1432),
.B(n_391),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1412),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1440),
.A2(n_1245),
.B1(n_1355),
.B2(n_1345),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1442),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1442),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1451),
.A2(n_1245),
.B1(n_1355),
.B2(n_1345),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1383),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1411),
.A2(n_437),
.B1(n_330),
.B2(n_393),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1404),
.B(n_1325),
.Y(n_1581)
);

AO31x2_ASAP7_75t_L g1582 ( 
.A1(n_1536),
.A2(n_1360),
.A3(n_1344),
.B(n_1246),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1432),
.A2(n_1335),
.B1(n_1316),
.B2(n_330),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1470),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1495),
.A2(n_1246),
.B(n_1354),
.C(n_1325),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1383),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1404),
.B(n_1325),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1458),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1535),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1396),
.B(n_1354),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1450),
.A2(n_437),
.B1(n_391),
.B2(n_393),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1450),
.A2(n_437),
.B1(n_391),
.B2(n_362),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1455),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1505),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1455),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1525),
.A2(n_1258),
.B1(n_364),
.B2(n_438),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1546),
.A2(n_435),
.B1(n_375),
.B2(n_378),
.Y(n_1597)
);

AOI222xp33_ASAP7_75t_L g1598 ( 
.A1(n_1421),
.A2(n_371),
.B1(n_383),
.B2(n_394),
.C1(n_395),
.C2(n_397),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1437),
.Y(n_1599)
);

CKINVDCx12_ASAP7_75t_R g1600 ( 
.A(n_1512),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1406),
.B(n_1307),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1535),
.B(n_1354),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1406),
.B(n_401),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1468),
.B(n_403),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1388),
.A2(n_447),
.B1(n_406),
.B2(n_407),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1452),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1427),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_SL g1608 ( 
.A1(n_1472),
.A2(n_1239),
.B(n_1258),
.Y(n_1608)
);

AOI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1417),
.A2(n_1239),
.B(n_1349),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1540),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1396),
.B(n_1343),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1468),
.B(n_405),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1479),
.A2(n_451),
.B1(n_416),
.B2(n_417),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1386),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1468),
.B(n_413),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1386),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1511),
.A2(n_1255),
.B(n_1246),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1396),
.B(n_1343),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1471),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1503),
.A2(n_1255),
.B(n_1241),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1374),
.B(n_419),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1513),
.A2(n_450),
.B1(n_422),
.B2(n_425),
.C(n_426),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1551),
.B(n_1255),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1389),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1374),
.B(n_420),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1537),
.B(n_434),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1503),
.A2(n_1255),
.B(n_1241),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1395),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1375),
.Y(n_1629)
);

INVx3_ASAP7_75t_SL g1630 ( 
.A(n_1395),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1373),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1396),
.B(n_1343),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1374),
.B(n_436),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1428),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1446),
.B(n_1413),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1521),
.A2(n_443),
.B1(n_445),
.B2(n_452),
.C(n_455),
.Y(n_1636)
);

OR2x6_ASAP7_75t_L g1637 ( 
.A(n_1474),
.B(n_1349),
.Y(n_1637)
);

CKINVDCx11_ASAP7_75t_R g1638 ( 
.A(n_1394),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1402),
.A2(n_1258),
.B1(n_456),
.B2(n_1349),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1426),
.A2(n_1258),
.B1(n_828),
.B2(n_676),
.Y(n_1640)
);

NOR4xp25_ASAP7_75t_L g1641 ( 
.A(n_1518),
.B(n_6),
.C(n_8),
.D(n_11),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1540),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1443),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1477),
.A2(n_1258),
.B1(n_828),
.B2(n_676),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1477),
.A2(n_1258),
.B1(n_676),
.B2(n_668),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1506),
.B(n_1241),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1508),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1379),
.A2(n_1241),
.B(n_632),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_SL g1649 ( 
.A(n_1516),
.B(n_13),
.C(n_14),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1507),
.B(n_16),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_R g1651 ( 
.A(n_1545),
.B(n_114),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1376),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1377),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1399),
.B(n_18),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1433),
.A2(n_676),
.B1(n_668),
.B2(n_656),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1535),
.B(n_122),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1527),
.B(n_817),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1435),
.A2(n_1457),
.B1(n_1462),
.B2(n_1445),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1466),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_SL g1660 ( 
.A(n_1499),
.B(n_23),
.C(n_25),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1510),
.B(n_26),
.Y(n_1661)
);

CKINVDCx6p67_ASAP7_75t_R g1662 ( 
.A(n_1394),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1407),
.B(n_1439),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1508),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1473),
.B(n_1510),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1480),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1490),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1540),
.Y(n_1668)
);

BUFx4f_ASAP7_75t_SL g1669 ( 
.A(n_1408),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1407),
.B(n_28),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1407),
.B(n_123),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1517),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1540),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1439),
.B(n_125),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1439),
.B(n_138),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1511),
.A2(n_817),
.B(n_656),
.Y(n_1676)
);

OAI222xp33_ASAP7_75t_L g1677 ( 
.A1(n_1493),
.A2(n_1475),
.B1(n_1384),
.B2(n_1547),
.C1(n_1499),
.C2(n_1492),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1520),
.A2(n_1485),
.B1(n_1384),
.B2(n_1502),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1384),
.A2(n_817),
.B1(n_710),
.B2(n_676),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1373),
.Y(n_1680)
);

INVx4_ASAP7_75t_SL g1681 ( 
.A(n_1458),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1526),
.B(n_148),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1400),
.A2(n_817),
.B1(n_710),
.B2(n_676),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1400),
.B(n_31),
.C(n_32),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1517),
.B(n_35),
.Y(n_1685)
);

AOI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1544),
.A2(n_1550),
.B(n_1536),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1460),
.A2(n_676),
.B1(n_668),
.B2(n_656),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1458),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1476),
.A2(n_668),
.B1(n_656),
.B2(n_37),
.C(n_38),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1529),
.B(n_35),
.Y(n_1690)
);

BUFx4f_ASAP7_75t_L g1691 ( 
.A(n_1408),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1428),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1414),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1529),
.B(n_36),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1526),
.B(n_153),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1519),
.B(n_36),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_R g1697 ( 
.A(n_1545),
.B(n_1530),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1415),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1415),
.Y(n_1699)
);

NAND2x1_ASAP7_75t_L g1700 ( 
.A(n_1458),
.B(n_656),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_R g1701 ( 
.A(n_1545),
.B(n_154),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1414),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1444),
.B(n_158),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1460),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1444),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1460),
.A2(n_668),
.B1(n_656),
.B2(n_46),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1400),
.A2(n_668),
.B1(n_656),
.B2(n_46),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1405),
.A2(n_668),
.B1(n_45),
.B2(n_47),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_L g1709 ( 
.A(n_1550),
.B(n_40),
.C(n_47),
.D(n_50),
.Y(n_1709)
);

INVx4_ASAP7_75t_SL g1710 ( 
.A(n_1458),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1405),
.A2(n_51),
.B1(n_53),
.B2(n_60),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1522),
.B(n_232),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1453),
.A2(n_202),
.B(n_221),
.Y(n_1713)
);

CKINVDCx6p67_ASAP7_75t_R g1714 ( 
.A(n_1428),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1428),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1428),
.B(n_1461),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1458),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1494),
.A2(n_196),
.B(n_220),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1461),
.B(n_62),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1541),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1476),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1476),
.B(n_66),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1509),
.B(n_74),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1483),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1469),
.Y(n_1725)
);

OAI22x1_ASAP7_75t_L g1726 ( 
.A1(n_1476),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1461),
.B(n_75),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1461),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1464),
.A2(n_1534),
.B1(n_1545),
.B2(n_1469),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1483),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1504),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1416),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_L g1733 ( 
.A1(n_1482),
.A2(n_81),
.B(n_83),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1483),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1483),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1444),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1461),
.B(n_165),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1509),
.B(n_87),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1464),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_1739)
);

AND2x6_ASAP7_75t_L g1740 ( 
.A(n_1522),
.B(n_1454),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1431),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1509),
.B(n_89),
.Y(n_1742)
);

OR2x6_ASAP7_75t_SL g1743 ( 
.A(n_1509),
.B(n_92),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1416),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1561),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1569),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1567),
.A2(n_1504),
.B1(n_1425),
.B2(n_1381),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1567),
.A2(n_1504),
.B1(n_1491),
.B2(n_1425),
.C(n_1534),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1649),
.A2(n_1580),
.B1(n_1727),
.B2(n_1719),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1629),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1562),
.B(n_1509),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1728),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1580),
.A2(n_1425),
.B1(n_1381),
.B2(n_1418),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1660),
.A2(n_1381),
.B1(n_1424),
.B2(n_1418),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1596),
.A2(n_1464),
.B1(n_1534),
.B2(n_1543),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1709),
.A2(n_1381),
.B1(n_1418),
.B2(n_1424),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1566),
.A2(n_1491),
.B1(n_1530),
.B2(n_1523),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1659),
.A2(n_1605),
.B1(n_1591),
.B2(n_1592),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_L g1759 ( 
.A(n_1605),
.B(n_1613),
.C(n_1597),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1555),
.B(n_1483),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1552),
.B(n_1416),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1597),
.A2(n_1523),
.B1(n_1530),
.B2(n_1543),
.C(n_1431),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1643),
.A2(n_1739),
.B1(n_1635),
.B2(n_1689),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1652),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1571),
.B(n_1530),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1659),
.A2(n_1491),
.B1(n_1543),
.B2(n_1454),
.C(n_97),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1579),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1591),
.A2(n_1418),
.B1(n_1424),
.B2(n_1489),
.Y(n_1768)
);

OAI21xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1731),
.A2(n_1539),
.B(n_1524),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1613),
.A2(n_1523),
.B1(n_1424),
.B2(n_1487),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1592),
.A2(n_1523),
.B1(n_1487),
.B2(n_1488),
.C(n_1489),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1598),
.A2(n_93),
.B(n_94),
.C(n_95),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1673),
.A2(n_1711),
.B1(n_1727),
.B2(n_1719),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1574),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1606),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1673),
.A2(n_1489),
.B1(n_1484),
.B2(n_1488),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1556),
.B(n_1416),
.Y(n_1777)
);

OAI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1743),
.A2(n_1487),
.B1(n_1484),
.B2(n_1488),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1641),
.A2(n_1454),
.B1(n_95),
.B2(n_98),
.C(n_99),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1684),
.A2(n_1497),
.B(n_1488),
.C(n_1489),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1653),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1626),
.B(n_166),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1607),
.A2(n_1624),
.B1(n_1584),
.B2(n_1619),
.C1(n_103),
.C2(n_104),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1661),
.B(n_1416),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1663),
.B(n_1482),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1583),
.A2(n_1514),
.B1(n_1484),
.B2(n_1487),
.Y(n_1786)
);

NAND2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1588),
.B(n_1514),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1572),
.B(n_1497),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1563),
.B(n_172),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1579),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1702),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1573),
.A2(n_1484),
.B1(n_1481),
.B2(n_1498),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1610),
.B(n_1496),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1663),
.B(n_1498),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1622),
.A2(n_1497),
.B1(n_1515),
.B2(n_1454),
.C(n_103),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1610),
.B(n_1496),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1631),
.Y(n_1797)
);

NAND2x1_ASAP7_75t_L g1798 ( 
.A(n_1588),
.B(n_1515),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1711),
.A2(n_1708),
.B1(n_1725),
.B2(n_1639),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1708),
.A2(n_1497),
.B1(n_1515),
.B2(n_1454),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1725),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1663),
.B(n_1481),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1603),
.A2(n_1515),
.B1(n_1478),
.B2(n_1524),
.Y(n_1803)
);

OAI21xp33_ASAP7_75t_L g1804 ( 
.A1(n_1731),
.A2(n_1398),
.B(n_1459),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1726),
.A2(n_93),
.B1(n_99),
.B2(n_101),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1553),
.A2(n_101),
.B1(n_106),
.B2(n_108),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1636),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.C(n_1538),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1706),
.A2(n_1459),
.B1(n_1430),
.B2(n_1429),
.C(n_1378),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1604),
.B(n_1430),
.Y(n_1809)
);

BUFx2_ASAP7_75t_R g1810 ( 
.A(n_1558),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1680),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1642),
.B(n_1409),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1586),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1704),
.A2(n_1398),
.B(n_1409),
.C(n_1378),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1612),
.B(n_1429),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1706),
.A2(n_1372),
.B1(n_1387),
.B2(n_1390),
.C(n_1448),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1560),
.B(n_1372),
.Y(n_1817)
);

AOI222xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1740),
.A2(n_585),
.B1(n_181),
.B2(n_182),
.C1(n_187),
.C2(n_194),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1680),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1565),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1717),
.A2(n_1387),
.B1(n_1390),
.B2(n_1478),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1599),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1557),
.A2(n_1548),
.B1(n_1539),
.B2(n_1531),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1721),
.A2(n_1423),
.B1(n_1391),
.B2(n_1392),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1733),
.A2(n_1449),
.B1(n_1448),
.B2(n_1423),
.C(n_1392),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_L g1826 ( 
.A1(n_1650),
.A2(n_1548),
.B1(n_195),
.B2(n_204),
.C(n_206),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1693),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1742),
.A2(n_1528),
.B1(n_1531),
.B2(n_1532),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1654),
.A2(n_1449),
.B1(n_1467),
.B2(n_1465),
.Y(n_1829)
);

OAI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1712),
.A2(n_177),
.B1(n_210),
.B2(n_212),
.C1(n_213),
.C2(n_217),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1723),
.A2(n_1738),
.B1(n_1722),
.B2(n_1633),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1678),
.B(n_1528),
.Y(n_1832)
);

OAI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1670),
.A2(n_1436),
.B(n_1467),
.C(n_1465),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1553),
.A2(n_1542),
.B1(n_1532),
.B2(n_1549),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1621),
.A2(n_1391),
.B1(n_1463),
.B2(n_1436),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1625),
.A2(n_1463),
.B1(n_1393),
.B2(n_1397),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1693),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1615),
.A2(n_1701),
.B1(n_1651),
.B2(n_1691),
.C(n_1718),
.Y(n_1838)
);

CKINVDCx6p67_ASAP7_75t_R g1839 ( 
.A(n_1630),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1696),
.B(n_219),
.Y(n_1840)
);

AOI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1623),
.A2(n_1441),
.B(n_1447),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1628),
.B(n_1542),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_SL g1843 ( 
.A(n_1637),
.B(n_1447),
.Y(n_1843)
);

AOI222xp33_ASAP7_75t_L g1844 ( 
.A1(n_1638),
.A2(n_1549),
.B1(n_585),
.B2(n_1441),
.C1(n_1397),
.C2(n_1393),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1601),
.A2(n_1410),
.B1(n_1434),
.B2(n_585),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_SL g1846 ( 
.A1(n_1585),
.A2(n_1657),
.B(n_1658),
.C(n_1694),
.Y(n_1846)
);

OA21x2_ASAP7_75t_L g1847 ( 
.A1(n_1585),
.A2(n_1617),
.B(n_1609),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1638),
.A2(n_1570),
.B1(n_1712),
.B2(n_1707),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1557),
.A2(n_1691),
.B1(n_1630),
.B2(n_1594),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1581),
.B(n_1587),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1642),
.B(n_1668),
.Y(n_1851)
);

OR2x6_ASAP7_75t_L g1852 ( 
.A(n_1637),
.B(n_1712),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1665),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1589),
.B(n_1602),
.Y(n_1854)
);

BUFx2_ASAP7_75t_SL g1855 ( 
.A(n_1728),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1658),
.A2(n_1671),
.B1(n_1685),
.B2(n_1690),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1634),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1669),
.A2(n_1637),
.B1(n_1645),
.B2(n_1568),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1714),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1671),
.A2(n_1675),
.B1(n_1674),
.B2(n_1656),
.Y(n_1860)
);

OAI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1646),
.A2(n_1687),
.B(n_1648),
.C(n_1640),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1640),
.A2(n_1716),
.B(n_1564),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1669),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1651),
.A2(n_1701),
.B1(n_1688),
.B2(n_1611),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1589),
.B(n_1602),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1671),
.A2(n_1674),
.B1(n_1675),
.B2(n_1656),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1645),
.A2(n_1568),
.B1(n_1668),
.B2(n_1644),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1602),
.Y(n_1868)
);

CKINVDCx6p67_ASAP7_75t_R g1869 ( 
.A(n_1565),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1716),
.A2(n_1618),
.B(n_1611),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1666),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1688),
.A2(n_1618),
.B1(n_1611),
.B2(n_1575),
.Y(n_1872)
);

OAI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1687),
.A2(n_1697),
.B1(n_1578),
.B2(n_1644),
.C(n_1720),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1677),
.A2(n_1729),
.B1(n_1735),
.B2(n_1734),
.C(n_1730),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1618),
.A2(n_1590),
.B1(n_1695),
.B2(n_1682),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1729),
.A2(n_1724),
.B1(n_1608),
.B2(n_1732),
.C(n_1744),
.Y(n_1876)
);

OA21x2_ASAP7_75t_L g1877 ( 
.A1(n_1698),
.A2(n_1699),
.B(n_1676),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1695),
.A2(n_1662),
.B1(n_1682),
.B2(n_1740),
.Y(n_1878)
);

AO22x2_ASAP7_75t_L g1879 ( 
.A1(n_1698),
.A2(n_1699),
.B1(n_1681),
.B2(n_1710),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1732),
.A2(n_1744),
.B1(n_1667),
.B2(n_1695),
.C(n_1703),
.Y(n_1880)
);

OAI221xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1600),
.A2(n_1655),
.B1(n_1697),
.B2(n_1705),
.C(n_1736),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_1634),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1590),
.B(n_1703),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1554),
.B(n_1559),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1632),
.A2(n_1655),
.B1(n_1703),
.B2(n_1741),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1559),
.Y(n_1886)
);

AND2x6_ASAP7_75t_SL g1887 ( 
.A(n_1737),
.B(n_1632),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1737),
.A2(n_1740),
.B1(n_1741),
.B2(n_1679),
.Y(n_1888)
);

AOI222xp33_ASAP7_75t_L g1889 ( 
.A1(n_1740),
.A2(n_1710),
.B1(n_1681),
.B2(n_1647),
.C1(n_1664),
.C2(n_1593),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1740),
.A2(n_1576),
.B1(n_1577),
.B2(n_1672),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1586),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1577),
.A2(n_1664),
.B1(n_1593),
.B2(n_1595),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1683),
.A2(n_1614),
.B1(n_1616),
.B2(n_1620),
.C(n_1627),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1715),
.B(n_1692),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1713),
.B(n_1616),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1595),
.A2(n_1672),
.B1(n_1647),
.B2(n_1627),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1715),
.B(n_1692),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1700),
.A2(n_1634),
.B1(n_1692),
.B2(n_1686),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1681),
.A2(n_1710),
.B1(n_1620),
.B2(n_1634),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1582),
.B(n_1692),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1582),
.B(n_1610),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1582),
.A2(n_1039),
.B1(n_1040),
.B2(n_1144),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1582),
.A2(n_1039),
.B1(n_1040),
.B2(n_1144),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1552),
.B(n_1571),
.Y(n_1904)
);

AOI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1567),
.A2(n_858),
.B1(n_1040),
.B2(n_1039),
.C(n_851),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1567),
.A2(n_1040),
.B1(n_1039),
.B2(n_858),
.C(n_851),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1561),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1556),
.Y(n_1908)
);

AOI222xp33_ASAP7_75t_L g1909 ( 
.A1(n_1567),
.A2(n_858),
.B1(n_1144),
.B2(n_1040),
.C1(n_1039),
.C2(n_628),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1552),
.B(n_1571),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1596),
.A2(n_1040),
.B1(n_1039),
.B2(n_858),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1567),
.A2(n_1039),
.B1(n_1040),
.B2(n_1144),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1567),
.A2(n_1039),
.B1(n_1040),
.B2(n_1144),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1567),
.A2(n_1039),
.B1(n_1040),
.B2(n_1382),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1567),
.A2(n_1039),
.B1(n_1040),
.B2(n_1382),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_SL g1916 ( 
.A1(n_1566),
.A2(n_1039),
.B1(n_1040),
.B2(n_1144),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1579),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1674),
.A2(n_994),
.B(n_870),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1562),
.B(n_1401),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1596),
.A2(n_1040),
.B1(n_1039),
.B2(n_858),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1751),
.B(n_1919),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1798),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1879),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1904),
.B(n_1910),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1791),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1745),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1877),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1817),
.B(n_1761),
.Y(n_1928)
);

BUFx8_ASAP7_75t_L g1929 ( 
.A(n_1863),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1746),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1767),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1767),
.Y(n_1932)
);

AOI322xp5_ASAP7_75t_L g1933 ( 
.A1(n_1905),
.A2(n_1912),
.A3(n_1913),
.B1(n_1758),
.B2(n_1920),
.C1(n_1911),
.C2(n_1805),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1877),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1765),
.B(n_1784),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1760),
.B(n_1777),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1802),
.B(n_1812),
.Y(n_1937)
);

OR2x6_ASAP7_75t_L g1938 ( 
.A(n_1852),
.B(n_1879),
.Y(n_1938)
);

NOR2x1_ASAP7_75t_R g1939 ( 
.A(n_1820),
.B(n_1801),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1901),
.B(n_1788),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1901),
.B(n_1775),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1906),
.A2(n_1915),
.B(n_1914),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1812),
.B(n_1843),
.Y(n_1943)
);

AOI33xp33_ASAP7_75t_L g1944 ( 
.A1(n_1912),
.A2(n_1913),
.A3(n_1758),
.B1(n_1805),
.B2(n_1763),
.B3(n_1773),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1907),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1900),
.B(n_1797),
.Y(n_1946)
);

NOR2x1_ASAP7_75t_L g1947 ( 
.A(n_1864),
.B(n_1838),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1879),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1811),
.B(n_1819),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1871),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1827),
.B(n_1837),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1790),
.B(n_1813),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1831),
.B(n_1750),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1831),
.B(n_1764),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1781),
.B(n_1890),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1890),
.B(n_1896),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1852),
.B(n_1832),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1793),
.B(n_1796),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1778),
.A2(n_1770),
.B(n_1757),
.Y(n_1959)
);

NOR2xp67_ASAP7_75t_L g1960 ( 
.A(n_1833),
.B(n_1842),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1896),
.B(n_1874),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1891),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1891),
.Y(n_1963)
);

AND2x4_ASAP7_75t_SL g1964 ( 
.A(n_1852),
.B(n_1899),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1908),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1917),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1917),
.B(n_1902),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1884),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1902),
.B(n_1903),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1793),
.B(n_1796),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1903),
.B(n_1850),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1847),
.B(n_1803),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1853),
.B(n_1800),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1787),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1787),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1886),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1785),
.B(n_1876),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1794),
.B(n_1809),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1829),
.B(n_1778),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1815),
.B(n_1854),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1895),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1779),
.B(n_1880),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1895),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1909),
.A2(n_1772),
.B(n_1759),
.C(n_1773),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1895),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1829),
.B(n_1753),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1810),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1769),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1892),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1865),
.B(n_1753),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1823),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1756),
.B(n_1878),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1834),
.B(n_1851),
.Y(n_1993)
);

AO21x2_ASAP7_75t_L g1994 ( 
.A1(n_1841),
.A2(n_1771),
.B(n_1804),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1754),
.B(n_1864),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1754),
.B(n_1756),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1792),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1916),
.A2(n_1799),
.B1(n_1749),
.B2(n_1807),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1892),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1878),
.B(n_1888),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1857),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1848),
.A2(n_1782),
.B1(n_1766),
.B2(n_1856),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1856),
.B(n_1846),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1893),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1828),
.B(n_1889),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1898),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1747),
.B(n_1851),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1748),
.B(n_1747),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1883),
.B(n_1868),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1780),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1768),
.B(n_1786),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1776),
.B(n_1768),
.Y(n_2012)
);

BUFx2_ASAP7_75t_SL g2013 ( 
.A(n_1882),
.Y(n_2013)
);

INVxp67_ASAP7_75t_SL g2014 ( 
.A(n_1825),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1857),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1776),
.B(n_1894),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1862),
.B(n_1861),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1835),
.B(n_1836),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1835),
.B(n_1836),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1897),
.B(n_1821),
.Y(n_2020)
);

NAND3xp33_ASAP7_75t_L g2021 ( 
.A(n_1783),
.B(n_1818),
.C(n_1806),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1821),
.B(n_1857),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1872),
.B(n_1870),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1857),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1824),
.B(n_1845),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1816),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1774),
.B(n_1872),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1752),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1887),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1808),
.Y(n_2030)
);

OAI31xp33_ASAP7_75t_L g2031 ( 
.A1(n_1984),
.A2(n_1830),
.A3(n_1795),
.B(n_1848),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1984),
.A2(n_1867),
.B1(n_1860),
.B2(n_1866),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_2010),
.A2(n_1762),
.B(n_1814),
.Y(n_2033)
);

OAI321xp33_ASAP7_75t_L g2034 ( 
.A1(n_1942),
.A2(n_1881),
.A3(n_1873),
.B1(n_1826),
.B2(n_1858),
.C(n_1755),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1942),
.A2(n_1860),
.B1(n_1866),
.B2(n_1789),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1927),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1945),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1927),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1965),
.B(n_1839),
.Y(n_2039)
);

NAND2xp33_ASAP7_75t_R g2040 ( 
.A(n_1987),
.B(n_1752),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1938),
.B(n_1918),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1940),
.B(n_1845),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1927),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_1944),
.B(n_1849),
.C(n_1840),
.Y(n_2044)
);

OAI221xp5_ASAP7_75t_SL g2045 ( 
.A1(n_1933),
.A2(n_1869),
.B1(n_1822),
.B2(n_1824),
.C(n_1844),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1934),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1945),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1928),
.B(n_1885),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_SL g2049 ( 
.A1(n_2021),
.A2(n_1875),
.B1(n_1859),
.B2(n_1855),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1945),
.Y(n_2050)
);

AOI31xp33_ASAP7_75t_L g2051 ( 
.A1(n_2021),
.A2(n_1939),
.A3(n_1998),
.B(n_1947),
.Y(n_2051)
);

INVxp67_ASAP7_75t_SL g2052 ( 
.A(n_1931),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1940),
.B(n_1935),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1933),
.A2(n_1859),
.B(n_1947),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_2002),
.A2(n_2017),
.B1(n_2004),
.B2(n_2003),
.C(n_2014),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1950),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1982),
.A2(n_1969),
.B1(n_2017),
.B2(n_2029),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1931),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1950),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_1932),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1937),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1928),
.B(n_1946),
.Y(n_2062)
);

OAI31xp33_ASAP7_75t_SL g2063 ( 
.A1(n_2014),
.A2(n_1961),
.A3(n_2005),
.B(n_2000),
.Y(n_2063)
);

OAI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2004),
.A2(n_2003),
.B(n_2030),
.C(n_1982),
.Y(n_2064)
);

NOR5xp2_ASAP7_75t_SL g2065 ( 
.A(n_2030),
.B(n_2029),
.C(n_1960),
.D(n_1939),
.E(n_2027),
.Y(n_2065)
);

INVx4_ASAP7_75t_L g2066 ( 
.A(n_2028),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1935),
.B(n_1978),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1921),
.B(n_1936),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1938),
.Y(n_2069)
);

NOR4xp25_ASAP7_75t_SL g2070 ( 
.A(n_1988),
.B(n_1981),
.C(n_1983),
.D(n_1948),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1965),
.B(n_1921),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2008),
.A2(n_2026),
.B(n_1961),
.C(n_1996),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1950),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_R g2074 ( 
.A(n_1988),
.B(n_2005),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1925),
.Y(n_2075)
);

OAI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2026),
.A2(n_2008),
.B1(n_2023),
.B2(n_2010),
.C(n_2011),
.Y(n_2076)
);

NOR4xp25_ASAP7_75t_SL g2077 ( 
.A(n_1981),
.B(n_1983),
.C(n_1948),
.D(n_2006),
.Y(n_2077)
);

NAND2x1_ASAP7_75t_L g2078 ( 
.A(n_1938),
.B(n_1957),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1938),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1925),
.Y(n_2080)
);

BUFx2_ASAP7_75t_L g2081 ( 
.A(n_1938),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1978),
.B(n_1941),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_SL g2083 ( 
.A1(n_1969),
.A2(n_1992),
.B1(n_2000),
.B2(n_2012),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2012),
.A2(n_1997),
.B1(n_2006),
.B2(n_1977),
.C(n_1971),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1926),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1941),
.B(n_1937),
.Y(n_2086)
);

INVx1_ASAP7_75t_SL g2087 ( 
.A(n_2013),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1937),
.B(n_1990),
.Y(n_2088)
);

OAI211xp5_ASAP7_75t_SL g2089 ( 
.A1(n_2027),
.A2(n_1973),
.B(n_2023),
.C(n_2011),
.Y(n_2089)
);

NAND2xp33_ASAP7_75t_R g2090 ( 
.A(n_1977),
.B(n_1943),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1926),
.Y(n_2091)
);

AND2x6_ASAP7_75t_L g2092 ( 
.A(n_1975),
.B(n_1958),
.Y(n_2092)
);

OAI211xp5_ASAP7_75t_SL g2093 ( 
.A1(n_1973),
.A2(n_1996),
.B(n_1979),
.C(n_1971),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1937),
.B(n_1990),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1992),
.A2(n_2016),
.B1(n_1995),
.B2(n_1954),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1957),
.A2(n_1995),
.B1(n_2013),
.B2(n_1964),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1943),
.B(n_1958),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1930),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1957),
.A2(n_1964),
.B1(n_1979),
.B2(n_1986),
.Y(n_2099)
);

OAI322xp33_ASAP7_75t_L g2100 ( 
.A1(n_1936),
.A2(n_1986),
.A3(n_1989),
.B1(n_1999),
.B2(n_1966),
.C1(n_1946),
.C2(n_1951),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1930),
.Y(n_2101)
);

AOI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_1997),
.A2(n_1953),
.B1(n_1954),
.B2(n_2016),
.C(n_2019),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1980),
.B(n_1970),
.Y(n_2103)
);

AOI21xp33_ASAP7_75t_SL g2104 ( 
.A1(n_1957),
.A2(n_1959),
.B(n_1923),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1980),
.B(n_1970),
.Y(n_2105)
);

AO21x2_ASAP7_75t_L g2106 ( 
.A1(n_1959),
.A2(n_1960),
.B(n_1994),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1953),
.B(n_1976),
.Y(n_2107)
);

OAI211xp5_ASAP7_75t_L g2108 ( 
.A1(n_1997),
.A2(n_1972),
.B(n_2019),
.C(n_2018),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1976),
.B(n_1968),
.Y(n_2109)
);

OAI221xp5_ASAP7_75t_L g2110 ( 
.A1(n_1957),
.A2(n_1985),
.B1(n_1991),
.B2(n_1989),
.C(n_1999),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_2039),
.B(n_1924),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2062),
.B(n_1952),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2037),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2088),
.B(n_1943),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2088),
.B(n_1943),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2037),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2047),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2047),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2094),
.B(n_1958),
.Y(n_2119)
);

INVx1_ASAP7_75t_SL g2120 ( 
.A(n_2062),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2094),
.B(n_1958),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2068),
.B(n_1963),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2050),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2103),
.B(n_1970),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2107),
.B(n_1952),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2058),
.B(n_1991),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2103),
.B(n_1970),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2050),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2060),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2052),
.B(n_1963),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2109),
.B(n_1962),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2056),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2069),
.B(n_1923),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2055),
.B(n_1924),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2105),
.B(n_1923),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_2078),
.B(n_1975),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2056),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2036),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2075),
.B(n_2108),
.Y(n_2139)
);

OR2x6_ASAP7_75t_L g2140 ( 
.A(n_2078),
.B(n_1985),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2105),
.B(n_2007),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2106),
.B(n_1991),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2086),
.B(n_2007),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2086),
.B(n_1993),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2059),
.Y(n_2145)
);

BUFx2_ASAP7_75t_L g2146 ( 
.A(n_2092),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2053),
.B(n_1993),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2059),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2038),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2087),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2073),
.Y(n_2151)
);

NOR2x1_ASAP7_75t_L g2152 ( 
.A(n_2106),
.B(n_2100),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2053),
.B(n_1993),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2073),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2067),
.B(n_1993),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2106),
.B(n_1972),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2069),
.B(n_1959),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2067),
.B(n_1985),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2082),
.B(n_2018),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2080),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2079),
.B(n_1922),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2080),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2082),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2079),
.B(n_1959),
.Y(n_2164)
);

AND2x4_ASAP7_75t_SL g2165 ( 
.A(n_2041),
.B(n_1975),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2081),
.B(n_2020),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_2071),
.B(n_2009),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2043),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2075),
.B(n_1962),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2085),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2085),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2081),
.B(n_1922),
.Y(n_2172)
);

NOR2x1_ASAP7_75t_SL g2173 ( 
.A(n_2041),
.B(n_1994),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2097),
.B(n_2020),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2097),
.B(n_1974),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2102),
.B(n_2091),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2043),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_2046),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2097),
.B(n_1974),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2051),
.B(n_2009),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_2046),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2041),
.B(n_1922),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2091),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2160),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2174),
.B(n_2041),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2174),
.B(n_2061),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_2134),
.B(n_2111),
.Y(n_2187)
);

AOI32xp33_ASAP7_75t_L g2188 ( 
.A1(n_2152),
.A2(n_2072),
.A3(n_2089),
.B1(n_2093),
.B2(n_2057),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2114),
.B(n_2061),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2160),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_2146),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_2139),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2114),
.B(n_2070),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2176),
.B(n_2084),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2176),
.B(n_2095),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2162),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2162),
.Y(n_2197)
);

NOR3xp33_ASAP7_75t_L g2198 ( 
.A(n_2152),
.B(n_2064),
.C(n_2076),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2170),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2122),
.B(n_2083),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2139),
.B(n_2120),
.Y(n_2201)
);

NOR2x1_ASAP7_75t_L g2202 ( 
.A(n_2150),
.B(n_2066),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2181),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2115),
.B(n_2104),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2122),
.B(n_2159),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2181),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2181),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2120),
.B(n_2048),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2157),
.B(n_2048),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2157),
.B(n_2033),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2159),
.B(n_2072),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2129),
.B(n_2167),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2164),
.B(n_2033),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2180),
.A2(n_2054),
.B(n_2031),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2170),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2171),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2181),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2164),
.B(n_2033),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2171),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2183),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2115),
.B(n_2104),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2129),
.B(n_2063),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2126),
.Y(n_2223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2224 ( 
.A1(n_2130),
.A2(n_2110),
.B(n_2065),
.C(n_2074),
.D(n_2099),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2112),
.B(n_2042),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2183),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_2126),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2112),
.B(n_2042),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2131),
.B(n_2101),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2166),
.B(n_2077),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_2146),
.B(n_2092),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2166),
.B(n_2092),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2131),
.B(n_2101),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2125),
.B(n_2098),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_2182),
.B(n_2092),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2125),
.B(n_2098),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2175),
.B(n_2092),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2138),
.Y(n_2238)
);

OAI21xp33_ASAP7_75t_L g2239 ( 
.A1(n_2156),
.A2(n_2032),
.B(n_2044),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2113),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2198),
.B(n_2150),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2209),
.B(n_2156),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2209),
.B(n_2201),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2195),
.B(n_2119),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2232),
.B(n_2140),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_2201),
.B(n_2142),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2239),
.B(n_2143),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_2188),
.B(n_2182),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2208),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2239),
.B(n_2143),
.Y(n_2250)
);

NAND5xp2_ASAP7_75t_SL g2251 ( 
.A(n_2214),
.B(n_2065),
.C(n_2035),
.D(n_2032),
.E(n_2173),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2232),
.B(n_2140),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2192),
.B(n_2141),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2235),
.B(n_2140),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2235),
.B(n_2204),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2235),
.B(n_2140),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2203),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2222),
.B(n_2141),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2235),
.B(n_2140),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2203),
.Y(n_2260)
);

NOR2x1p5_ASAP7_75t_L g2261 ( 
.A(n_2211),
.B(n_2182),
.Y(n_2261)
);

CKINVDCx14_ASAP7_75t_R g2262 ( 
.A(n_2187),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2208),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2212),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2194),
.B(n_2158),
.Y(n_2265)
);

NOR2x1p5_ASAP7_75t_L g2266 ( 
.A(n_2191),
.B(n_2200),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2184),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2203),
.Y(n_2268)
);

BUFx2_ASAP7_75t_L g2269 ( 
.A(n_2202),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2214),
.A2(n_2034),
.B(n_2045),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_2225),
.B(n_2119),
.Y(n_2271)
);

AND2x2_ASAP7_75t_SL g2272 ( 
.A(n_2224),
.B(n_2165),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2184),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2190),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2188),
.B(n_2158),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2190),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_2202),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2185),
.A2(n_2096),
.B1(n_2182),
.B2(n_1994),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2191),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2204),
.B(n_2175),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2228),
.B(n_2155),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2210),
.B(n_2142),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2196),
.Y(n_2283)
);

OR2x2_ASAP7_75t_L g2284 ( 
.A(n_2210),
.B(n_2130),
.Y(n_2284)
);

NOR2x1_ASAP7_75t_L g2285 ( 
.A(n_2230),
.B(n_2113),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2196),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2205),
.B(n_2155),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2234),
.B(n_2147),
.Y(n_2288)
);

INVxp67_ASAP7_75t_L g2289 ( 
.A(n_2230),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2197),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2197),
.Y(n_2291)
);

AOI31xp33_ASAP7_75t_L g2292 ( 
.A1(n_2224),
.A2(n_2040),
.A3(n_2049),
.B(n_2090),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2213),
.B(n_2169),
.Y(n_2293)
);

AND2x4_ASAP7_75t_SL g2294 ( 
.A(n_2231),
.B(n_2133),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2221),
.B(n_2179),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2185),
.B(n_2121),
.Y(n_2296)
);

OAI32xp33_ASAP7_75t_L g2297 ( 
.A1(n_2241),
.A2(n_2213),
.A3(n_2218),
.B1(n_2191),
.B2(n_2193),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2262),
.B(n_2229),
.Y(n_2298)
);

AOI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_2272),
.A2(n_2218),
.B(n_2193),
.Y(n_2299)
);

OAI21xp33_ASAP7_75t_L g2300 ( 
.A1(n_2272),
.A2(n_2233),
.B(n_2221),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2264),
.B(n_2223),
.Y(n_2301)
);

NOR3xp33_ASAP7_75t_L g2302 ( 
.A(n_2270),
.B(n_2289),
.C(n_2292),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2248),
.A2(n_2191),
.B(n_2136),
.Y(n_2303)
);

NOR4xp25_ASAP7_75t_L g2304 ( 
.A(n_2275),
.B(n_2238),
.C(n_2220),
.D(n_2226),
.Y(n_2304)
);

AOI31xp33_ASAP7_75t_L g2305 ( 
.A1(n_2251),
.A2(n_2136),
.A3(n_2231),
.B(n_2227),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2244),
.B(n_2236),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2255),
.B(n_2231),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_2249),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2267),
.Y(n_2309)
);

OAI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2278),
.A2(n_2136),
.B1(n_2215),
.B2(n_2216),
.C(n_2220),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2266),
.A2(n_2231),
.B1(n_2165),
.B2(n_1964),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2267),
.Y(n_2312)
);

CKINVDCx14_ASAP7_75t_R g2313 ( 
.A(n_2269),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2265),
.B(n_2186),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2247),
.B(n_2186),
.Y(n_2315)
);

OAI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2266),
.A2(n_2165),
.B1(n_2133),
.B2(n_2163),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2250),
.B(n_2135),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2279),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2261),
.A2(n_2258),
.B1(n_2269),
.B2(n_2285),
.Y(n_2319)
);

NAND3xp33_ASAP7_75t_L g2320 ( 
.A(n_2263),
.B(n_2238),
.C(n_2219),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2261),
.A2(n_2296),
.B1(n_2251),
.B2(n_2253),
.Y(n_2321)
);

OAI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2277),
.A2(n_2237),
.B1(n_2133),
.B2(n_1975),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2271),
.B(n_2135),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2277),
.A2(n_2237),
.B(n_2189),
.Y(n_2324)
);

OAI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2243),
.A2(n_2025),
.B(n_1956),
.C(n_2238),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2243),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2281),
.B(n_2147),
.Y(n_2327)
);

O2A1O1Ixp5_ASAP7_75t_L g2328 ( 
.A1(n_2255),
.A2(n_2172),
.B(n_2161),
.C(n_2206),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2279),
.Y(n_2329)
);

AOI21xp33_ASAP7_75t_SL g2330 ( 
.A1(n_2245),
.A2(n_2172),
.B(n_2161),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2287),
.B(n_2153),
.Y(n_2331)
);

AOI22x1_ASAP7_75t_L g2332 ( 
.A1(n_2245),
.A2(n_2161),
.B1(n_2172),
.B2(n_2133),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2273),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2288),
.B(n_2280),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2280),
.B(n_2153),
.Y(n_2335)
);

A2O1A1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_2284),
.A2(n_1956),
.B(n_2025),
.C(n_2022),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2284),
.A2(n_2161),
.B(n_2172),
.Y(n_2337)
);

NOR2xp67_ASAP7_75t_SL g2338 ( 
.A(n_2252),
.B(n_2028),
.Y(n_2338)
);

OAI21xp33_ASAP7_75t_L g2339 ( 
.A1(n_2302),
.A2(n_2259),
.B(n_2256),
.Y(n_2339)
);

NAND4xp75_ASAP7_75t_L g2340 ( 
.A(n_2299),
.B(n_2259),
.C(n_2256),
.D(n_2254),
.Y(n_2340)
);

OAI32xp33_ASAP7_75t_SL g2341 ( 
.A1(n_2320),
.A2(n_2246),
.A3(n_2293),
.B1(n_2242),
.B2(n_2282),
.Y(n_2341)
);

AOI21xp33_ASAP7_75t_L g2342 ( 
.A1(n_2297),
.A2(n_2246),
.B(n_2293),
.Y(n_2342)
);

HB1xp67_ASAP7_75t_L g2343 ( 
.A(n_2308),
.Y(n_2343)
);

O2A1O1Ixp33_ASAP7_75t_L g2344 ( 
.A1(n_2313),
.A2(n_2273),
.B(n_2291),
.C(n_2276),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2307),
.B(n_2294),
.Y(n_2345)
);

AOI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2304),
.A2(n_2297),
.B1(n_2319),
.B2(n_2321),
.C(n_2300),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2313),
.A2(n_2294),
.B1(n_2252),
.B2(n_2254),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_2307),
.B(n_2318),
.Y(n_2348)
);

O2A1O1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2305),
.A2(n_2336),
.B(n_2310),
.C(n_2298),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2303),
.B(n_2295),
.Y(n_2350)
);

AOI33xp33_ASAP7_75t_L g2351 ( 
.A1(n_2309),
.A2(n_2276),
.A3(n_2291),
.B1(n_2290),
.B2(n_2286),
.B3(n_2283),
.Y(n_2351)
);

OAI211xp5_ASAP7_75t_L g2352 ( 
.A1(n_2325),
.A2(n_2242),
.B(n_2290),
.C(n_2286),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2298),
.A2(n_1994),
.B1(n_2283),
.B2(n_2274),
.Y(n_2353)
);

OAI21xp33_ASAP7_75t_L g2354 ( 
.A1(n_2326),
.A2(n_2295),
.B(n_2274),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2312),
.Y(n_2355)
);

OAI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_2311),
.A2(n_2189),
.B1(n_2199),
.B2(n_2215),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2336),
.A2(n_2282),
.B(n_2268),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2316),
.A2(n_2092),
.B1(n_2022),
.B2(n_2199),
.Y(n_2358)
);

AOI22xp33_ASAP7_75t_L g2359 ( 
.A1(n_2301),
.A2(n_1967),
.B1(n_2268),
.B2(n_2260),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2333),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2318),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2329),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2330),
.B(n_2173),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2329),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2315),
.Y(n_2365)
);

A2O1A1Ixp33_ASAP7_75t_L g2366 ( 
.A1(n_2328),
.A2(n_2324),
.B(n_2337),
.C(n_2306),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2332),
.A2(n_2260),
.B(n_2257),
.Y(n_2367)
);

OAI21xp5_ASAP7_75t_L g2368 ( 
.A1(n_2332),
.A2(n_2257),
.B(n_2226),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2338),
.A2(n_2092),
.B1(n_2219),
.B2(n_2216),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2343),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2346),
.B(n_2314),
.Y(n_2371)
);

NAND4xp75_ASAP7_75t_L g2372 ( 
.A(n_2342),
.B(n_2334),
.C(n_2317),
.D(n_2335),
.Y(n_2372)
);

XNOR2xp5_ASAP7_75t_L g2373 ( 
.A(n_2340),
.B(n_2323),
.Y(n_2373)
);

NOR2x1_ASAP7_75t_L g2374 ( 
.A(n_2361),
.B(n_2322),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2339),
.B(n_2327),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2355),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2348),
.Y(n_2377)
);

NOR2x1_ASAP7_75t_L g2378 ( 
.A(n_2362),
.B(n_2240),
.Y(n_2378)
);

OAI321xp33_ASAP7_75t_L g2379 ( 
.A1(n_2349),
.A2(n_2331),
.A3(n_2338),
.B1(n_2240),
.B2(n_1967),
.C(n_1974),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2348),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2360),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2351),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2351),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2364),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2365),
.B(n_2217),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2348),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2354),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2347),
.B(n_2217),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2344),
.B(n_2144),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2366),
.B(n_2217),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_2345),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2345),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2356),
.A2(n_2207),
.B1(n_2206),
.B2(n_1929),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2366),
.B(n_2144),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_2391),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2377),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2377),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2380),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2380),
.B(n_2350),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2370),
.B(n_2352),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2386),
.B(n_2353),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2392),
.B(n_2353),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2378),
.Y(n_2403)
);

AOI211x1_ASAP7_75t_L g2404 ( 
.A1(n_2382),
.A2(n_2368),
.B(n_2341),
.C(n_2367),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2387),
.B(n_2359),
.Y(n_2405)
);

AOI211xp5_ASAP7_75t_L g2406 ( 
.A1(n_2371),
.A2(n_2357),
.B(n_2363),
.C(n_2358),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2384),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2383),
.A2(n_2373),
.B(n_2390),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2379),
.B(n_2359),
.Y(n_2409)
);

AOI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2404),
.A2(n_2390),
.B1(n_2375),
.B2(n_2394),
.C(n_2376),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2398),
.Y(n_2411)
);

AOI32xp33_ASAP7_75t_L g2412 ( 
.A1(n_2406),
.A2(n_2374),
.A3(n_2388),
.B1(n_2389),
.B2(n_2381),
.Y(n_2412)
);

O2A1O1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_2408),
.A2(n_2388),
.B(n_2385),
.C(n_2363),
.Y(n_2413)
);

A2O1A1Ixp33_ASAP7_75t_SL g2414 ( 
.A1(n_2398),
.A2(n_2397),
.B(n_2396),
.C(n_2407),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_SL g2415 ( 
.A(n_2395),
.B(n_2400),
.C(n_2409),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2405),
.B(n_2372),
.Y(n_2416)
);

OAI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2409),
.A2(n_2393),
.B1(n_2369),
.B2(n_2385),
.C(n_2207),
.Y(n_2417)
);

NOR2xp67_ASAP7_75t_L g2418 ( 
.A(n_2403),
.B(n_2207),
.Y(n_2418)
);

AOI221x1_ASAP7_75t_L g2419 ( 
.A1(n_2401),
.A2(n_2206),
.B1(n_2169),
.B2(n_2116),
.C(n_2148),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2400),
.B(n_1929),
.C(n_2015),
.Y(n_2420)
);

AOI221xp5_ASAP7_75t_L g2421 ( 
.A1(n_2402),
.A2(n_2128),
.B1(n_2148),
.B2(n_2123),
.C(n_2151),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_L g2422 ( 
.A(n_2399),
.B(n_1929),
.C(n_2024),
.Y(n_2422)
);

AOI211xp5_ASAP7_75t_L g2423 ( 
.A1(n_2410),
.A2(n_2399),
.B(n_2121),
.C(n_2179),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2411),
.Y(n_2424)
);

NAND2x1_ASAP7_75t_L g2425 ( 
.A(n_2411),
.B(n_2066),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2412),
.B(n_2127),
.Y(n_2426)
);

NOR3x2_ASAP7_75t_L g2427 ( 
.A(n_2414),
.B(n_1929),
.C(n_1949),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2415),
.A2(n_2015),
.B1(n_2024),
.B2(n_2028),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2416),
.B(n_2413),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2420),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2424),
.B(n_2418),
.Y(n_2431)
);

XNOR2xp5_ASAP7_75t_L g2432 ( 
.A(n_2427),
.B(n_2422),
.Y(n_2432)
);

OR2x2_ASAP7_75t_L g2433 ( 
.A(n_2429),
.B(n_2426),
.Y(n_2433)
);

NAND3xp33_ASAP7_75t_SL g2434 ( 
.A(n_2430),
.B(n_2417),
.C(n_2421),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2423),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2428),
.Y(n_2436)
);

AND2x4_ASAP7_75t_L g2437 ( 
.A(n_2425),
.B(n_2419),
.Y(n_2437)
);

XNOR2xp5_ASAP7_75t_L g2438 ( 
.A(n_2427),
.B(n_2124),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2431),
.Y(n_2439)
);

NAND5xp2_ASAP7_75t_L g2440 ( 
.A(n_2435),
.B(n_2124),
.C(n_2127),
.D(n_1955),
.E(n_1968),
.Y(n_2440)
);

NOR4xp75_ASAP7_75t_L g2441 ( 
.A(n_2434),
.B(n_2001),
.C(n_2028),
.D(n_1922),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2437),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2432),
.B(n_2118),
.Y(n_2443)
);

NAND3xp33_ASAP7_75t_SL g2444 ( 
.A(n_2433),
.B(n_2436),
.C(n_2437),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2439),
.B(n_2438),
.Y(n_2445)
);

NOR2xp67_ASAP7_75t_L g2446 ( 
.A(n_2442),
.B(n_2066),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2443),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2441),
.Y(n_2448)
);

OAI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2445),
.A2(n_2444),
.B(n_2440),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2449),
.A2(n_2445),
.B(n_2448),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2450),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2450),
.Y(n_2452)
);

OAI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2451),
.A2(n_2446),
.B(n_2447),
.Y(n_2453)
);

AOI221xp5_ASAP7_75t_L g2454 ( 
.A1(n_2452),
.A2(n_2178),
.B1(n_2118),
.B2(n_2151),
.C(n_2117),
.Y(n_2454)
);

AOI222xp33_ASAP7_75t_L g2455 ( 
.A1(n_2453),
.A2(n_2454),
.B1(n_2178),
.B2(n_2123),
.C1(n_2154),
.C2(n_2117),
.Y(n_2455)
);

AND2x2_ASAP7_75t_SL g2456 ( 
.A(n_2453),
.B(n_2024),
.Y(n_2456)
);

AOI322xp5_ASAP7_75t_L g2457 ( 
.A1(n_2456),
.A2(n_2116),
.A3(n_2154),
.B1(n_2128),
.B2(n_2132),
.C1(n_2137),
.C2(n_2145),
.Y(n_2457)
);

AOI221xp5_ASAP7_75t_L g2458 ( 
.A1(n_2457),
.A2(n_2455),
.B1(n_2132),
.B2(n_2145),
.C(n_2137),
.Y(n_2458)
);

AOI211xp5_ASAP7_75t_L g2459 ( 
.A1(n_2458),
.A2(n_2177),
.B(n_2168),
.C(n_2149),
.Y(n_2459)
);


endmodule