module fake_jpeg_4797_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx10_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_9),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_30),
.B(n_15),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_14),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.C(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_22),
.B1(n_5),
.B2(n_4),
.Y(n_34)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_24),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_39),
.C(n_8),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_8),
.C(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_8),
.B2(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_32),
.C(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_44),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_43),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_45),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B(n_48),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_25),
.C(n_21),
.Y(n_54)
);


endmodule