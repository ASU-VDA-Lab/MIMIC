module fake_jpeg_16511_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

AND2x4_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_51),
.B1(n_24),
.B2(n_22),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_62),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_36),
.C(n_37),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_68),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_39),
.B1(n_26),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_54),
.B1(n_31),
.B2(n_49),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_77),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_37),
.C(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_25),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_39),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_37),
.C(n_34),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_31),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_83),
.Y(n_122)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_57),
.B1(n_58),
.B2(n_20),
.C(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_39),
.B1(n_55),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_99),
.B1(n_101),
.B2(n_79),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_64),
.B(n_73),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_1),
.B(n_2),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_34),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_72),
.B(n_38),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_74),
.B1(n_80),
.B2(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_31),
.B1(n_53),
.B2(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_94),
.B1(n_89),
.B2(n_95),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_88),
.Y(n_133)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_62),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_120),
.B(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_25),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_24),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_102),
.C(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_129),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_115),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_125),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_133),
.B1(n_107),
.B2(n_103),
.C(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_95),
.B1(n_101),
.B2(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_1),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_99),
.B(n_82),
.C(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_140),
.C(n_110),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_93),
.B(n_21),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_104),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_21),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_111),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_155),
.C(n_131),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_122),
.C(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_156),
.B(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_116),
.C(n_109),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_163),
.B(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_155),
.C(n_151),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_133),
.B(n_123),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_127),
.B1(n_125),
.B2(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_23),
.B1(n_4),
.B2(n_2),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_132),
.B(n_134),
.C(n_135),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_144),
.B(n_146),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_109),
.C(n_113),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_29),
.C(n_23),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_177),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_146),
.B(n_109),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_23),
.C(n_3),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_159),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_175),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_178),
.B(n_9),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_170),
.C(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_192),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_169),
.B1(n_160),
.B2(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_9),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_186),
.B1(n_184),
.B2(n_4),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_10),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_11),
.C(n_12),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_195),
.C(n_199),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_11),
.Y(n_206)
);


endmodule