module real_jpeg_4376_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_8;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

INVx13_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

A2O1A1Ixp33_ASAP7_75t_L g3 ( 
.A1(n_1),
.A2(n_4),
.B(n_7),
.C(n_10),
.Y(n_3)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_8),
.Y(n_7)
);

INVx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx13_ASAP7_75t_L g4 ( 
.A(n_5),
.Y(n_4)
);

INVx8_ASAP7_75t_L g5 ( 
.A(n_6),
.Y(n_5)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);


endmodule