module fake_netlist_6_725_n_109 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_109);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_109;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

AND2x6_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_17),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_24),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_19),
.B1(n_30),
.B2(n_29),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_20),
.C(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_42),
.B1(n_41),
.B2(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_33),
.B(n_34),
.Y(n_54)
);

OAI22x1_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_32),
.Y(n_56)
);

AOI221xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_32),
.B1(n_2),
.B2(n_4),
.C(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_33),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_33),
.B(n_14),
.Y(n_59)
);

AO21x2_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_49),
.B(n_48),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_44),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_49),
.B(n_48),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_45),
.B(n_33),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_44),
.B(n_46),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_61),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_66),
.B(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AO31x2_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_60),
.A3(n_66),
.B(n_65),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_65),
.B(n_61),
.C(n_66),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_73),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.Y(n_86)
);

NAND4xp25_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_69),
.C(n_76),
.D(n_6),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp67_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_80),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_69),
.B1(n_85),
.B2(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_84),
.B1(n_80),
.B2(n_72),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI211xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_46),
.B(n_4),
.C(n_7),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_93),
.C(n_92),
.Y(n_96)
);

AOI222xp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_90),
.B1(n_45),
.B2(n_92),
.C1(n_10),
.C2(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_47),
.Y(n_98)
);

OAI211xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_1),
.B(n_8),
.C(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_72),
.B1(n_75),
.B2(n_64),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_75),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_100),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_102),
.B1(n_60),
.B2(n_47),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_105),
.B1(n_60),
.B2(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_47),
.B1(n_60),
.B2(n_64),
.Y(n_109)
);


endmodule