module fake_jpeg_11476_n_613 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_62),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_68),
.A2(n_22),
.B1(n_54),
.B2(n_29),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_8),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_75),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_87),
.Y(n_127)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_28),
.B(n_6),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_112),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_108),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_24),
.B(n_10),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_118),
.Y(n_167)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_37),
.A2(n_11),
.B(n_13),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_17),
.B(n_37),
.Y(n_143)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_42),
.B(n_49),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_29),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_137),
.B(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_32),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_142),
.B(n_186),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_36),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_79),
.A2(n_37),
.B1(n_55),
.B2(n_38),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_156),
.A2(n_183),
.B(n_48),
.Y(n_238)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_58),
.B(n_32),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_95),
.Y(n_171)
);

CKINVDCx6p67_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_179),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_59),
.A2(n_55),
.B1(n_35),
.B2(n_34),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_175),
.A2(n_75),
.B1(n_82),
.B2(n_88),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_99),
.A2(n_20),
.B1(n_37),
.B2(n_51),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_194),
.B1(n_68),
.B2(n_122),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_58),
.B(n_47),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_184),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_20),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_56),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_62),
.B(n_56),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_22),
.B1(n_45),
.B2(n_27),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_63),
.B(n_45),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_65),
.Y(n_191)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_95),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_102),
.A2(n_37),
.B1(n_55),
.B2(n_38),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_80),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_205),
.A2(n_206),
.B1(n_262),
.B2(n_158),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_86),
.B1(n_76),
.B2(n_81),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_226),
.Y(n_288)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_215),
.B(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_218),
.A2(n_241),
.B(n_185),
.Y(n_304)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_219),
.Y(n_315)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_117),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_140),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_225),
.B(n_229),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_168),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_201),
.B1(n_197),
.B2(n_196),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_228),
.A2(n_127),
.B1(n_165),
.B2(n_198),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_49),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_128),
.Y(n_230)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_152),
.A2(n_46),
.B1(n_60),
.B2(n_96),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_149),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_233),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_140),
.B(n_46),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_240),
.Y(n_291)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_250),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_137),
.B(n_18),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_170),
.B(n_18),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_175),
.A2(n_85),
.B1(n_109),
.B2(n_104),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_242),
.A2(n_243),
.B1(n_253),
.B2(n_261),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_120),
.B1(n_103),
.B2(n_54),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_202),
.Y(n_244)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_251),
.Y(n_293)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_152),
.A2(n_27),
.B1(n_55),
.B2(n_38),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_263),
.B1(n_272),
.B2(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_129),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g252 ( 
.A(n_154),
.Y(n_252)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_150),
.A2(n_134),
.B1(n_139),
.B2(n_148),
.Y(n_253)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

CKINVDCx9p33_ASAP7_75t_R g323 ( 
.A(n_254),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_0),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_123),
.B(n_0),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_258),
.Y(n_331)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_129),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_151),
.A2(n_176),
.B1(n_166),
.B2(n_38),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_178),
.A2(n_35),
.B1(n_51),
.B2(n_43),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_159),
.A2(n_35),
.B1(n_51),
.B2(n_43),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_181),
.Y(n_265)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_125),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_270),
.Y(n_297)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_124),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_133),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_3),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_159),
.A2(n_35),
.B1(n_51),
.B2(n_43),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_138),
.B1(n_136),
.B2(n_169),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_207),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_330),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_287),
.B1(n_321),
.B2(n_322),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_157),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_313),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_285),
.A2(n_289),
.B1(n_305),
.B2(n_310),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_227),
.A2(n_242),
.B1(n_221),
.B2(n_228),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_292),
.Y(n_336)
);

OR2x4_ASAP7_75t_L g302 ( 
.A(n_218),
.B(n_127),
.Y(n_302)
);

HAxp5_ASAP7_75t_SL g348 ( 
.A(n_302),
.B(n_254),
.CON(n_348),
.SN(n_348)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_214),
.B(n_157),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_303),
.B(n_307),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_218),
.A2(n_187),
.B1(n_177),
.B2(n_160),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_204),
.B(n_132),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_221),
.A2(n_213),
.B1(n_219),
.B2(n_208),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_236),
.B(n_135),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_237),
.B(n_173),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_320),
.B(n_244),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_237),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_240),
.A2(n_144),
.B1(n_43),
.B2(n_153),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_268),
.A2(n_48),
.B1(n_11),
.B2(n_14),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_323),
.B1(n_267),
.B2(n_259),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_217),
.B(n_3),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_4),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_211),
.B(n_216),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_285),
.A2(n_265),
.B1(n_250),
.B2(n_239),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_364),
.B1(n_325),
.B2(n_322),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_323),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_334),
.B(n_337),
.Y(n_389)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_280),
.A2(n_241),
.B(n_271),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_338),
.A2(n_350),
.B(n_297),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_286),
.Y(n_341)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_223),
.C(n_220),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_370),
.C(n_361),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_352),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_293),
.C(n_291),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_296),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_353),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_275),
.A2(n_211),
.B(n_222),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_233),
.B1(n_244),
.B2(n_248),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_351),
.A2(n_355),
.B1(n_358),
.B2(n_368),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_211),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_286),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_304),
.A2(n_211),
.B(n_231),
.C(n_252),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_362),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_312),
.A2(n_246),
.B1(n_203),
.B2(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_321),
.A2(n_210),
.B1(n_203),
.B2(n_230),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_319),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_359),
.B(n_325),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_280),
.B(n_252),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_361),
.B(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_264),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_363),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_281),
.A2(n_305),
.B1(n_313),
.B2(n_275),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_247),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_369),
.Y(n_384)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_280),
.A2(n_269),
.B1(n_270),
.B2(n_234),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_278),
.B(n_209),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_224),
.C(n_272),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_278),
.B(n_326),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_372),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_279),
.B(n_258),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_326),
.B(n_274),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_315),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_287),
.A2(n_48),
.B1(n_52),
.B2(n_11),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_375),
.A2(n_315),
.B1(n_309),
.B2(n_316),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_371),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_345),
.A2(n_288),
.B1(n_282),
.B2(n_283),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_398),
.B1(n_401),
.B2(n_392),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_391),
.C(n_393),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_407),
.B1(n_412),
.B2(n_352),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_298),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_302),
.Y(n_393)
);

AOI21x1_ASAP7_75t_SL g428 ( 
.A1(n_394),
.A2(n_410),
.B(n_354),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_404),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_345),
.A2(n_282),
.B1(n_315),
.B2(n_299),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_319),
.C(n_316),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_403),
.C(n_373),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_409),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_319),
.C(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_406),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_282),
.B1(n_311),
.B2(n_317),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_350),
.A2(n_309),
.B(n_290),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_336),
.B(n_353),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_317),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_338),
.A2(n_306),
.B(n_314),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_354),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_372),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_349),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_380),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_413),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_387),
.A2(n_351),
.B1(n_358),
.B2(n_355),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_429),
.B1(n_431),
.B2(n_435),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_416),
.Y(n_464)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_419),
.B(n_335),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_422),
.A2(n_437),
.B1(n_444),
.B2(n_446),
.Y(n_467)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_426),
.Y(n_463)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_440),
.B(n_408),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_359),
.B1(n_360),
.B2(n_362),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_343),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_430),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_411),
.A2(n_364),
.B1(n_373),
.B2(n_346),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_434),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_391),
.B(n_344),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_390),
.B(n_344),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_376),
.B(n_341),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_393),
.B(n_365),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_441),
.C(n_442),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_410),
.B(n_380),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_386),
.B(n_373),
.C(n_366),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_347),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_447),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_390),
.B(n_343),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_357),
.B(n_332),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_445),
.A2(n_389),
.B(n_384),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_374),
.B1(n_334),
.B2(n_340),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_367),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_448),
.A2(n_452),
.B(n_472),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_449),
.B(n_473),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_422),
.A2(n_388),
.B1(n_398),
.B2(n_379),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_453),
.A2(n_415),
.B1(n_445),
.B2(n_446),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_399),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_456),
.B(n_476),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_429),
.A2(n_388),
.B1(n_379),
.B2(n_402),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_458),
.A2(n_459),
.B1(n_469),
.B2(n_417),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_413),
.A2(n_406),
.B1(n_400),
.B2(n_403),
.Y(n_459)
);

AO22x1_ASAP7_75t_L g462 ( 
.A1(n_440),
.A2(n_400),
.B1(n_381),
.B2(n_405),
.Y(n_462)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_425),
.C(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_474),
.C(n_478),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_381),
.B1(n_405),
.B2(n_377),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_306),
.C(n_301),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_290),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_341),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_301),
.C(n_300),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_421),
.B(n_420),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_428),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_449),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_468),
.B(n_443),
.Y(n_482)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_483),
.A2(n_486),
.B1(n_494),
.B2(n_497),
.Y(n_512)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_438),
.B1(n_418),
.B2(n_427),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_493),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_466),
.Y(n_488)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_448),
.A2(n_458),
.B(n_450),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_489),
.A2(n_462),
.B(n_463),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_363),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_455),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_453),
.A2(n_414),
.B1(n_424),
.B2(n_426),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_455),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_501),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_496),
.A2(n_294),
.B1(n_328),
.B2(n_311),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_452),
.A2(n_414),
.B1(n_432),
.B2(n_434),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_468),
.B(n_423),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_498),
.A2(n_499),
.B1(n_450),
.B2(n_461),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_477),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_460),
.C(n_456),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_460),
.C(n_474),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_502),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_340),
.Y(n_503)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_363),
.Y(n_504)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_457),
.B(n_329),
.Y(n_506)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_506),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_513),
.B(n_485),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_515),
.C(n_516),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_469),
.C(n_473),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_476),
.C(n_459),
.Y(n_516)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_462),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_529),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_494),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_475),
.C(n_454),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_532),
.C(n_495),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_329),
.Y(n_525)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_525),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_527),
.A2(n_496),
.B1(n_486),
.B2(n_497),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_284),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_501),
.B(n_284),
.C(n_300),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_546),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_528),
.Y(n_538)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_538),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_524),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_539),
.B(n_543),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_514),
.B(n_480),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_541),
.Y(n_555)
);

FAx1_ASAP7_75t_SL g541 ( 
.A(n_516),
.B(n_505),
.CI(n_481),
.CON(n_541),
.SN(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_530),
.A2(n_484),
.B1(n_490),
.B2(n_493),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_520),
.B1(n_531),
.B2(n_508),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_489),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_544),
.B(n_549),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_545),
.A2(n_552),
.B1(n_536),
.B2(n_522),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_487),
.C(n_505),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_510),
.C(n_532),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_510),
.Y(n_563)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_517),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_485),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_550),
.B(n_551),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_483),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_512),
.B(n_503),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_552),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_534),
.A2(n_523),
.B(n_509),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_556),
.A2(n_561),
.B(n_277),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_557),
.B(n_565),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_535),
.B(n_539),
.C(n_546),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_566),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_548),
.A2(n_509),
.B(n_508),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_567),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_535),
.B(n_511),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_543),
.B(n_522),
.C(n_520),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_537),
.Y(n_567)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_568),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_506),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_547),
.C(n_541),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_574),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_556),
.A2(n_531),
.B(n_525),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_572),
.A2(n_581),
.B(n_561),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_518),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_518),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_575),
.B(n_577),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_331),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_566),
.B(n_331),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_557),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_568),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_572),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_587),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_564),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_591),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_580),
.B(n_560),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_589),
.B(n_590),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_555),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_564),
.B(n_578),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_592),
.A2(n_578),
.B(n_585),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_594),
.B(n_598),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_591),
.A2(n_554),
.B(n_563),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_596),
.A2(n_290),
.B(n_276),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_554),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_567),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_599),
.B(n_588),
.Y(n_601)
);

OAI21x1_ASAP7_75t_SL g604 ( 
.A1(n_601),
.A2(n_602),
.B(n_603),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_593),
.A2(n_277),
.B1(n_328),
.B2(n_276),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_600),
.A2(n_597),
.B(n_595),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_605),
.B(n_4),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g606 ( 
.A(n_600),
.B(n_4),
.C(n_5),
.Y(n_606)
);

O2A1O1Ixp5_ASAP7_75t_L g608 ( 
.A1(n_606),
.A2(n_4),
.B(n_5),
.C(n_52),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_607),
.B(n_608),
.C(n_5),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_609),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_604),
.C(n_52),
.Y(n_611)
);

BUFx24_ASAP7_75t_SL g612 ( 
.A(n_611),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_SL g613 ( 
.A(n_612),
.B(n_5),
.C(n_52),
.Y(n_613)
);


endmodule