module fake_jpeg_3623_n_167 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_15),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_73),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_60),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_62),
.B1(n_60),
.B2(n_56),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_62),
.B1(n_59),
.B2(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_87),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_57),
.B1(n_46),
.B2(n_44),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_44),
.Y(n_98)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_50),
.B1(n_46),
.B2(n_49),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_52),
.C(n_48),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_43),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_52),
.B(n_49),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_68),
.C(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_40),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_97),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_63),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AND2x4_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_68),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_5),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_23),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_86),
.B1(n_84),
.B2(n_8),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_115),
.Y(n_137)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_7),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_99),
.B1(n_90),
.B2(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_6),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_24),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_22),
.B1(n_38),
.B2(n_37),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_90),
.B(n_21),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_129),
.B(n_26),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_18),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_136),
.C(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_132),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_120),
.B(n_116),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_134),
.B1(n_138),
.B2(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_7),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_127),
.B1(n_133),
.B2(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_25),
.C(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_142),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_27),
.C(n_34),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_146),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_39),
.C(n_33),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_29),
.B1(n_32),
.B2(n_14),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_16),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_129),
.B1(n_137),
.B2(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_13),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_155),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_152),
.B(n_16),
.C(n_17),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_17),
.Y(n_167)
);


endmodule