module real_jpeg_7589_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_0),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_0),
.B(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_2),
.B(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_4),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_7),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_13),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_13),
.B(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_122),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_120),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_104),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_17),
.B(n_104),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_61),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_46),
.B2(n_47),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.C(n_37),
.Y(n_20)
);

FAx1_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_33),
.CI(n_37),
.CON(n_105),
.SN(n_105)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_22),
.Y(n_137)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_24),
.Y(n_135)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_24),
.Y(n_157)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_35),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_77),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_73),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B1(n_102),
.B2(n_103),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_98),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.C(n_118),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_176),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_105),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.C(n_116),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_116),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_173),
.B(n_177),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_149),
.B(n_172),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_138),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_138),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_129),
.C(n_136),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_133),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_144),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_166),
.B(n_171),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_159),
.B(n_165),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_158),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_156),
.Y(n_167)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);


endmodule