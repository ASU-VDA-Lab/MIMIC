module real_jpeg_27803_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_262, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_262;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_16),
.B1(n_53),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_16),
.B1(n_43),
.B2(n_44),
.Y(n_203)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_1),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_5),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_22),
.B(n_26),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_5),
.B(n_29),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_5),
.A2(n_6),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_8),
.B(n_25),
.C(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_9),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_184)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_10),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_254),
.B(n_257),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_66),
.B(n_253),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_30),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_14),
.B(n_30),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_14),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_19),
.B1(n_27),
.B2(n_29),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_15),
.A2(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_17),
.A2(n_23),
.B(n_34),
.C(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_45),
.Y(n_46)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_27),
.B(n_35),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_61),
.C(n_62),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_31),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.C(n_48),
.Y(n_31)
);

AOI211xp5_ASAP7_75t_L g75 ( 
.A1(n_32),
.A2(n_76),
.B(n_78),
.C(n_83),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_32),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_32),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_32),
.A2(n_84),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_32),
.A2(n_84),
.B1(n_198),
.B2(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_32),
.A2(n_84),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_32),
.A2(n_198),
.B(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_32),
.A2(n_84),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_32),
.A2(n_84),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_32),
.B(n_48),
.C(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_32),
.B(n_240),
.C(n_241),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_34),
.A2(n_44),
.B(n_56),
.C(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_34),
.B(n_52),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_34),
.B(n_137),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_34),
.A2(n_43),
.B(n_45),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_36),
.A2(n_48),
.B1(n_49),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_36),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_38),
.A2(n_81),
.B1(n_128),
.B2(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_48),
.A2(n_49),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_52),
.A2(n_57),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_52),
.A2(n_57),
.B1(n_60),
.B2(n_203),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_53),
.B(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_61),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_247),
.B(n_252),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_225),
.A3(n_242),
.B1(n_245),
.B2(n_246),
.C(n_262),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_209),
.B(n_224),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_190),
.B(n_208),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_115),
.B(n_172),
.C(n_189),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_105),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_72),
.B(n_105),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_94),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_85),
.B2(n_86),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_74),
.B(n_86),
.C(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_82),
.B1(n_87),
.B2(n_93),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_82),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_76),
.A2(n_82),
.B1(n_122),
.B2(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_101),
.C(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_76),
.A2(n_82),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_155),
.C(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_76),
.B(n_87),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_76),
.A2(n_82),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_76),
.B(n_181),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_84),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_79),
.A2(n_82),
.B(n_149),
.C(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_79),
.A2(n_80),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_79),
.B(n_84),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_101),
.C(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_80),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_80),
.B(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_83),
.A2(n_104),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_88),
.A2(n_92),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_104),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_95),
.A2(n_96),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_95),
.A2(n_96),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_102),
.B1(n_125),
.B2(n_129),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_102),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_102),
.B1(n_113),
.B2(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_139),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_107),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_109),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_171),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_164),
.B(n_170),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_151),
.B(n_163),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_142),
.B(n_150),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_130),
.B(n_141),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_174),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_179),
.B1(n_185),
.B2(n_186),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_185),
.C(n_187),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_192),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_205),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_197),
.C(n_205),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_195),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_206),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_204),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_201),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.C(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_227),
.C(n_233),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_227),
.CI(n_233),
.CON(n_244),
.SN(n_244)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);


endmodule