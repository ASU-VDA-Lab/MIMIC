module real_jpeg_12806_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_311, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_311;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_3),
.A2(n_38),
.B1(n_44),
.B2(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_38),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_38),
.B1(n_149),
.B2(n_161),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_7),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_7),
.A2(n_44),
.B1(n_47),
.B2(n_153),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_7),
.A2(n_101),
.B1(n_102),
.B2(n_153),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_7),
.A2(n_149),
.B1(n_153),
.B2(n_161),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_46),
.B1(n_101),
.B2(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_9),
.A2(n_46),
.B1(n_149),
.B2(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_30),
.C(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_31),
.B1(n_44),
.B2(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_10),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_48),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_31),
.B1(n_101),
.B2(n_102),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_58),
.B(n_102),
.C(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_31),
.B1(n_149),
.B2(n_161),
.Y(n_166)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_248),
.C(n_304),
.Y(n_12)
);

OA21x2_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_303),
.B(n_308),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_295),
.B(n_302),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_257),
.B(n_292),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_238),
.B(n_256),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_217),
.B(n_237),
.Y(n_17)
);

AOI321xp33_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_177),
.A3(n_210),
.B1(n_215),
.B2(n_216),
.C(n_311),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_140),
.B(n_176),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_117),
.B(n_139),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_94),
.B(n_116),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_72),
.B(n_93),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_26),
.B(n_90),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_36),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_28),
.A2(n_33),
.B(n_36),
.Y(n_112)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_30),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_47),
.B(n_59),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_31),
.B(n_102),
.C(n_130),
.Y(n_148)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_33),
.A2(n_90),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_36),
.A2(n_152),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_42),
.B(n_69),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_42),
.A2(n_174),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_43),
.B(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_48),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_48),
.Y(n_175)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_51),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_52),
.Y(n_174)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_60),
.C(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_56),
.B(n_107),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_56),
.A2(n_104),
.B(n_107),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_56),
.A2(n_170),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_59),
.B1(n_101),
.B2(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_71),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_86),
.B(n_92),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_80),
.B(n_85),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_108),
.C(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_102),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_103),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_105),
.B(n_134),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_105),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_109),
.A2(n_175),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_109),
.B(n_121),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_111),
.A2(n_112),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_111),
.A2(n_112),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_112),
.B(n_234),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_112),
.A2(n_245),
.B(n_247),
.Y(n_261)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_138),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_138),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_137),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_126),
.B(n_145),
.C(n_155),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.CI(n_132),
.CON(n_126),
.SN(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_129),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_129),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_131),
.B1(n_149),
.B2(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_133),
.B(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_142),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_156),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_154),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_169),
.C(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_164),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_162),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_163),
.A2(n_166),
.B(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_163),
.A2(n_181),
.B(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_182),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_170),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_172),
.A2(n_173),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_172),
.A2(n_173),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_173),
.B(n_265),
.C(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_173),
.B(n_289),
.C(n_291),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_204),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_204),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_189),
.C(n_200),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_187),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_181),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_185),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_200),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_197),
.C(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_196),
.A2(n_249),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_196),
.B(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_197),
.A2(n_199),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_300),
.C(n_301),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_219),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_236),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_232),
.B2(n_233),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_233),
.C(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_225),
.C(n_230),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_243),
.C(n_251),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B(n_255),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_263),
.B1(n_264),
.B2(n_274),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_261),
.C(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_275),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_266),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_278),
.C(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_297),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_307),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);


endmodule