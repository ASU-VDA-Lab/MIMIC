module fake_netlist_1_11717_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx3_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OAI21x1_ASAP7_75t_L g12 ( .A1(n_1), .A2(n_5), .B(n_3), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_2), .B(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
NOR3xp33_ASAP7_75t_SL g17 ( .A(n_15), .B(n_0), .C(n_1), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_10), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_16), .A2(n_12), .B(n_11), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_14), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
O2A1O1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_18), .B(n_17), .C(n_20), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
OA22x2_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_21), .B1(n_12), .B2(n_14), .Y(n_30) );
AOI21xp5_ASAP7_75t_SL g31 ( .A1(n_28), .A2(n_10), .B(n_18), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_19), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_13), .Y(n_33) );
NAND3x2_ASAP7_75t_L g34 ( .A(n_30), .B(n_2), .C(n_4), .Y(n_34) );
NAND3xp33_ASAP7_75t_L g35 ( .A(n_34), .B(n_30), .C(n_21), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
XOR2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_33), .Y(n_37) );
AOI22xp33_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_35), .B1(n_6), .B2(n_9), .Y(n_38) );
endmodule