module real_aes_9087_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_0), .A2(n_160), .B(n_472), .C(n_475), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_1), .B(n_466), .Y(n_476) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_2), .B(n_88), .C(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
INVx1_ASAP7_75t_L g158 ( .A(n_3), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_4), .B(n_161), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_5), .A2(n_461), .B(n_534), .Y(n_533) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_6), .A2(n_183), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_7), .A2(n_39), .B1(n_148), .B2(n_206), .Y(n_246) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_8), .A2(n_20), .B1(n_436), .B2(n_722), .C1(n_723), .C2(n_726), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_8), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_9), .B(n_183), .Y(n_191) );
AND2x6_ASAP7_75t_L g163 ( .A(n_10), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_11), .A2(n_163), .B(n_452), .C(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_12), .B(n_40), .Y(n_104) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_15), .B(n_144), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_16), .B(n_161), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_17), .B(n_135), .Y(n_193) );
AO32x2_ASAP7_75t_L g244 ( .A1(n_18), .A2(n_134), .A3(n_177), .B1(n_183), .B2(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_19), .A2(n_30), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_19), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_21), .B(n_148), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_22), .B(n_135), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_23), .A2(n_54), .B1(n_148), .B2(n_206), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g208 ( .A1(n_24), .A2(n_80), .B1(n_144), .B2(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_25), .B(n_148), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_26), .A2(n_177), .B(n_452), .C(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_27), .A2(n_177), .B(n_452), .C(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_28), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_29), .B(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_30), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_30), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_31), .A2(n_461), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_32), .B(n_179), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_33), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_35), .A2(n_458), .B(n_501), .C(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_36), .B(n_148), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_37), .B(n_179), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_38), .B(n_228), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_41), .B(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_42), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_43), .B(n_161), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_44), .B(n_461), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_45), .A2(n_458), .B(n_501), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_46), .B(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g473 ( .A(n_47), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_48), .A2(n_89), .B1(n_206), .B2(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g526 ( .A(n_49), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_50), .B(n_148), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_51), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_52), .B(n_461), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_53), .B(n_156), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g197 ( .A1(n_55), .A2(n_59), .B1(n_144), .B2(n_148), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_56), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_57), .B(n_148), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_58), .B(n_148), .Y(n_225) );
INVx1_ASAP7_75t_L g164 ( .A(n_60), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_61), .A2(n_101), .B1(n_110), .B2(n_730), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_62), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_63), .B(n_466), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_64), .A2(n_150), .B(n_156), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_65), .B(n_148), .Y(n_159) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_67), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_68), .B(n_161), .Y(n_504) );
AO32x2_ASAP7_75t_L g203 ( .A1(n_69), .A2(n_177), .A3(n_183), .B1(n_204), .B2(n_209), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_70), .B(n_162), .Y(n_517) );
INVx1_ASAP7_75t_L g173 ( .A(n_71), .Y(n_173) );
INVx1_ASAP7_75t_L g216 ( .A(n_72), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_73), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_74), .B(n_485), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_75), .A2(n_452), .B(n_454), .C(n_458), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_76), .B(n_144), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_77), .Y(n_535) );
INVx1_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_79), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_81), .B(n_206), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_82), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_83), .B(n_144), .Y(n_220) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_85), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_86), .B(n_176), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_87), .B(n_144), .Y(n_187) );
OR2x2_ASAP7_75t_L g118 ( .A(n_88), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g439 ( .A(n_88), .B(n_120), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_88), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_90), .A2(n_99), .B1(n_144), .B2(n_145), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_91), .B(n_461), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_92), .Y(n_503) );
INVxp67_ASAP7_75t_L g538 ( .A(n_93), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_94), .B(n_144), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_95), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g455 ( .A(n_96), .Y(n_455) );
INVx1_ASAP7_75t_L g513 ( .A(n_97), .Y(n_513) );
AND2x2_ASAP7_75t_L g528 ( .A(n_98), .B(n_179), .Y(n_528) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g732 ( .A(n_103), .Y(n_732) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g120 ( .A(n_104), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_116), .B(n_434), .Y(n_110) );
BUFx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g729 ( .A(n_115), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_431), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g433 ( .A(n_118), .Y(n_433) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_119), .B(n_443), .Y(n_725) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g442 ( .A(n_120), .B(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_127), .B2(n_430), .Y(n_122) );
INVx1_ASAP7_75t_L g430 ( .A(n_123), .Y(n_430) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR5x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_321), .C(n_379), .D(n_415), .E(n_422), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_267), .C(n_291), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_199), .B1(n_233), .B2(n_238), .C(n_248), .Y(n_129) );
OAI21xp5_ASAP7_75t_SL g401 ( .A1(n_130), .A2(n_402), .B(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_180), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_131), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
INVx2_ASAP7_75t_L g237 ( .A(n_132), .Y(n_237) );
AND2x2_ASAP7_75t_L g250 ( .A(n_132), .B(n_182), .Y(n_250) );
AND2x2_ASAP7_75t_L g304 ( .A(n_132), .B(n_181), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_132), .B(n_167), .Y(n_319) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_165), .Y(n_132) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_133), .A2(n_168), .B(n_178), .Y(n_167) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_134), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_136), .B(n_137), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_154), .B(n_163), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_147), .C(n_150), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_143), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_143), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx3_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_148), .Y(n_457) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
AND2x6_ASAP7_75t_L g452 ( .A(n_149), .B(n_453), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_150), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_151), .A2(n_219), .B(n_220), .Y(n_218) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g485 ( .A(n_152), .Y(n_485) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
INVx1_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g453 ( .A(n_153), .Y(n_453) );
AND2x2_ASAP7_75t_L g462 ( .A(n_153), .B(n_157), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_159), .C(n_160), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g172 ( .A1(n_155), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_155), .A2(n_484), .B(n_486), .Y(n_483) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_189), .B(n_190), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_176), .B1(n_196), .B2(n_197), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_160), .A2(n_176), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_161), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_186), .B(n_187), .Y(n_185) );
O2A1O1Ixp5_ASAP7_75t_SL g214 ( .A1(n_161), .A2(n_215), .B(n_216), .C(n_217), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_161), .B(n_538), .Y(n_537) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_162), .A2(n_176), .B1(n_205), .B2(n_208), .Y(n_204) );
BUFx3_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_163), .A2(n_185), .B(n_188), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_163), .A2(n_214), .B(n_218), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_163), .A2(n_224), .B(n_229), .Y(n_223) );
INVx4_ASAP7_75t_SL g459 ( .A(n_163), .Y(n_459) );
AND2x4_ASAP7_75t_L g461 ( .A(n_163), .B(n_462), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_163), .B(n_462), .Y(n_514) );
AND2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_278), .Y(n_337) );
AND2x2_ASAP7_75t_L g370 ( .A(n_166), .B(n_182), .Y(n_370) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g277 ( .A(n_167), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g290 ( .A(n_167), .B(n_182), .Y(n_290) );
AND2x2_ASAP7_75t_L g297 ( .A(n_167), .B(n_278), .Y(n_297) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_167), .Y(n_306) );
AND2x2_ASAP7_75t_L g313 ( .A(n_167), .B(n_181), .Y(n_313) );
INVx1_ASAP7_75t_L g344 ( .A(n_167), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_177), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_175), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g474 ( .A(n_176), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g194 ( .A(n_177), .B(n_195), .C(n_198), .Y(n_194) );
INVx2_ASAP7_75t_L g209 ( .A(n_179), .Y(n_209) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_179), .A2(n_213), .B(n_221), .Y(n_212) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_179), .A2(n_223), .B(n_232), .Y(n_222) );
INVx1_ASAP7_75t_L g491 ( .A(n_179), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_179), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_179), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g320 ( .A(n_180), .Y(n_320) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_192), .Y(n_180) );
INVx2_ASAP7_75t_L g276 ( .A(n_181), .Y(n_276) );
AND2x2_ASAP7_75t_L g298 ( .A(n_181), .B(n_237), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_181), .B(n_344), .Y(n_349) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_182), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g421 ( .A(n_182), .B(n_385), .Y(n_421) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_191), .Y(n_182) );
INVx4_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_183), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_183), .A2(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g235 ( .A(n_192), .Y(n_235) );
INVx3_ASAP7_75t_L g336 ( .A(n_192), .Y(n_336) );
OR2x2_ASAP7_75t_L g366 ( .A(n_192), .B(n_367), .Y(n_366) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_192), .B(n_276), .Y(n_392) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
INVx1_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
AO21x1_ASAP7_75t_L g278 ( .A1(n_195), .A2(n_198), .B(n_279), .Y(n_278) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_198), .A2(n_450), .B(n_463), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_198), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g466 ( .A(n_198), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_198), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_198), .A2(n_512), .B(n_519), .Y(n_511) );
AOI33xp33_ASAP7_75t_L g412 ( .A1(n_199), .A2(n_250), .A3(n_264), .B1(n_336), .B2(n_413), .B3(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_210), .Y(n_200) );
OR2x2_ASAP7_75t_L g265 ( .A(n_201), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_201), .B(n_262), .Y(n_324) );
OR2x2_ASAP7_75t_L g377 ( .A(n_201), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g303 ( .A(n_202), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g328 ( .A(n_202), .B(n_210), .Y(n_328) );
AND2x2_ASAP7_75t_L g395 ( .A(n_202), .B(n_240), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_202), .A2(n_295), .B(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
AND2x2_ASAP7_75t_L g274 ( .A(n_203), .B(n_244), .Y(n_274) );
AND2x2_ASAP7_75t_L g323 ( .A(n_203), .B(n_243), .Y(n_323) );
INVx2_ASAP7_75t_L g475 ( .A(n_207), .Y(n_475) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_207), .Y(n_505) );
INVx1_ASAP7_75t_L g488 ( .A(n_209), .Y(n_488) );
INVx2_ASAP7_75t_SL g365 ( .A(n_210), .Y(n_365) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
INVx2_ASAP7_75t_L g285 ( .A(n_211), .Y(n_285) );
INVx1_ASAP7_75t_L g416 ( .A(n_211), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_211), .B(n_310), .Y(n_429) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
OR2x2_ASAP7_75t_L g262 ( .A(n_212), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_222), .Y(n_240) );
AND2x2_ASAP7_75t_L g257 ( .A(n_222), .B(n_243), .Y(n_257) );
INVx1_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
INVx1_ASAP7_75t_L g270 ( .A(n_222), .Y(n_270) );
AND2x2_ASAP7_75t_L g295 ( .A(n_222), .B(n_244), .Y(n_295) );
INVx2_ASAP7_75t_L g311 ( .A(n_222), .Y(n_311) );
AND2x2_ASAP7_75t_L g404 ( .A(n_222), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_222), .B(n_285), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g259 ( .A(n_235), .Y(n_259) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_235), .B(n_319), .Y(n_385) );
INVx1_ASAP7_75t_SL g345 ( .A(n_236), .Y(n_345) );
INVx2_ASAP7_75t_L g266 ( .A(n_237), .Y(n_266) );
AND2x2_ASAP7_75t_L g335 ( .A(n_237), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g351 ( .A(n_237), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g413 ( .A(n_239), .Y(n_413) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g268 ( .A(n_241), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g371 ( .A(n_241), .B(n_361), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_241), .A2(n_382), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
INVx1_ASAP7_75t_L g333 ( .A(n_242), .Y(n_333) );
OR2x2_ASAP7_75t_L g397 ( .A(n_243), .B(n_256), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_243), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g310 ( .A(n_244), .B(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_L g317 ( .A(n_244), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .B1(n_258), .B2(n_260), .Y(n_248) );
OR2x2_ASAP7_75t_L g327 ( .A(n_249), .B(n_277), .Y(n_327) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_250), .A2(n_369), .B1(n_371), .B2(n_372), .C1(n_373), .C2(n_376), .Y(n_368) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_257), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g315 ( .A(n_254), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_256), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_256), .Y(n_340) );
AND2x2_ASAP7_75t_L g388 ( .A(n_256), .B(n_257), .Y(n_388) );
INVx1_ASAP7_75t_L g406 ( .A(n_256), .Y(n_406) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g372 ( .A(n_259), .B(n_298), .Y(n_372) );
AND2x2_ASAP7_75t_L g414 ( .A(n_259), .B(n_290), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_261), .B(n_309), .Y(n_396) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_262), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g289 ( .A(n_266), .B(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g357 ( .A(n_266), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_275), .C(n_280), .Y(n_267) );
INVxp67_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_269), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_269), .B(n_316), .Y(n_411) );
BUFx3_ASAP7_75t_L g375 ( .A(n_270), .Y(n_375) );
INVx1_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g301 ( .A(n_273), .B(n_295), .Y(n_301) );
INVx1_ASAP7_75t_SL g341 ( .A(n_274), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g331 ( .A(n_276), .Y(n_331) );
AND2x2_ASAP7_75t_L g354 ( .A(n_276), .B(n_337), .Y(n_354) );
INVx1_ASAP7_75t_SL g325 ( .A(n_277), .Y(n_325) );
INVx1_ASAP7_75t_L g352 ( .A(n_278), .Y(n_352) );
AOI31xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .A3(n_283), .B(n_286), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g347 ( .A(n_285), .Y(n_347) );
BUFx2_ASAP7_75t_L g361 ( .A(n_285), .Y(n_361) );
AND2x2_ASAP7_75t_L g389 ( .A(n_285), .B(n_310), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g362 ( .A(n_289), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_290), .B(n_357), .Y(n_403) );
AND2x2_ASAP7_75t_L g410 ( .A(n_290), .B(n_336), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_296), .B(n_299), .C(n_314), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_296), .A2(n_323), .B1(n_324), .B2(n_325), .C(n_326), .Y(n_322) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g330 ( .A(n_297), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
OAI32xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_302), .A3(n_305), .B1(n_307), .B2(n_312), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_301), .A2(n_354), .B(n_355), .C(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OAI21xp5_ASAP7_75t_SL g417 ( .A1(n_309), .A2(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g378 ( .A(n_310), .Y(n_378) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_316), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g364 ( .A(n_316), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g381 ( .A(n_318), .Y(n_381) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND4xp25_ASAP7_75t_SL g321 ( .A(n_322), .B(n_334), .C(n_353), .D(n_368), .Y(n_321) );
AND2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g382 ( .A(n_323), .B(n_375), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_325), .B(n_357), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_329), .B2(n_332), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_327), .A2(n_378), .B1(n_409), .B2(n_411), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_327), .A2(n_416), .B(n_417), .C(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g386 ( .A(n_328), .Y(n_386) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_330), .A2(n_364), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_386), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_338), .C(n_342), .Y(n_334) );
INVx1_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_339), .A2(n_343), .B1(n_346), .B2(n_348), .Y(n_342) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g369 ( .A(n_351), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_363), .B2(n_366), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_361), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_372), .Y(n_426) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND5xp2_ASAP7_75t_L g379 ( .A(n_380), .B(n_387), .C(n_401), .D(n_407), .E(n_412), .Y(n_379) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_390), .C(n_393), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI31xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .A3(n_397), .B(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g422 ( .A1(n_409), .A2(n_411), .B1(n_423), .B2(n_426), .C1(n_427), .C2(n_428), .Y(n_422) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_431), .B(n_435), .C(n_729), .Y(n_434) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_441), .B2(n_444), .Y(n_437) );
INVx2_ASAP7_75t_L g727 ( .A(n_438), .Y(n_727) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_440), .A2(n_444), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g728 ( .A(n_441), .Y(n_728) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR3x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_630), .C(n_679), .Y(n_444) );
NAND5xp2_ASAP7_75t_L g445 ( .A(n_446), .B(n_564), .C(n_593), .D(n_601), .E(n_616), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_492), .B(n_508), .C(n_548), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_477), .Y(n_447) );
AND2x2_ASAP7_75t_L g559 ( .A(n_448), .B(n_556), .Y(n_559) );
AND2x2_ASAP7_75t_L g592 ( .A(n_448), .B(n_478), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_448), .B(n_496), .Y(n_685) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_465), .Y(n_448) );
INVx2_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
BUFx2_ASAP7_75t_L g659 ( .A(n_449), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx5_ASAP7_75t_L g470 ( .A(n_452), .Y(n_470) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_459), .A2(n_469), .B(n_470), .C(n_471), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_459), .A2(n_470), .B(n_535), .C(n_536), .Y(n_534) );
BUFx2_ASAP7_75t_L g481 ( .A(n_461), .Y(n_481) );
AND2x2_ASAP7_75t_L g477 ( .A(n_465), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g557 ( .A(n_465), .Y(n_557) );
AND2x2_ASAP7_75t_L g643 ( .A(n_465), .B(n_556), .Y(n_643) );
AND2x2_ASAP7_75t_L g698 ( .A(n_465), .B(n_495), .Y(n_698) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_476), .Y(n_465) );
INVx2_ASAP7_75t_L g501 ( .A(n_470), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g615 ( .A(n_477), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_477), .B(n_496), .Y(n_662) );
INVx5_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
AND2x4_ASAP7_75t_L g577 ( .A(n_478), .B(n_557), .Y(n_577) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_478), .Y(n_599) );
AND2x2_ASAP7_75t_L g674 ( .A(n_478), .B(n_659), .Y(n_674) );
AND2x2_ASAP7_75t_L g677 ( .A(n_478), .B(n_497), .Y(n_677) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
AOI21xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_488), .Y(n_479) );
INVx2_ASAP7_75t_L g487 ( .A(n_485), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_487), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_487), .A2(n_505), .B(n_526), .C(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_492), .B(n_557), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_492), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
AND2x2_ASAP7_75t_L g582 ( .A(n_494), .B(n_557), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_494), .B(n_497), .Y(n_600) );
INVx1_ASAP7_75t_L g620 ( .A(n_494), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_494), .B(n_556), .Y(n_665) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_494), .Y(n_707) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_496), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_496), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_496), .A2(n_552), .B(n_613), .C(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g628 ( .A(n_496), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g632 ( .A(n_496), .B(n_556), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_496), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_496), .B(n_557), .Y(n_647) );
AND2x2_ASAP7_75t_L g697 ( .A(n_496), .B(n_698), .Y(n_697) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g561 ( .A(n_497), .Y(n_561) );
AND2x2_ASAP7_75t_L g602 ( .A(n_497), .B(n_555), .Y(n_602) );
AND2x2_ASAP7_75t_L g614 ( .A(n_497), .B(n_589), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_497), .B(n_643), .Y(n_661) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_506), .Y(n_497) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_529), .Y(n_508) );
INVx1_ASAP7_75t_L g550 ( .A(n_509), .Y(n_550) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
OR2x2_ASAP7_75t_L g552 ( .A(n_510), .B(n_521), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_510), .B(n_559), .C(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_510), .B(n_531), .Y(n_569) );
OR2x2_ASAP7_75t_L g584 ( .A(n_510), .B(n_572), .Y(n_584) );
AND2x2_ASAP7_75t_L g590 ( .A(n_510), .B(n_540), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_510), .B(n_721), .Y(n_720) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_511), .B(n_531), .Y(n_587) );
AND2x2_ASAP7_75t_L g626 ( .A(n_511), .B(n_541), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_511), .B(n_540), .Y(n_654) );
OR2x2_ASAP7_75t_L g657 ( .A(n_511), .B(n_540), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
INVx5_ASAP7_75t_SL g572 ( .A(n_521), .Y(n_572) );
OR2x2_ASAP7_75t_L g578 ( .A(n_521), .B(n_530), .Y(n_578) );
AND2x2_ASAP7_75t_L g594 ( .A(n_521), .B(n_595), .Y(n_594) );
AOI321xp33_ASAP7_75t_L g601 ( .A1(n_521), .A2(n_602), .A3(n_603), .B1(n_604), .B2(n_610), .C(n_612), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_521), .B(n_529), .Y(n_611) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
OR2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_569), .Y(n_671) );
AND2x2_ASAP7_75t_L g693 ( .A(n_521), .B(n_590), .Y(n_693) );
AND2x2_ASAP7_75t_L g712 ( .A(n_521), .B(n_531), .Y(n_712) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_531), .B(n_540), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_531), .B(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g589 ( .A(n_531), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_531), .B(n_590), .Y(n_595) );
INVxp67_ASAP7_75t_L g625 ( .A(n_531), .Y(n_625) );
OR2x2_ASAP7_75t_L g667 ( .A(n_531), .B(n_572), .Y(n_667) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_531) );
OR2x2_ASAP7_75t_L g549 ( .A(n_540), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_SL g563 ( .A(n_540), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_540), .B(n_552), .Y(n_596) );
AND2x2_ASAP7_75t_L g645 ( .A(n_540), .B(n_589), .Y(n_645) );
AND2x2_ASAP7_75t_L g683 ( .A(n_540), .B(n_572), .Y(n_683) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_541), .B(n_572), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B(n_554), .C(n_558), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_549), .A2(n_551), .B1(n_676), .B2(n_678), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_551), .A2(n_574), .B1(n_629), .B2(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_SL g703 ( .A(n_552), .Y(n_703) );
INVx1_ASAP7_75t_SL g603 ( .A(n_553), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_555), .B(n_575), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_555), .A2(n_596), .B1(n_603), .B2(n_617), .C1(n_621), .C2(n_627), .Y(n_616) );
AND2x2_ASAP7_75t_L g706 ( .A(n_555), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g581 ( .A(n_556), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_556), .B(n_576), .Y(n_651) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_556), .Y(n_688) );
AND2x2_ASAP7_75t_L g691 ( .A(n_556), .B(n_600), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_556), .B(n_707), .Y(n_717) );
INVx1_ASAP7_75t_L g608 ( .A(n_557), .Y(n_608) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_557), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_559), .A2(n_700), .B(n_701), .C(n_704), .Y(n_699) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_561), .B(n_623), .C(n_626), .Y(n_622) );
OR2x2_ASAP7_75t_L g650 ( .A(n_561), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_561), .B(n_577), .Y(n_678) );
OR2x2_ASAP7_75t_L g583 ( .A(n_563), .B(n_584), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B(n_573), .C(n_585), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_566), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g672 ( .A(n_567), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_568), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g586 ( .A(n_571), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_572), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g640 ( .A(n_572), .B(n_590), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_572), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_572), .B(n_589), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .B1(n_579), .B2(n_583), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_575), .B(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_577), .B(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_578), .A2(n_642), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_641) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g696 ( .A(n_581), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_581), .B(n_698), .Y(n_709) );
INVx1_ASAP7_75t_L g629 ( .A(n_582), .Y(n_629) );
INVx1_ASAP7_75t_L g700 ( .A(n_583), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_584), .A2(n_667), .B(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_591), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_597), .Y(n_593) );
INVx1_ASAP7_75t_L g633 ( .A(n_594), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_595), .A2(n_681), .B1(n_684), .B2(n_686), .C(n_689), .Y(n_680) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_603), .A2(n_693), .B1(n_694), .B2(n_696), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g669 ( .A(n_605), .Y(n_669) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp67_ASAP7_75t_SL g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g673 ( .A(n_609), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g638 ( .A(n_614), .Y(n_638) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_619), .B(n_643), .Y(n_695) );
INVxp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_625), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_626), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g718 ( .A(n_626), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_633), .B(n_634), .C(n_668), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B(n_641), .C(n_660), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g721 ( .A(n_645), .Y(n_721) );
AND2x2_ASAP7_75t_L g658 ( .A(n_647), .B(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B1(n_656), .B2(n_658), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OR2x2_ASAP7_75t_L g666 ( .A(n_654), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g719 ( .A(n_655), .Y(n_719) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI31xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .A3(n_663), .B(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_672), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_677), .Y(n_676) );
NAND5xp2_ASAP7_75t_L g679 ( .A(n_680), .B(n_692), .C(n_699), .D(n_713), .E(n_716), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_691), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_716) );
INVx1_ASAP7_75t_SL g715 ( .A(n_693), .Y(n_715) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B(n_710), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
endmodule