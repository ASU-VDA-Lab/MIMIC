module fake_jpeg_28501_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx11_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx12_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_13),
.B1(n_10),
.B2(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_14),
.B1(n_34),
.B2(n_41),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_19),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_14),
.B(n_19),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI32xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_26),
.A3(n_32),
.B1(n_25),
.B2(n_21),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_37),
.B(n_43),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_49),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_61),
.C(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_51),
.B(n_50),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_40),
.B(n_53),
.C(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_54),
.C(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVxp33_ASAP7_75t_SL g68 ( 
.A(n_67),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_65),
.Y(n_69)
);


endmodule