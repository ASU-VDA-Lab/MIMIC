module fake_jpeg_19739_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_29),
.B1(n_19),
.B2(n_20),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_30),
.B(n_22),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_21),
.B(n_26),
.Y(n_87)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_47),
.B1(n_58),
.B2(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_70),
.Y(n_94)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_71),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_25),
.B1(n_35),
.B2(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_75),
.Y(n_99)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_31),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_34),
.B(n_36),
.C(n_38),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_34),
.B(n_51),
.C(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_84),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_40),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_53),
.B1(n_43),
.B2(n_33),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_0),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_34),
.B1(n_21),
.B2(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_45),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_101),
.Y(n_137)
);

HB1xp67_ASAP7_75t_SL g123 ( 
.A(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_98),
.B1(n_100),
.B2(n_107),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_34),
.B1(n_43),
.B2(n_33),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_86),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_102),
.B1(n_74),
.B2(n_81),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_82),
.B1(n_83),
.B2(n_72),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_34),
.B1(n_33),
.B2(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_16),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_9),
.B1(n_15),
.B2(n_2),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_85),
.C(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_28),
.B1(n_17),
.B2(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_0),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_61),
.B(n_65),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_117),
.B(n_124),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_80),
.B1(n_75),
.B2(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_61),
.B1(n_69),
.B2(n_64),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_131),
.B1(n_97),
.B2(n_96),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_60),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_129),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_86),
.C(n_81),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_141),
.C(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_136),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_7),
.B1(n_15),
.B2(n_2),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_140),
.B(n_5),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_28),
.B1(n_17),
.B2(n_0),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_113),
.B1(n_112),
.B2(n_105),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_88),
.A2(n_28),
.B1(n_17),
.B2(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_93),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_28),
.C(n_17),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_6),
.C(n_2),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_108),
.B(n_101),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_148),
.B1(n_156),
.B2(n_161),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_153),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_95),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_155),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_139),
.B(n_95),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_106),
.C(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_97),
.B1(n_92),
.B2(n_100),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_105),
.C(n_114),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_131),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_1),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_3),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_4),
.B(n_5),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_170),
.Y(n_180)
);

AOI22x1_ASAP7_75t_SL g168 ( 
.A1(n_115),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_139),
.B1(n_127),
.B2(n_122),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_129),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_147),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_195),
.C(n_183),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_191),
.CI(n_194),
.CON(n_201),
.SN(n_201)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_138),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_135),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_130),
.C(n_12),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_11),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_187),
.B(n_194),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_195),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_190),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_153),
.CI(n_144),
.CON(n_208),
.SN(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_159),
.C(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_182),
.C(n_152),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_156),
.B1(n_148),
.B2(n_167),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_186),
.B1(n_177),
.B2(n_150),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_145),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_193),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_151),
.C(n_192),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_198),
.C(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_143),
.B1(n_215),
.B2(n_150),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_168),
.B(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_227),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_186),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_197),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_244),
.C(n_217),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_238),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_230),
.B(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_207),
.B1(n_213),
.B2(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_202),
.C(n_201),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_201),
.C(n_200),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_250),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_199),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_249),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_214),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_253),
.Y(n_259)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_227),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_222),
.B1(n_212),
.B2(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_249),
.A2(n_155),
.B1(n_196),
.B2(n_223),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_231),
.B(n_200),
.Y(n_263)
);

OAI211xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_206),
.B(n_165),
.C(n_216),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_248),
.CI(n_247),
.CON(n_265),
.SN(n_265)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_269),
.C(n_158),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_267),
.A3(n_268),
.B1(n_169),
.B2(n_171),
.C1(n_149),
.C2(n_161),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_252),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_235),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_261),
.B(n_260),
.C(n_187),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_271),
.A3(n_272),
.B1(n_264),
.B2(n_158),
.C1(n_13),
.C2(n_12),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_164),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_11),
.B(n_13),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_275),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_13),
.Y(n_278)
);


endmodule