module real_aes_11486_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g582 ( .A(n_0), .B(n_58), .Y(n_582) );
AND2x2_ASAP7_75t_L g599 ( .A(n_0), .B(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_0), .Y(n_635) );
INVx1_ASAP7_75t_L g673 ( .A(n_0), .Y(n_673) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_1), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_2), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_3), .B(n_121), .Y(n_205) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_4), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_5), .Y(n_685) );
INVx1_ASAP7_75t_L g573 ( .A(n_6), .Y(n_573) );
OR2x2_ASAP7_75t_L g499 ( .A(n_7), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g532 ( .A(n_7), .Y(n_532) );
BUFx2_ASAP7_75t_L g493 ( .A(n_8), .Y(n_493) );
OR2x2_ASAP7_75t_L g581 ( .A(n_8), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g585 ( .A(n_8), .Y(n_585) );
INVx1_ASAP7_75t_L g598 ( .A(n_8), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_9), .A2(n_12), .B1(n_520), .B2(n_525), .C(n_529), .Y(n_519) );
INVx1_ASAP7_75t_L g607 ( .A(n_9), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_10), .B(n_118), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_11), .B(n_104), .Y(n_196) );
INVx1_ASAP7_75t_L g601 ( .A(n_12), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_13), .B(n_104), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_14), .B(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_14), .Y(n_719) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_15), .Y(n_683) );
AND2x2_ASAP7_75t_L g172 ( .A(n_16), .B(n_173), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_17), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_17), .Y(n_485) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_19), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_20), .B(n_182), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g133 ( .A(n_21), .B(n_134), .Y(n_133) );
NAND2xp33_ASAP7_75t_L g194 ( .A(n_22), .B(n_134), .Y(n_194) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_23), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_24), .Y(n_233) );
INVx1_ASAP7_75t_L g500 ( .A(n_25), .Y(n_500) );
INVx1_ASAP7_75t_L g533 ( .A(n_25), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_26), .B(n_120), .Y(n_139) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_27), .Y(n_693) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_28), .A2(n_51), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_29), .A2(n_136), .B(n_177), .C(n_179), .Y(n_176) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_30), .A2(n_45), .B1(n_554), .B2(n_556), .C(n_559), .Y(n_553) );
INVx1_ASAP7_75t_L g647 ( .A(n_30), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_31), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g112 ( .A(n_32), .B(n_113), .Y(n_112) );
NAND2xp33_ASAP7_75t_L g154 ( .A(n_33), .B(n_148), .Y(n_154) );
AND2x6_ASAP7_75t_L g83 ( .A(n_34), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_34), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_34), .B(n_676), .Y(n_723) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_35), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_36), .A2(n_68), .B1(n_541), .B2(n_548), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_36), .A2(n_68), .B1(n_620), .B2(n_626), .C(n_630), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_37), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_38), .B(n_178), .Y(n_193) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_39), .B(n_148), .Y(n_206) );
INVx1_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_40), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_41), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_42), .B(n_148), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_43), .A2(n_64), .B1(n_563), .B2(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g655 ( .A(n_43), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_44), .A2(n_54), .B1(n_535), .B2(n_538), .Y(n_534) );
INVx1_ASAP7_75t_L g590 ( .A(n_44), .Y(n_590) );
INVx1_ASAP7_75t_L g649 ( .A(n_45), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_47), .Y(n_496) );
AND2x2_ASAP7_75t_L g181 ( .A(n_48), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_49), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g580 ( .A(n_50), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_52), .Y(n_138) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_53), .B(n_92), .Y(n_214) );
INVx1_ASAP7_75t_L g612 ( .A(n_54), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_55), .B(n_132), .Y(n_153) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_55), .Y(n_713) );
BUFx10_ASAP7_75t_L g709 ( .A(n_56), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_57), .B(n_91), .Y(n_190) );
INVx2_ASAP7_75t_L g600 ( .A(n_58), .Y(n_600) );
NAND2xp33_ASAP7_75t_L g220 ( .A(n_59), .B(n_118), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_60), .B(n_134), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_61), .Y(n_180) );
INVx2_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_63), .Y(n_239) );
INVx1_ASAP7_75t_L g641 ( .A(n_64), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_65), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_66), .B(n_125), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_67), .Y(n_201) );
INVx1_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_70), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_71), .Y(n_506) );
AND2x2_ASAP7_75t_L g242 ( .A(n_72), .B(n_104), .Y(n_242) );
INVx2_ASAP7_75t_L g579 ( .A(n_73), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_74), .B(n_182), .Y(n_221) );
INVx1_ASAP7_75t_L g503 ( .A(n_75), .Y(n_503) );
BUFx3_ASAP7_75t_L g510 ( .A(n_75), .Y(n_510) );
INVx1_ASAP7_75t_L g505 ( .A(n_76), .Y(n_505) );
BUFx3_ASAP7_75t_L g517 ( .A(n_76), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_483), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx8_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
NOR2xp67_ASAP7_75t_L g163 ( .A(n_82), .B(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_82), .A2(n_231), .B(n_237), .Y(n_230) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g721 ( .A1(n_86), .A2(n_722), .B(n_723), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_87), .A2(n_168), .B(n_172), .Y(n_167) );
BUFx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx3_ASAP7_75t_L g122 ( .A(n_88), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_88), .A2(n_153), .B(n_154), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_88), .Y(n_191) );
BUFx12f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
O2A1O1Ixp33_ASAP7_75t_L g109 ( .A1(n_89), .A2(n_110), .B(n_111), .C(n_112), .Y(n_109) );
INVx5_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx5_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx2_ASAP7_75t_L g216 ( .A(n_92), .Y(n_216) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
INVx2_ASAP7_75t_L g121 ( .A(n_93), .Y(n_121) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_93), .Y(n_170) );
INVx1_ASAP7_75t_L g175 ( .A(n_93), .Y(n_175) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NOR3x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_336), .C(n_419), .Y(n_95) );
NAND4xp75_ASAP7_75t_L g96 ( .A(n_97), .B(n_271), .C(n_302), .D(n_317), .Y(n_96) );
NOR2x1_ASAP7_75t_L g97 ( .A(n_98), .B(n_208), .Y(n_97) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_157), .Y(n_98) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_99), .A2(n_293), .B(n_300), .Y(n_292) );
INVx2_ASAP7_75t_L g339 ( .A(n_99), .Y(n_339) );
AND2x2_ASAP7_75t_L g399 ( .A(n_99), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_127), .Y(n_99) );
AND2x4_ASAP7_75t_L g315 ( .A(n_100), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g394 ( .A(n_100), .B(n_262), .Y(n_394) );
INVx2_ASAP7_75t_L g424 ( .A(n_100), .Y(n_424) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g295 ( .A(n_102), .Y(n_295) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_102), .Y(n_346) );
OAI21x1_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_108), .B(n_124), .Y(n_102) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_103), .A2(n_129), .B(n_140), .Y(n_128) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_103), .A2(n_199), .B(n_207), .Y(n_198) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_103), .A2(n_129), .B(n_140), .Y(n_248) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_103), .A2(n_108), .B(n_124), .Y(n_264) );
BUFx4f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g144 ( .A(n_104), .Y(n_144) );
INVx4_ASAP7_75t_L g165 ( .A(n_104), .Y(n_165) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_104), .A2(n_212), .B(n_221), .Y(n_211) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_104), .A2(n_212), .B(n_221), .Y(n_251) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_104), .A2(n_212), .B(n_221), .Y(n_299) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g126 ( .A(n_105), .Y(n_126) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g183 ( .A(n_106), .Y(n_183) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_123), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_110), .A2(n_688), .B1(n_689), .B2(n_694), .Y(n_687) );
INVx1_ASAP7_75t_L g694 ( .A(n_110), .Y(n_694) );
INVx5_ASAP7_75t_L g219 ( .A(n_113), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B(n_119), .C(n_122), .Y(n_114) );
O2A1O1Ixp5_ASAP7_75t_L g137 ( .A1(n_116), .A2(n_122), .B(n_138), .C(n_139), .Y(n_137) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g132 ( .A(n_118), .Y(n_132) );
INVx2_ASAP7_75t_SL g178 ( .A(n_118), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_118), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
INVx2_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_L g200 ( .A1(n_122), .A2(n_201), .B(n_202), .C(n_203), .Y(n_200) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_123), .A2(n_130), .B(n_137), .Y(n_129) );
OAI21x1_ASAP7_75t_L g187 ( .A1(n_123), .A2(n_188), .B(n_192), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_123), .A2(n_200), .B(n_204), .Y(n_199) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_123), .A2(n_213), .B(n_217), .Y(n_212) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g321 ( .A(n_127), .Y(n_321) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_127), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_141), .Y(n_127) );
INVx2_ASAP7_75t_L g225 ( .A(n_128), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_135), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_134), .B(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_135), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_135), .A2(n_214), .B(n_215), .Y(n_213) );
CKINVDCx6p67_ASAP7_75t_R g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_SL g236 ( .A(n_136), .Y(n_236) );
INVx2_ASAP7_75t_L g226 ( .A(n_141), .Y(n_226) );
OR2x2_ASAP7_75t_L g287 ( .A(n_141), .B(n_264), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_141), .B(n_225), .Y(n_316) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_156), .Y(n_142) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_143), .A2(n_187), .B(n_196), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_143), .A2(n_145), .B(n_156), .Y(n_253) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_155), .Y(n_145) );
AOI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_151), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_148), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx1_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_151), .A2(n_218), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_184), .Y(n_158) );
OR2x2_ASAP7_75t_L g387 ( .A(n_159), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g418 ( .A(n_159), .Y(n_418) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g227 ( .A(n_160), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g451 ( .A(n_160), .B(n_304), .Y(n_451) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_161), .B(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g397 ( .A(n_161), .Y(n_397) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_161), .Y(n_466) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g258 ( .A(n_162), .Y(n_258) );
AOI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_181), .Y(n_162) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_165), .A2(n_230), .B(n_242), .Y(n_229) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_165), .A2(n_230), .B(n_242), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_176), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g240 ( .A(n_169), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_SL g259 ( .A(n_184), .Y(n_259) );
INVx1_ASAP7_75t_L g382 ( .A(n_184), .Y(n_382) );
OR2x2_ASAP7_75t_L g470 ( .A(n_184), .B(n_286), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_184), .B(n_354), .Y(n_479) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_197), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g228 ( .A(n_186), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g275 ( .A(n_186), .B(n_197), .Y(n_275) );
INVx1_ASAP7_75t_L g290 ( .A(n_186), .Y(n_290) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_186), .Y(n_326) );
AND2x2_ASAP7_75t_L g362 ( .A(n_186), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g390 ( .A(n_186), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp33_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_238), .B(n_240), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
BUFx3_ASAP7_75t_L g343 ( .A(n_197), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_197), .B(n_257), .Y(n_448) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g269 ( .A(n_198), .Y(n_269) );
OAI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_227), .B(n_243), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
INVx2_ASAP7_75t_L g282 ( .A(n_211), .Y(n_282) );
INVx2_ASAP7_75t_L g314 ( .A(n_211), .Y(n_314) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_211), .Y(n_400) );
AND2x2_ASAP7_75t_L g452 ( .A(n_211), .B(n_252), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g234 ( .A(n_219), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_222), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g345 ( .A(n_223), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
AND2x2_ASAP7_75t_L g263 ( .A(n_224), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g332 ( .A(n_224), .B(n_299), .Y(n_332) );
AND2x2_ASAP7_75t_L g378 ( .A(n_224), .B(n_299), .Y(n_378) );
INVx1_ASAP7_75t_L g385 ( .A(n_224), .Y(n_385) );
OR2x2_ASAP7_75t_L g450 ( .A(n_224), .B(n_250), .Y(n_450) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g262 ( .A(n_226), .Y(n_262) );
AND2x2_ASAP7_75t_L g283 ( .A(n_226), .B(n_248), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_227), .A2(n_334), .B1(n_339), .B2(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g270 ( .A(n_228), .Y(n_270) );
OR2x2_ASAP7_75t_L g334 ( .A(n_228), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g276 ( .A(n_229), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g301 ( .A(n_229), .B(n_258), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_234), .B(n_236), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_254), .B1(n_260), .B2(n_265), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_245), .A2(n_288), .B1(n_358), .B2(n_359), .Y(n_357) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
AND2x2_ASAP7_75t_L g435 ( .A(n_246), .B(n_279), .Y(n_435) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_247), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_247), .B(n_295), .Y(n_445) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
INVx1_ASAP7_75t_L g286 ( .A(n_250), .Y(n_286) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g309 ( .A(n_251), .Y(n_309) );
BUFx2_ASAP7_75t_L g376 ( .A(n_251), .Y(n_376) );
INVx1_ASAP7_75t_L g444 ( .A(n_251), .Y(n_444) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g280 ( .A(n_253), .B(n_264), .Y(n_280) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_259), .Y(n_254) );
AND2x2_ASAP7_75t_L g356 ( .A(n_255), .B(n_343), .Y(n_356) );
AND2x4_ASAP7_75t_L g427 ( .A(n_255), .B(n_275), .Y(n_427) );
INVx1_ASAP7_75t_L g442 ( .A(n_255), .Y(n_442) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_256), .Y(n_461) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_257), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g354 ( .A(n_257), .Y(n_354) );
INVx1_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
INVx1_ASAP7_75t_L g363 ( .A(n_258), .Y(n_363) );
INVx1_ASAP7_75t_L g358 ( .A(n_260), .Y(n_358) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_262), .B(n_295), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_264), .Y(n_371) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g379 ( .A(n_267), .B(n_335), .Y(n_379) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVxp67_ASAP7_75t_L g417 ( .A(n_268), .Y(n_417) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g325 ( .A(n_269), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_269), .B(n_270), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_269), .B(n_354), .Y(n_360) );
AND2x2_ASAP7_75t_L g389 ( .A(n_269), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_269), .B(n_397), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_278), .B(n_284), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g431 ( .A(n_274), .Y(n_431) );
NAND2xp67_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g348 ( .A(n_275), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_275), .B(n_301), .Y(n_411) );
AND2x4_ASAP7_75t_L g323 ( .A(n_276), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g350 ( .A(n_276), .Y(n_350) );
INVx1_ASAP7_75t_L g335 ( .A(n_277), .Y(n_335) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g330 ( .A(n_279), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g340 ( .A(n_279), .Y(n_340) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B(n_292), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_285), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_413) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g410 ( .A(n_286), .Y(n_410) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
OR2x2_ASAP7_75t_L g395 ( .A(n_289), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x2_ASAP7_75t_L g426 ( .A(n_294), .B(n_378), .Y(n_426) );
INVx1_ASAP7_75t_L g468 ( .A(n_294), .Y(n_468) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
AND2x2_ASAP7_75t_L g423 ( .A(n_296), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_297), .Y(n_458) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_299), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g381 ( .A(n_301), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_301), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_301), .B(n_434), .Y(n_433) );
NAND2x1_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_312), .Y(n_305) );
INVxp33_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
AND2x2_ASAP7_75t_L g476 ( .A(n_308), .B(n_394), .Y(n_476) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2x1_ASAP7_75t_SL g449 ( .A(n_311), .B(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g437 ( .A(n_312), .Y(n_437) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_343), .Y(n_342) );
AO22x1_ASAP7_75t_L g327 ( .A1(n_315), .A2(n_328), .B1(n_330), .B2(n_333), .Y(n_327) );
AND2x2_ASAP7_75t_L g374 ( .A(n_316), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g467 ( .A(n_316), .B(n_468), .Y(n_467) );
O2A1O1Ixp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B(n_323), .C(n_327), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_319), .A2(n_399), .B1(n_401), .B2(n_403), .C(n_408), .Y(n_398) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g415 ( .A(n_320), .B(n_392), .Y(n_415) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_322), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g482 ( .A(n_332), .Y(n_482) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g474 ( .A(n_335), .Y(n_474) );
NAND4xp75_ASAP7_75t_L g336 ( .A(n_337), .B(n_364), .C(n_398), .D(n_412), .Y(n_336) );
AOI221x1_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B1(n_344), .B2(n_347), .C(n_357), .Y(n_337) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g434 ( .A(n_343), .Y(n_434) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
OAI211xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_349), .B(n_351), .C(n_355), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_348), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g416 ( .A(n_352), .Y(n_416) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_380), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_372), .B(n_379), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_367), .A2(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_368), .B(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
BUFx2_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
NAND2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_386), .Y(n_380) );
AND2x2_ASAP7_75t_L g464 ( .A(n_382), .B(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_383), .A2(n_431), .B(n_455), .C(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_389), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g407 ( .A(n_390), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_392), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_394), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_418), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND4xp75_ASAP7_75t_L g419 ( .A(n_420), .B(n_436), .C(n_453), .D(n_462), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_427), .B(n_428), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g455 ( .A(n_424), .Y(n_455) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AO22x1_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_432), .B2(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_443), .B(n_446), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_441), .A2(n_476), .B1(n_477), .B2(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_449), .B1(n_451), .B2(n_452), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_455), .A2(n_457), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g472 ( .A(n_460), .Y(n_472) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_475), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B1(n_469), .B2(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B1(n_674), .B2(n_679), .C(n_716), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_486), .A2(n_717), .B1(n_719), .B2(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_587), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_494), .B1(n_573), .B2(n_574), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x6_ASAP7_75t_L g633 ( .A(n_493), .B(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g494 ( .A(n_495), .B(n_512), .C(n_552), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_506), .B2(n_507), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_496), .A2(n_570), .B1(n_638), .B2(n_663), .Y(n_662) );
INVx6_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx2_ASAP7_75t_L g511 ( .A(n_499), .Y(n_511) );
OR2x2_ASAP7_75t_L g514 ( .A(n_499), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g544 ( .A(n_500), .Y(n_544) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g516 ( .A(n_503), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g509 ( .A(n_505), .B(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_506), .A2(n_518), .B1(n_650), .B2(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_509), .Y(n_537) );
INVx2_ASAP7_75t_SL g555 ( .A(n_509), .Y(n_555) );
INVx2_ASAP7_75t_L g523 ( .A(n_510), .Y(n_523) );
AND2x2_ASAP7_75t_L g528 ( .A(n_510), .B(n_517), .Y(n_528) );
AND2x4_ASAP7_75t_L g569 ( .A(n_511), .B(n_527), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_518), .B1(n_519), .B2(n_534), .C(n_540), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_516), .Y(n_539) );
INVx2_ASAP7_75t_L g524 ( .A(n_517), .Y(n_524) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx6_ASAP7_75t_L g565 ( .A(n_522), .Y(n_565) );
AND2x2_ASAP7_75t_L g586 ( .A(n_522), .B(n_543), .Y(n_586) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g551 ( .A(n_523), .Y(n_551) );
INVx1_ASAP7_75t_L g547 ( .A(n_524), .Y(n_547) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g571 ( .A(n_527), .B(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_528), .Y(n_558) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x4_ASAP7_75t_L g543 ( .A(n_531), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_533), .Y(n_561) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x4_ASAP7_75t_L g549 ( .A(n_543), .B(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g572 ( .A(n_543), .Y(n_572) );
AND2x4_ASAP7_75t_L g712 ( .A(n_543), .B(n_545), .Y(n_712) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g707 ( .A(n_546), .Y(n_707) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_562), .B1(n_567), .B2(n_570), .C(n_571), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g704 ( .A(n_561), .Y(n_704) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_583), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .Y(n_576) );
BUFx2_ASAP7_75t_L g640 ( .A(n_577), .Y(n_640) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g595 ( .A(n_579), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g605 ( .A(n_579), .Y(n_605) );
AND2x2_ASAP7_75t_L g611 ( .A(n_579), .B(n_580), .Y(n_611) );
INVx2_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
INVx1_ASAP7_75t_L g646 ( .A(n_579), .Y(n_646) );
INVx2_ASAP7_75t_L g596 ( .A(n_580), .Y(n_596) );
INVx1_ASAP7_75t_L g618 ( .A(n_580), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
INVx1_ASAP7_75t_L g645 ( .A(n_580), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_580), .B(n_616), .Y(n_654) );
INVx3_ASAP7_75t_L g625 ( .A(n_581), .Y(n_625) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_619), .C(n_632), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_606), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_601), .B2(n_602), .Y(n_589) );
BUFx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g659 ( .A(n_594), .Y(n_659) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g604 ( .A(n_596), .B(n_605), .Y(n_604) );
AND2x6_ASAP7_75t_L g602 ( .A(n_597), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g608 ( .A(n_597), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g613 ( .A(n_597), .B(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g670 ( .A(n_598), .Y(n_670) );
INVx1_ASAP7_75t_L g636 ( .A(n_600), .Y(n_636) );
INVx1_ASAP7_75t_L g672 ( .A(n_600), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_603), .B(n_625), .Y(n_631) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_612), .B2(n_613), .Y(n_606) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g629 ( .A(n_616), .Y(n_629) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2x1_ASAP7_75t_SL g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_625), .B(n_628), .Y(n_627) );
BUFx4f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .A3(n_648), .B1(n_660), .B2(n_662), .B3(n_667), .Y(n_632) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B1(n_642), .B2(n_647), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_645), .B(n_646), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_655), .B2(n_656), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
CKINVDCx8_ASAP7_75t_R g667 ( .A(n_668), .Y(n_667) );
INVx5_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x6_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_676), .B(n_678), .Y(n_700) );
INVx1_ASAP7_75t_SL g722 ( .A(n_676), .Y(n_722) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_696), .B1(n_713), .B2(n_714), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_680), .A2(n_713), .B1(n_715), .B2(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_687), .B2(n_695), .Y(n_680) );
CKINVDCx14_ASAP7_75t_R g695 ( .A(n_681), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx8_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx8_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_699), .Y(n_718) );
OR2x6_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OR2x4_ASAP7_75t_L g715 ( .A(n_700), .B(n_702), .Y(n_715) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI31xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .A3(n_708), .B(n_710), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx6_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
endmodule