module fake_jpeg_3582_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_1),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_60),
.B1(n_61),
.B2(n_57),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_83),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_60),
.C(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_67),
.B1(n_48),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_67),
.B1(n_52),
.B2(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_51),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_53),
.B1(n_65),
.B2(n_62),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_63),
.B(n_49),
.C(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_11),
.Y(n_120)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_59),
.B1(n_54),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_11),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_89),
.B1(n_84),
.B2(n_43),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_14),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_6),
.B(n_7),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_12),
.B(n_13),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_119),
.B1(n_104),
.B2(n_107),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_28),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_116),
.B1(n_96),
.B2(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_35),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_27),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_33),
.C(n_32),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_25),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_132),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_95),
.B1(n_31),
.B2(n_30),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_143),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_29),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_148),
.C(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_140),
.C(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_14),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_21),
.B1(n_22),
.B2(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_123),
.C(n_113),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_112),
.B(n_16),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_15),
.C(n_17),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_19),
.C(n_20),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_163),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_19),
.B(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

AO22x1_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_133),
.B1(n_145),
.B2(n_135),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_166),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_21),
.B1(n_22),
.B2(n_154),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_156),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_150),
.C(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_151),
.C(n_168),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_161),
.A3(n_177),
.B1(n_154),
.B2(n_171),
.C1(n_176),
.C2(n_174),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_189),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_157),
.A3(n_159),
.B1(n_160),
.B2(n_162),
.C1(n_177),
.C2(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_180),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_188),
.C(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_193),
.B(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);


endmodule