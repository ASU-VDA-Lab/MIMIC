module real_jpeg_10339_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_266, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_266;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_1),
.A2(n_20),
.B1(n_40),
.B2(n_41),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_20),
.B1(n_55),
.B2(n_56),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_10),
.B(n_25),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_54)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_40),
.B(n_54),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_40),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_10),
.B(n_56),
.Y(n_148)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_11),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_10),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_10),
.A2(n_29),
.B1(n_55),
.B2(n_56),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_74),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_10),
.A2(n_24),
.B(n_39),
.C(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_22),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_23),
.B(n_26),
.C(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_26),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_11),
.A2(n_26),
.B(n_29),
.C(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_106),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_105),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_16),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_66),
.C(n_75),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_17),
.B(n_66),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_32),
.B1(n_33),
.B2(n_65),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_18),
.A2(n_65),
.B1(n_94),
.B2(n_103),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_18),
.A2(n_65),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_18),
.B(n_119),
.C(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_18),
.A2(n_65),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_18),
.B(n_230),
.C(n_232),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_19),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_23),
.B(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_96),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_24),
.A2(n_38),
.B(n_39),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_29),
.A2(n_41),
.B(n_59),
.C(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_29),
.B(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_29),
.B(n_54),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_29),
.A2(n_40),
.B(n_44),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B(n_45),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_36),
.A2(n_72),
.B1(n_74),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_46),
.A2(n_71),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_47),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_51),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_64),
.C(n_65),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_53),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_68),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_54),
.A2(n_60),
.B1(n_88),
.B2(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_55),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_69),
.A2(n_70),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_69),
.A2(n_70),
.B1(n_95),
.B2(n_102),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_70),
.B(n_137),
.C(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_70),
.B(n_102),
.C(n_222),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_72),
.B(n_74),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_75),
.A2(n_76),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_89),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_89),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_77),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_77),
.A2(n_85),
.B1(n_124),
.B2(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_79),
.B(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_83),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_81),
.A2(n_82),
.B1(n_139),
.B2(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_82),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_138),
.B(n_140),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_84),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_95),
.A2(n_102),
.B1(n_119),
.B2(n_174),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_111),
.C(n_119),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_129),
.B(n_264),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_126),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_108),
.B(n_126),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_120),
.C(n_121),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_109),
.A2(n_110),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_111),
.A2(n_112),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_114),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_117),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_116),
.A2(n_117),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_157),
.C(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_184),
.C(n_191),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_143),
.B1(n_149),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_119),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_143),
.C(n_179),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_119),
.A2(n_174),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_120),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

AOI321xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_239),
.A3(n_252),
.B1(n_258),
.B2(n_263),
.C(n_266),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_211),
.C(n_236),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_193),
.B(n_210),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_181),
.B(n_192),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_169),
.B(n_180),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_160),
.B(n_168),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_150),
.B(n_159),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_142),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_152),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_143),
.A2(n_149),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_149),
.B(n_216),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B(n_158),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_167),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_179),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_183),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_195),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_203),
.C(n_209),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_213),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_213),
.B(n_223),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_219),
.CI(n_220),
.CON(n_213),
.SN(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_235),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.C(n_235),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_259),
.B(n_262),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_249),
.C(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule