module fake_netlist_1_3978_n_443 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_443, n_188);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_443;
output n_188;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g65 ( .A(n_5), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_21), .Y(n_66) );
INVxp67_ASAP7_75t_SL g67 ( .A(n_36), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_8), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_37), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_48), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_26), .Y(n_71) );
CKINVDCx20_ASAP7_75t_R g72 ( .A(n_25), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_0), .Y(n_73) );
INVxp33_ASAP7_75t_SL g74 ( .A(n_10), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_59), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_14), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_40), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_29), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_24), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_42), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g81 ( .A(n_64), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_39), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_56), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_31), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_63), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_34), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_54), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_61), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_10), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_46), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_60), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_66), .Y(n_97) );
INVx3_ASAP7_75t_L g98 ( .A(n_88), .Y(n_98) );
INVx3_ASAP7_75t_L g99 ( .A(n_88), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_91), .Y(n_100) );
AND2x6_ASAP7_75t_L g101 ( .A(n_66), .B(n_27), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_68), .B(n_0), .Y(n_103) );
NAND2xp33_ASAP7_75t_SL g104 ( .A(n_72), .B(n_1), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_91), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_96), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_76), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_76), .Y(n_113) );
INVx5_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_87), .B(n_1), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_94), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_79), .B(n_2), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_109), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_108), .B(n_94), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_97), .B(n_68), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_100), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_97), .B(n_73), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_102), .B(n_83), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_102), .B(n_73), .Y(n_128) );
AND2x6_ASAP7_75t_L g129 ( .A(n_107), .B(n_95), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_109), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_109), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_100), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_113), .B(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_107), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_100), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_105), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_110), .B(n_85), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_101), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_105), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_122), .B(n_116), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g148 ( .A(n_144), .B(n_110), .C(n_112), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_123), .B(n_111), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_123), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_128), .B(n_111), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_136), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
AND2x6_ASAP7_75t_SL g159 ( .A(n_125), .B(n_115), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_129), .A2(n_101), .B1(n_112), .B2(n_107), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_126), .B(n_114), .Y(n_161) );
CKINVDCx6p67_ASAP7_75t_R g162 ( .A(n_129), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_142), .B(n_114), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_129), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_121), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_130), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_130), .B(n_114), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_131), .Y(n_173) );
INVx1_ASAP7_75t_SL g174 ( .A(n_131), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_133), .B(n_114), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_135), .B(n_114), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_135), .Y(n_178) );
INVx2_ASAP7_75t_R g179 ( .A(n_166), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_158), .B(n_103), .Y(n_180) );
NAND2x1_ASAP7_75t_L g181 ( .A(n_149), .B(n_101), .Y(n_181) );
BUFx12f_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_178), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_158), .B(n_103), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_178), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
UNKNOWN g188 ( );
INVx5_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_150), .A2(n_118), .B1(n_92), .B2(n_119), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_150), .A2(n_101), .B1(n_104), .B2(n_65), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_106), .B(n_119), .C(n_90), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_148), .A2(n_106), .B(n_77), .C(n_96), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_153), .B(n_93), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_149), .B(n_101), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_156), .A2(n_74), .B1(n_101), .B2(n_67), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_152), .B(n_99), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_154), .B(n_99), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_157), .B(n_99), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
BUFx12f_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_155), .B(n_99), .Y(n_206) );
BUFx4f_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_183), .B(n_98), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_183), .A2(n_168), .B1(n_165), .B2(n_167), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_180), .B(n_160), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_209), .A2(n_167), .B(n_163), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_189), .B(n_166), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_203), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_185), .B(n_169), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_203), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_197), .B(n_169), .Y(n_219) );
BUFx10_ASAP7_75t_L g220 ( .A(n_195), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_180), .B(n_146), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_189), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_188), .A2(n_161), .B1(n_117), .B2(n_77), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g224 ( .A1(n_182), .A2(n_98), .B1(n_95), .B2(n_90), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_204), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_193), .A2(n_140), .B(n_132), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_198), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_207), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_189), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_198), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_229), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_229), .Y(n_235) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_192), .B(n_204), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_215), .B(n_186), .Y(n_237) );
AOI221xp5_ASAP7_75t_L g238 ( .A1(n_224), .A2(n_184), .B1(n_190), .B2(n_194), .C(n_206), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_228), .A2(n_207), .B1(n_186), .B2(n_196), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_215), .B(n_206), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_233), .A2(n_205), .B1(n_182), .B2(n_191), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_218), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_218), .B(n_199), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_230), .A2(n_197), .B1(n_205), .B2(n_208), .Y(n_245) );
BUFx4f_ASAP7_75t_SL g246 ( .A(n_210), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_230), .A2(n_197), .B1(n_208), .B2(n_200), .Y(n_247) );
INVx6_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_225), .A2(n_202), .B(n_84), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_223), .A2(n_201), .B1(n_98), .B2(n_117), .C(n_105), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_232), .B(n_187), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_242), .Y(n_255) );
AOI22xp5_ASAP7_75t_SL g256 ( .A1(n_245), .A2(n_232), .B1(n_217), .B2(n_226), .Y(n_256) );
OAI222xp33_ASAP7_75t_L g257 ( .A1(n_246), .A2(n_231), .B1(n_222), .B2(n_211), .C1(n_219), .C2(n_212), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_232), .B1(n_219), .B2(n_222), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_253), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_244), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g263 ( .A1(n_248), .A2(n_232), .B1(n_216), .B2(n_217), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_241), .B(n_201), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_244), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_254), .B(n_220), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_250), .B(n_105), .C(n_117), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
OAI221xp5_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_98), .B1(n_78), .B2(n_117), .C(n_181), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_254), .B(n_227), .Y(n_274) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_240), .A2(n_82), .B(n_89), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_240), .B(n_227), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_236), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_271), .Y(n_278) );
OAI33xp33_ASAP7_75t_L g279 ( .A1(n_259), .A2(n_86), .A3(n_243), .B1(n_247), .B2(n_138), .B3(n_140), .Y(n_279) );
BUFx2_ASAP7_75t_SL g280 ( .A(n_272), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_264), .B(n_249), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_265), .B(n_145), .C(n_127), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_260), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_261), .B(n_249), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_276), .B(n_236), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_276), .B(n_236), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_267), .B(n_249), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_274), .B(n_217), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_274), .B(n_226), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_270), .Y(n_291) );
NAND4xp25_ASAP7_75t_L g292 ( .A(n_268), .B(n_251), .C(n_138), .D(n_132), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_272), .B(n_227), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_263), .A2(n_248), .B1(n_231), .B2(n_222), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_262), .B(n_227), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_255), .B(n_226), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_277), .B(n_2), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_3), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
AO31x2_ASAP7_75t_L g304 ( .A1(n_256), .A2(n_231), .A3(n_222), .B(n_124), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_273), .B(n_4), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_257), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_269), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_276), .B(n_4), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_291), .B(n_231), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_306), .A2(n_214), .B(n_187), .C(n_181), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_308), .B(n_5), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_289), .B(n_220), .Y(n_314) );
OAI31xp33_ASAP7_75t_L g315 ( .A1(n_305), .A2(n_195), .A3(n_214), .B(n_8), .Y(n_315) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_282), .B(n_127), .C(n_134), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_291), .B(n_219), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_289), .B(n_219), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_289), .Y(n_319) );
NOR2xp33_ASAP7_75t_R g320 ( .A(n_308), .B(n_248), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_280), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
NAND2xp33_ASAP7_75t_SL g323 ( .A(n_302), .B(n_214), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_298), .B(n_248), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_290), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_286), .B(n_6), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_288), .B(n_7), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_298), .B(n_7), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_293), .B(n_9), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_297), .B(n_11), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_300), .Y(n_333) );
AOI31xp33_ASAP7_75t_L g334 ( .A1(n_281), .A2(n_214), .A3(n_195), .B(n_12), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_286), .B(n_12), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_290), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_298), .B(n_208), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_290), .Y(n_338) );
NOR2xp33_ASAP7_75t_R g339 ( .A(n_301), .B(n_13), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_305), .B(n_124), .C(n_176), .D(n_175), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_299), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_284), .B(n_145), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_287), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_295), .B(n_208), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_285), .B(n_179), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_285), .B(n_15), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_279), .B(n_16), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_311), .B(n_303), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_334), .A2(n_307), .B1(n_294), .B2(n_296), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_321), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_334), .A2(n_296), .B(n_294), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_321), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_344), .B(n_17), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_340), .A2(n_219), .B1(n_127), .B2(n_134), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_336), .B(n_304), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_329), .B(n_127), .C(n_134), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_127), .B1(n_134), .B2(n_139), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_320), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_335), .B(n_18), .Y(n_363) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_315), .B(n_327), .C(n_313), .D(n_343), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_319), .B(n_304), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_339), .B(n_304), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_348), .A2(n_145), .B(n_141), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_326), .B(n_19), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_341), .B(n_145), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_338), .B(n_141), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_328), .B(n_141), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_314), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_331), .B(n_141), .Y(n_375) );
OAI21xp33_ASAP7_75t_L g376 ( .A1(n_322), .A2(n_134), .B(n_139), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_318), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_318), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_208), .B1(n_141), .B2(n_139), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_347), .B(n_20), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_315), .A2(n_177), .B(n_172), .Y(n_382) );
AOI322xp5_ASAP7_75t_L g383 ( .A1(n_323), .A2(n_139), .A3(n_23), .B1(n_32), .B2(n_33), .C1(n_35), .C2(n_38), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_309), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_317), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_325), .A2(n_22), .B1(n_41), .B2(n_43), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_354), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_370), .B(n_316), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_362), .A2(n_374), .B(n_352), .C(n_366), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_356), .B(n_346), .Y(n_390) );
NAND2xp33_ASAP7_75t_SL g391 ( .A(n_366), .B(n_337), .Y(n_391) );
BUFx8_ASAP7_75t_SL g392 ( .A(n_378), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_373), .B(n_310), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_357), .A2(n_44), .B(n_45), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_377), .B(n_47), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_358), .A2(n_49), .B(n_50), .C(n_51), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_368), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_376), .B(n_52), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_365), .B(n_53), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_360), .A2(n_170), .B(n_175), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_364), .B(n_57), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_357), .A2(n_151), .B1(n_171), .B2(n_62), .C(n_58), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_359), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_385), .Y(n_409) );
NAND4xp75_ASAP7_75t_L g410 ( .A(n_406), .B(n_355), .C(n_384), .D(n_381), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_391), .A2(n_385), .B1(n_363), .B2(n_361), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_406), .A2(n_408), .B1(n_393), .B2(n_389), .Y(n_412) );
XOR2x2_ASAP7_75t_L g413 ( .A(n_387), .B(n_363), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_404), .B(n_369), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_408), .A2(n_367), .B1(n_386), .B2(n_372), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_394), .A2(n_380), .B1(n_371), .B2(n_375), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g417 ( .A1(n_398), .A2(n_380), .B(n_383), .C(n_382), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_399), .B(n_171), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_390), .A2(n_173), .B1(n_174), .B2(n_409), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_392), .B(n_405), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_410), .B(n_400), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_417), .A2(n_388), .B(n_398), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_420), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_416), .A2(n_402), .B1(n_407), .B2(n_397), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_421), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_413), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_412), .A2(n_395), .B1(n_403), .B2(n_411), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_419), .A2(n_418), .B1(n_415), .B2(n_414), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_414), .A2(n_389), .B1(n_412), .B2(n_391), .C(n_417), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_417), .A2(n_389), .B1(n_396), .B2(n_408), .C(n_412), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_412), .A2(n_389), .B1(n_410), .B2(n_362), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_431), .B(n_427), .Y(n_433) );
INVx3_ASAP7_75t_SL g434 ( .A(n_424), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_426), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_432), .Y(n_436) );
OAI222xp33_ASAP7_75t_L g437 ( .A1(n_433), .A2(n_430), .B1(n_423), .B2(n_422), .C1(n_425), .C2(n_429), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_435), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_438), .B(n_436), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_437), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_439), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_441), .A2(n_440), .B1(n_439), .B2(n_434), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_442), .A2(n_423), .B(n_428), .Y(n_443) );
endmodule