module fake_netlist_1_2567_n_42 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_4), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
BUFx10_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_2), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_1), .Y(n_20) );
NAND2xp33_ASAP7_75t_L g21 ( .A(n_16), .B(n_11), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_19), .B(n_0), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_17), .B(n_3), .Y(n_24) );
NAND2xp5_ASAP7_75t_SL g25 ( .A(n_17), .B(n_5), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_17), .Y(n_26) );
OAI21xp33_ASAP7_75t_L g27 ( .A1(n_12), .A2(n_5), .B(n_6), .Y(n_27) );
OR2x6_ASAP7_75t_L g28 ( .A(n_24), .B(n_14), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_22), .Y(n_29) );
AO31x2_ASAP7_75t_L g30 ( .A1(n_23), .A2(n_17), .A3(n_13), .B(n_15), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_22), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_26), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_27), .B1(n_20), .B2(n_18), .C1(n_24), .C2(n_25), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
OAI211xp5_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_21), .B(n_28), .C(n_34), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_35), .B(n_36), .Y(n_38) );
BUFx12f_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_38), .Y(n_40) );
XOR2xp5_ASAP7_75t_L g41 ( .A(n_40), .B(n_6), .Y(n_41) );
OAI221xp5_ASAP7_75t_R g42 ( .A1(n_41), .A2(n_39), .B1(n_30), .B2(n_8), .C(n_7), .Y(n_42) );
endmodule