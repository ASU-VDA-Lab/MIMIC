module real_jpeg_11350_n_22 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_22);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_22;

wire n_43;
wire n_54;
wire n_37;
wire n_57;
wire n_65;
wire n_35;
wire n_33;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_31;
wire n_58;
wire n_52;
wire n_67;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_71;
wire n_42;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_70;
wire n_41;
wire n_27;
wire n_32;
wire n_56;
wire n_26;
wire n_48;
wire n_30;

AOI321xp33_ASAP7_75t_L g24 ( 
.A1(n_0),
.A2(n_25),
.A3(n_32),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

NOR4xp25_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_2),
.C(n_5),
.D(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_14),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_28),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_10),
.B1(n_11),
.B2(n_54),
.C(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_9),
.B(n_62),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_26),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

OAI221xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_18),
.B1(n_26),
.B2(n_29),
.C(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

OAI222xp33_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_12),
.B1(n_16),
.B2(n_37),
.C1(n_38),
.C2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_12),
.B(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_21),
.B1(n_38),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

OAI221xp5_ASAP7_75t_L g44 ( 
.A1(n_19),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_30),
.B(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_40),
.A3(n_43),
.B1(n_44),
.B2(n_51),
.Y(n_23)
);

OAI31xp33_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_31),
.A3(n_53),
.B(n_58),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_29),
.A2(n_55),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_53),
.B(n_58),
.Y(n_52)
);

AOI211xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_42),
.B(n_61),
.C(n_68),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_38),
.A3(n_42),
.B1(n_68),
.B2(n_70),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_41),
.B(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_59),
.A3(n_60),
.B1(n_62),
.B2(n_69),
.C1(n_71),
.C2(n_72),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR5xp2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.C(n_65),
.D(n_66),
.E(n_67),
.Y(n_62)
);


endmodule