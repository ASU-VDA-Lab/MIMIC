module fake_jpeg_26636_n_119 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_46),
.B1(n_18),
.B2(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_16),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_49),
.Y(n_60)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_13),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_62),
.B(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_46),
.B1(n_19),
.B2(n_15),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_24),
.B(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_37),
.B1(n_42),
.B2(n_49),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_75),
.B1(n_58),
.B2(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_48),
.B1(n_42),
.B2(n_21),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_70),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_74),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_43),
.C(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_60),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_79),
.C(n_81),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_60),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_59),
.C(n_58),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_56),
.B1(n_59),
.B2(n_62),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_71),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_93),
.B1(n_96),
.B2(n_77),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_69),
.B(n_58),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AOI21x1_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_74),
.B(n_64),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_95),
.B(n_21),
.C(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_63),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_40),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_15),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_103),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_1),
.C(n_2),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_25),
.A3(n_14),
.B1(n_45),
.B2(n_86),
.C(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_107),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_101),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_2),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_102),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_7),
.B(n_9),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.C(n_114),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_9),
.Y(n_119)
);


endmodule