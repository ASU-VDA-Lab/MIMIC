module fake_jpeg_27358_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_22),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx2_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_26),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_15),
.B1(n_13),
.B2(n_19),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_64),
.B1(n_65),
.B2(n_30),
.Y(n_79)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_38),
.B1(n_46),
.B2(n_33),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_32),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_36),
.C(n_34),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_48),
.C(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_28),
.B1(n_42),
.B2(n_46),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_80),
.B1(n_50),
.B2(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_83),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_47),
.C(n_50),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_30),
.B1(n_15),
.B2(n_23),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_77),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_60),
.B(n_47),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_94),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_62),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_47),
.B(n_14),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_80),
.B1(n_72),
.B2(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_100),
.B1(n_78),
.B2(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_102),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_51),
.B1(n_59),
.B2(n_54),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_47),
.B(n_32),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_82),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_31),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_31),
.C(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_124),
.B1(n_88),
.B2(n_104),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_118),
.B1(n_96),
.B2(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_81),
.B1(n_71),
.B2(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_66),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_93),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_101),
.B(n_82),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_73),
.B1(n_15),
.B2(n_27),
.Y(n_175)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_135),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_142),
.B1(n_147),
.B2(n_152),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_87),
.B1(n_94),
.B2(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_153),
.B1(n_15),
.B2(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_95),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_110),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_114),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_101),
.B1(n_87),
.B2(n_94),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_122),
.B(n_73),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_22),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_86),
.B1(n_67),
.B2(n_77),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_77),
.C(n_31),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_107),
.C(n_115),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_67),
.B1(n_59),
.B2(n_54),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_67),
.B1(n_73),
.B2(n_13),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_105),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_130),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_161),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_121),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_160),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_124),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_165),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_120),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_167),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_108),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_170),
.C(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_176),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_108),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_132),
.B(n_153),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_174),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_16),
.B1(n_18),
.B2(n_12),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_18),
.B(n_13),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_19),
.B1(n_14),
.B2(n_16),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_180),
.B1(n_18),
.B2(n_12),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_19),
.B1(n_14),
.B2(n_16),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_200),
.B(n_201),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_129),
.B1(n_132),
.B2(n_150),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_191),
.B1(n_201),
.B2(n_25),
.Y(n_210)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_151),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_198),
.B1(n_172),
.B2(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_12),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_29),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_0),
.B(n_1),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_12),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_164),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_182),
.B1(n_192),
.B2(n_200),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_155),
.C(n_156),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_181),
.C(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_196),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_175),
.B1(n_159),
.B2(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_220),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_0),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_217),
.Y(n_235)
);

FAx1_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_195),
.CI(n_190),
.CON(n_214),
.SN(n_214)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_25),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_29),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_182),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_207),
.C(n_187),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_229),
.C(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_199),
.C(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_213),
.C(n_214),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_191),
.C(n_184),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_188),
.C(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_236),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_27),
.C(n_20),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_249),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_243),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_214),
.C(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_247),
.C(n_20),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_21),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_21),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_27),
.C(n_20),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_1),
.B(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_258),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_3),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_R g271 ( 
.A(n_254),
.B(n_256),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_21),
.Y(n_267)
);

FAx1_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_4),
.CI(n_5),
.CON(n_256),
.SN(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_20),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_21),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_20),
.C(n_21),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_4),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_269),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_246),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_271),
.B1(n_268),
.B2(n_267),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_21),
.C(n_5),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_4),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_261),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_8),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_259),
.C(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_8),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_274),
.B(n_277),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_278),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

AOI321xp33_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_276),
.C(n_273),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_9),
.C(n_10),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_9),
.B(n_11),
.Y(n_288)
);


endmodule