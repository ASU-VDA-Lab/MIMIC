module fake_jpeg_16384_n_239 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_0),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_44),
.Y(n_64)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_54),
.Y(n_61)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_23),
.B1(n_14),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_20),
.B1(n_22),
.B2(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_18),
.Y(n_74)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_20),
.B2(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_35),
.B1(n_23),
.B2(n_14),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_69),
.B1(n_46),
.B2(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_67),
.B1(n_25),
.B2(n_24),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_20),
.B1(n_17),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_51),
.B1(n_41),
.B2(n_44),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_22),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_34),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_89),
.B1(n_92),
.B2(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_90),
.B1(n_76),
.B2(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_64),
.C(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_47),
.C(n_21),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_22),
.B(n_15),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_47),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_43),
.B1(n_33),
.B2(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_96),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_75),
.B1(n_71),
.B2(n_60),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_43),
.B1(n_41),
.B2(n_48),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_97),
.B1(n_93),
.B2(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_67),
.B1(n_69),
.B2(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_111),
.B1(n_85),
.B2(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_61),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_18),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_114),
.B(n_88),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_116),
.B1(n_90),
.B2(n_93),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_24),
.B(n_15),
.C(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_113),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_81),
.C(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_58),
.Y(n_134)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_132),
.B1(n_98),
.B2(n_115),
.Y(n_146)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_89),
.B(n_96),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_89),
.B(n_78),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_82),
.B(n_83),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_128),
.A2(n_129),
.B(n_111),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_47),
.B1(n_73),
.B2(n_36),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_73),
.B1(n_58),
.B2(n_52),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_73),
.B1(n_58),
.B2(n_52),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_108),
.B(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_146),
.B1(n_149),
.B2(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_157),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_151),
.C(n_120),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_124),
.A3(n_127),
.B1(n_129),
.B2(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_153),
.B(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_112),
.B1(n_99),
.B2(n_104),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_101),
.C(n_110),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_101),
.B(n_73),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_73),
.B1(n_52),
.B2(n_42),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_7),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_125),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_121),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_162),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_169),
.C(n_173),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_172),
.B(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_118),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_155),
.CI(n_146),
.CON(n_182),
.SN(n_182)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_131),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_123),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_123),
.C(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_151),
.C(n_141),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_183),
.C(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_8),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_147),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_156),
.C(n_145),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_7),
.B(n_12),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_26),
.C(n_1),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_168),
.C(n_159),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_170),
.B1(n_172),
.B2(n_10),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_26),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_26),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_26),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_8),
.B(n_12),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_6),
.B(n_11),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_2),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_198),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_177),
.B(n_186),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_182),
.B(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_184),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_179),
.C(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_194),
.B1(n_182),
.B2(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_212),
.B(n_222),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_196),
.B1(n_6),
.B2(n_5),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_221),
.C(n_208),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_5),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_3),
.B(n_4),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_6),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_10),
.C(n_11),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_11),
.C(n_4),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_231),
.C(n_225),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_3),
.C(n_4),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_233),
.A2(n_230),
.B(n_223),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_3),
.B(n_26),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_3),
.B(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_26),
.Y(n_239)
);


endmodule