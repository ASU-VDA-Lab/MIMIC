module fake_jpeg_7886_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_30),
.B1(n_21),
.B2(n_35),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_32),
.B1(n_16),
.B2(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_54),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_30),
.B1(n_19),
.B2(n_31),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_53),
.A2(n_29),
.A3(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_30),
.B1(n_21),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_76),
.B1(n_32),
.B2(n_29),
.Y(n_111)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_16),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_30),
.B1(n_21),
.B2(n_33),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_33),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_8),
.B(n_15),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_27),
.B1(n_16),
.B2(n_26),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_106),
.B1(n_34),
.B2(n_23),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_24),
.B1(n_20),
.B2(n_59),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_91),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_95),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_103),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_SL g136 ( 
.A(n_99),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_26),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_14),
.B(n_11),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_25),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_73),
.A3(n_51),
.B1(n_19),
.B2(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_27),
.B1(n_29),
.B2(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_75),
.Y(n_134)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_134),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_41),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_77),
.C(n_83),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_139),
.B1(n_96),
.B2(n_82),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_140),
.Y(n_150)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_132),
.Y(n_164)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_137),
.Y(n_180)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_59),
.B1(n_75),
.B2(n_24),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_89),
.A2(n_20),
.B1(n_34),
.B2(n_23),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_41),
.C(n_39),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_23),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_100),
.B1(n_106),
.B2(n_105),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_105),
.B1(n_91),
.B2(n_81),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_155),
.C(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_81),
.B1(n_90),
.B2(n_97),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_77),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_159),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_88),
.B1(n_92),
.B2(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_113),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_134),
.B1(n_140),
.B2(n_124),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_171),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_78),
.B1(n_80),
.B2(n_114),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_173),
.Y(n_201)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_23),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_78),
.B1(n_34),
.B2(n_19),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_19),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_34),
.B1(n_19),
.B2(n_9),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_135),
.B1(n_137),
.B2(n_126),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_126),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_1),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_122),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_183),
.C(n_188),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_119),
.C(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_189),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_117),
.B(n_145),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_202),
.B(n_177),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_130),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_208),
.C(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_191),
.B(n_192),
.Y(n_240)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_199),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_205),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_150),
.B(n_19),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_148),
.B1(n_175),
.B2(n_152),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_7),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_13),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_212),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_1),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_1),
.C(n_2),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_231),
.B1(n_236),
.B2(n_238),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_148),
.B1(n_156),
.B2(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_216),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_261)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_221),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_227),
.B(n_228),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_155),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_186),
.B(n_211),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_167),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_213),
.C(n_196),
.Y(n_250)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_241),
.B1(n_10),
.B2(n_3),
.Y(n_262)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_190),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_246),
.C(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_200),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_222),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_184),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_234),
.B(n_221),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_184),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_196),
.C(n_181),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_208),
.C(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_202),
.C(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_259),
.C(n_218),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_204),
.C(n_147),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_228),
.B1(n_217),
.B2(n_6),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_234),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_223),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_265),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_256),
.C(n_250),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_272),
.B(n_273),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_215),
.B1(n_224),
.B2(n_240),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_236),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_251),
.B(n_257),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_243),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_278),
.B(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_242),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_251),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_229),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_295),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_265),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_276),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_258),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_244),
.C(n_249),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_253),
.C(n_248),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_267),
.C(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_278),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_272),
.B1(n_277),
.B2(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_292),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_276),
.CI(n_271),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_305),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_275),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_275),
.B(n_261),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_310),
.C(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_233),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_316),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_247),
.B(n_233),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_299),
.B(n_298),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_302),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_301),
.B1(n_302),
.B2(n_307),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_289),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_300),
.CI(n_303),
.CON(n_321),
.SN(n_321)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_322),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_300),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_320),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_325),
.B(n_321),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_325),
.Y(n_334)
);

OAI31xp33_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_331),
.A3(n_329),
.B(n_328),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_326),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_10),
.Y(n_337)
);

OAI311xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_4),
.A3(n_6),
.B1(n_332),
.C1(n_324),
.Y(n_338)
);


endmodule