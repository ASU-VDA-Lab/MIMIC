module fake_jpeg_2782_n_699 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_699);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_699;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_5),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_63),
.Y(n_223)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_22),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_78),
.Y(n_149)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_22),
.A2(n_19),
.B1(n_17),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_68),
.A2(n_37),
.B1(n_28),
.B2(n_31),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_72),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_73),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_74),
.Y(n_205)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_76),
.Y(n_220)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_77),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_88),
.Y(n_156)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_82),
.Y(n_222)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_96),
.Y(n_214)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_113),
.Y(n_177)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_20),
.Y(n_108)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_59),
.Y(n_109)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_42),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_20),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_24),
.B(n_44),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_37),
.Y(n_184)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_53),
.Y(n_146)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_38),
.Y(n_130)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_23),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_132),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_28),
.B1(n_53),
.B2(n_25),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_143),
.A2(n_182),
.B1(n_212),
.B2(n_54),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_146),
.B(n_23),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_78),
.A2(n_34),
.B(n_44),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_147),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_SL g158 ( 
.A(n_115),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_97),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_161),
.B(n_166),
.C(n_174),
.Y(n_277)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_103),
.A2(n_40),
.B(n_34),
.C(n_31),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_165),
.A2(n_57),
.B(n_54),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_72),
.B(n_25),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_171),
.A2(n_175),
.B1(n_217),
.B2(n_225),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_112),
.B(n_26),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_173),
.B(n_184),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_104),
.B(n_53),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_64),
.A2(n_25),
.B1(n_40),
.B2(n_26),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_63),
.A2(n_25),
.B1(n_46),
.B2(n_33),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_60),
.B(n_46),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_191),
.B(n_208),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_120),
.B(n_41),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_41),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_102),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_99),
.B(n_32),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_209),
.B(n_0),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_71),
.A2(n_46),
.B1(n_41),
.B2(n_32),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_94),
.B(n_49),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_228),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_61),
.B(n_49),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_57),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_73),
.A2(n_48),
.B1(n_32),
.B2(n_33),
.Y(n_217)
);

BUFx16f_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g304 ( 
.A(n_218),
.Y(n_304)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_116),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_62),
.A2(n_49),
.B1(n_48),
.B2(n_33),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_96),
.B(n_48),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_127),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_234),
.B(n_239),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_235),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_236),
.Y(n_353)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_237),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g238 ( 
.A1(n_143),
.A2(n_77),
.B1(n_93),
.B2(n_82),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_238),
.A2(n_275),
.B1(n_276),
.B2(n_280),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_127),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_242),
.A2(n_245),
.B(n_273),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_74),
.B1(n_89),
.B2(n_65),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_246),
.A2(n_247),
.B1(n_267),
.B2(n_212),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_147),
.A2(n_70),
.B1(n_101),
.B2(n_98),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_150),
.Y(n_250)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_250),
.Y(n_342)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_162),
.Y(n_251)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_251),
.Y(n_369)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_149),
.A2(n_118),
.B1(n_117),
.B2(n_114),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_253),
.B(n_291),
.Y(n_349)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_181),
.Y(n_255)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_257),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_136),
.B(n_111),
.C(n_107),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_259),
.B(n_288),
.C(n_155),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_268),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_265),
.Y(n_368)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_266),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_156),
.A2(n_142),
.B1(n_177),
.B2(n_135),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_148),
.Y(n_270)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_168),
.Y(n_272)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_149),
.B(n_54),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_217),
.A2(n_106),
.B1(n_126),
.B2(n_125),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_164),
.A2(n_122),
.B1(n_67),
.B2(n_76),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_191),
.B(n_57),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_279),
.B(n_294),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_182),
.A2(n_130),
.B1(n_47),
.B2(n_81),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_202),
.Y(n_282)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_284),
.Y(n_334)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_151),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_166),
.B(n_47),
.Y(n_285)
);

AOI22x1_ASAP7_75t_L g351 ( 
.A1(n_285),
.A2(n_295),
.B1(n_176),
.B2(n_58),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_138),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_299),
.Y(n_320)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_197),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_287),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_144),
.B(n_90),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_172),
.A2(n_180),
.B1(n_187),
.B2(n_193),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_289),
.A2(n_229),
.B1(n_222),
.B2(n_205),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_203),
.A2(n_47),
.B1(n_45),
.B2(n_90),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_139),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_292),
.Y(n_364)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_194),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_137),
.B(n_85),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_176),
.A2(n_23),
.B(n_45),
.C(n_85),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_167),
.B(n_170),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_300),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_140),
.A2(n_45),
.B1(n_58),
.B2(n_16),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_298),
.A2(n_169),
.B1(n_133),
.B2(n_139),
.Y(n_335)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_207),
.B(n_15),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_206),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_305),
.Y(n_329)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_308),
.Y(n_358)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_159),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_192),
.B(n_15),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_310),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_178),
.B(n_14),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_158),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_311),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_197),
.B(n_229),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_316),
.B(n_319),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_218),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_248),
.A2(n_210),
.B1(n_134),
.B2(n_214),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_321),
.A2(n_362),
.B1(n_372),
.B2(n_308),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_254),
.B(n_221),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_323),
.B(n_344),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_260),
.A2(n_188),
.B1(n_190),
.B2(n_211),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_219),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_267),
.B(n_210),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_356),
.Y(n_414)
);

AOI32xp33_ASAP7_75t_L g350 ( 
.A1(n_268),
.A2(n_307),
.A3(n_277),
.B1(n_258),
.B2(n_253),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_274),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_361),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_276),
.A2(n_157),
.B1(n_195),
.B2(n_223),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_245),
.B(n_285),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_134),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_1),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_256),
.A2(n_157),
.B1(n_223),
.B2(n_154),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_285),
.A2(n_189),
.B(n_214),
.C(n_58),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_363),
.B(n_3),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_295),
.A2(n_222),
.B1(n_205),
.B2(n_58),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_371),
.A2(n_291),
.B(n_282),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_238),
.A2(n_246),
.B1(n_289),
.B2(n_259),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_288),
.B(n_58),
.C(n_14),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_306),
.C(n_284),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_230),
.B(n_298),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_378),
.A2(n_405),
.B(n_363),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_261),
.B1(n_257),
.B2(n_251),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_288),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_410),
.C(n_412),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_383),
.A2(n_362),
.B1(n_344),
.B2(n_355),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_316),
.A2(n_230),
.B1(n_305),
.B2(n_250),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_388),
.B1(n_403),
.B2(n_407),
.Y(n_434)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_347),
.A2(n_264),
.B1(n_262),
.B2(n_235),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_390),
.A2(n_392),
.B(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_319),
.Y(n_433)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_394),
.Y(n_442)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_357),
.B(n_241),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_SL g435 ( 
.A(n_395),
.B(n_319),
.Y(n_435)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_320),
.B(n_243),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_398),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_249),
.C(n_232),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_319),
.C(n_332),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_400),
.Y(n_458)
);

AO21x2_ASAP7_75t_SL g401 ( 
.A1(n_351),
.A2(n_244),
.B(n_236),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_401),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_372),
.A2(n_271),
.B1(n_293),
.B2(n_265),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_356),
.A2(n_349),
.B(n_345),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_278),
.B(n_301),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_334),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_406),
.B(n_409),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_333),
.A2(n_292),
.B1(n_263),
.B2(n_233),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_333),
.A2(n_255),
.B1(n_272),
.B2(n_287),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_408),
.A2(n_415),
.B1(n_426),
.B2(n_364),
.Y(n_431)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_304),
.C(n_240),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_314),
.B(n_13),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_423),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_323),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_349),
.A2(n_252),
.B1(n_240),
.B2(n_13),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_418),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_304),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_417),
.B(n_348),
.C(n_340),
.Y(n_457)
);

AO21x2_ASAP7_75t_L g419 ( 
.A1(n_321),
.A2(n_1),
.B(n_3),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_420),
.Y(n_437)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_1),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_332),
.B(n_304),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_348),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_338),
.B(n_370),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_349),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_404),
.B(n_337),
.CI(n_350),
.CON(n_427),
.SN(n_427)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_427),
.B(n_459),
.CI(n_393),
.CON(n_490),
.SN(n_490)
);

OAI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_430),
.A2(n_396),
.B1(n_391),
.B2(n_409),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_431),
.A2(n_445),
.B1(n_401),
.B2(n_405),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_433),
.B(n_435),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_436),
.A2(n_461),
.B(n_463),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_395),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_314),
.B1(n_338),
.B2(n_373),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_447),
.B1(n_453),
.B2(n_468),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_444),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_381),
.A2(n_338),
.B1(n_370),
.B2(n_355),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_374),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_452),
.C(n_455),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_383),
.A2(n_359),
.B1(n_358),
.B2(n_352),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_325),
.A3(n_365),
.B1(n_322),
.B2(n_359),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_322),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_381),
.A2(n_352),
.B1(n_339),
.B2(n_317),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_382),
.B(n_334),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_464),
.C(n_389),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_399),
.B(n_334),
.C(n_368),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_387),
.B(n_367),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g486 ( 
.A(n_460),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_381),
.A2(n_367),
.B(n_364),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_378),
.A2(n_346),
.B(n_324),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_410),
.B(n_340),
.C(n_331),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_389),
.A2(n_339),
.B1(n_330),
.B2(n_343),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_389),
.B1(n_408),
.B2(n_414),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_472),
.A2(n_481),
.B1(n_493),
.B2(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_413),
.Y(n_473)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_432),
.B(n_411),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_474),
.Y(n_534)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_466),
.Y(n_475)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_475),
.Y(n_528)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_478),
.A2(n_482),
.B1(n_484),
.B2(n_485),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_479),
.B(n_495),
.C(n_507),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_462),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_480),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_467),
.A2(n_413),
.B1(n_403),
.B2(n_407),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_401),
.B1(n_419),
.B2(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_434),
.A2(n_401),
.B1(n_402),
.B2(n_397),
.Y(n_484)
);

AOI22x1_ASAP7_75t_L g485 ( 
.A1(n_445),
.A2(n_397),
.B1(n_377),
.B2(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_492),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_430),
.A2(n_419),
.B1(n_415),
.B2(n_426),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_488),
.A2(n_496),
.B1(n_504),
.B2(n_505),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_489),
.B(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_449),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_443),
.A2(n_395),
.B1(n_419),
.B2(n_418),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_441),
.B(n_422),
.C(n_423),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_456),
.A2(n_377),
.B1(n_379),
.B2(n_431),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_463),
.A2(n_419),
.B1(n_388),
.B2(n_421),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_499),
.B(n_502),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_500),
.A2(n_442),
.B1(n_394),
.B2(n_369),
.Y(n_533)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_439),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_501),
.B(n_442),
.Y(n_532)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_447),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_437),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_459),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_437),
.A2(n_386),
.B1(n_420),
.B2(n_400),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_434),
.A2(n_461),
.B1(n_465),
.B2(n_468),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_441),
.B(n_331),
.C(n_328),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_433),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_509),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_446),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_452),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_519),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_492),
.A2(n_428),
.B1(n_453),
.B2(n_427),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_512),
.A2(n_514),
.B1(n_529),
.B2(n_530),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_497),
.A2(n_428),
.B1(n_427),
.B2(n_429),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_486),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_522),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_489),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_505),
.A2(n_444),
.B1(n_429),
.B2(n_450),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_521),
.A2(n_523),
.B1(n_533),
.B2(n_496),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_469),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_502),
.A2(n_457),
.B1(n_455),
.B2(n_458),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_525),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_506),
.A2(n_435),
.B(n_464),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_527),
.A2(n_475),
.B(n_342),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_497),
.A2(n_458),
.B1(n_448),
.B2(n_440),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_503),
.A2(n_439),
.B1(n_442),
.B2(n_416),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_507),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_543),
.C(n_487),
.Y(n_547)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_532),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_330),
.Y(n_535)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_369),
.Y(n_537)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_537),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_342),
.Y(n_538)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_538),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_476),
.B(n_491),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_477),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_494),
.B(n_470),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_541),
.B(n_353),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_491),
.B(n_346),
.C(n_328),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_469),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_488),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_478),
.A2(n_343),
.B1(n_353),
.B2(n_366),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_484),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_547),
.B(n_567),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_548),
.A2(n_562),
.B1(n_574),
.B2(n_528),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_520),
.Y(n_549)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_549),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_517),
.B(n_508),
.C(n_509),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_550),
.B(n_552),
.C(n_555),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_517),
.B(n_472),
.C(n_490),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_511),
.C(n_519),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_526),
.A2(n_482),
.B1(n_498),
.B2(n_504),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_556),
.A2(n_568),
.B(n_7),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_539),
.B(n_490),
.C(n_483),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_557),
.B(n_561),
.C(n_566),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_481),
.Y(n_559)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_559),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_563),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_493),
.C(n_485),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_501),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_485),
.C(n_506),
.Y(n_566)
);

XNOR2x1_ASAP7_75t_L g569 ( 
.A(n_525),
.B(n_366),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_569),
.B(n_575),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_514),
.B(n_512),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_570),
.B(n_513),
.Y(n_583)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_573),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_513),
.A2(n_318),
.B1(n_4),
.B2(n_5),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g575 ( 
.A(n_510),
.B(n_318),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_534),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_579),
.Y(n_584)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_540),
.Y(n_578)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_578),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_535),
.B(n_3),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_516),
.B(n_3),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_6),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_583),
.B(n_587),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_554),
.A2(n_572),
.B1(n_521),
.B2(n_515),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_585),
.A2(n_591),
.B1(n_598),
.B2(n_548),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_515),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_565),
.B(n_510),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_599),
.Y(n_618)
);

OAI22x1_ASAP7_75t_L g591 ( 
.A1(n_554),
.A2(n_533),
.B1(n_542),
.B2(n_524),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_543),
.C(n_524),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_593),
.B(n_594),
.C(n_596),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_558),
.B(n_516),
.C(n_537),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_547),
.B(n_546),
.C(n_536),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_572),
.A2(n_540),
.B1(n_545),
.B2(n_528),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_565),
.B(n_545),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_600),
.A2(n_605),
.B1(n_579),
.B2(n_571),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_566),
.A2(n_538),
.B(n_318),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_601),
.A2(n_602),
.B(n_576),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_553),
.A2(n_3),
.B(n_5),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_555),
.B(n_5),
.C(n_6),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_603),
.B(n_601),
.C(n_576),
.Y(n_625)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_604),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_562),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_607),
.A2(n_568),
.B1(n_551),
.B2(n_578),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_608),
.A2(n_614),
.B1(n_622),
.B2(n_8),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_609),
.Y(n_631)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_592),
.Y(n_610)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_598),
.Y(n_611)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_611),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_612),
.A2(n_605),
.B1(n_583),
.B2(n_588),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_551),
.Y(n_613)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_613),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_597),
.B(n_570),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_615),
.B(n_603),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_585),
.A2(n_561),
.B(n_564),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_616),
.A2(n_628),
.B(n_7),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_SL g617 ( 
.A(n_590),
.B(n_575),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_617),
.B(n_623),
.Y(n_637)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_595),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_621),
.Y(n_634)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_600),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_591),
.A2(n_559),
.B1(n_564),
.B2(n_571),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_593),
.B(n_567),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_582),
.B(n_557),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_624),
.B(n_8),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_625),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_626),
.B(n_630),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_588),
.A2(n_569),
.B(n_587),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g630 ( 
.A1(n_584),
.A2(n_552),
.B1(n_574),
.B2(n_9),
.C(n_10),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_623),
.Y(n_657)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_633),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_616),
.A2(n_589),
.B(n_602),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_635),
.A2(n_640),
.B(n_629),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_612),
.A2(n_589),
.B1(n_594),
.B2(n_596),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_641),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_620),
.B(n_586),
.C(n_599),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_638),
.B(n_620),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_611),
.A2(n_582),
.B(n_586),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_609),
.B(n_7),
.Y(n_641)
);

OAI21x1_ASAP7_75t_SL g664 ( 
.A1(n_643),
.A2(n_9),
.B(n_10),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_644),
.B(n_625),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_8),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_646),
.B(n_647),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_613),
.B(n_8),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_650),
.A2(n_628),
.B1(n_627),
.B2(n_626),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_639),
.A2(n_621),
.B1(n_619),
.B2(n_610),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_651),
.B(n_652),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_653),
.B(n_654),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_649),
.B(n_635),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_657),
.B(n_659),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_658),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_638),
.B(n_629),
.C(n_618),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_660),
.A2(n_643),
.B(n_634),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_650),
.A2(n_622),
.B1(n_608),
.B2(n_617),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_661),
.B(n_662),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_9),
.C(n_10),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_664),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_639),
.A2(n_9),
.B1(n_648),
.B2(n_645),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_665),
.B(n_642),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_636),
.B(n_9),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_666),
.B(n_641),
.Y(n_667)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_667),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_659),
.B(n_648),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_670),
.B(n_673),
.Y(n_682)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_671),
.Y(n_686)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_633),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_672),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_656),
.B(n_645),
.C(n_631),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_674),
.B(n_653),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_674),
.B(n_656),
.C(n_655),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_679),
.B(n_683),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_669),
.B(n_631),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_684),
.A2(n_685),
.B(n_668),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_655),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_682),
.A2(n_675),
.B(n_676),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_687),
.A2(n_691),
.B(n_677),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_673),
.B(n_672),
.Y(n_688)
);

OAI211xp5_ASAP7_75t_L g694 ( 
.A1(n_688),
.A2(n_689),
.B(n_663),
.C(n_647),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_681),
.A2(n_634),
.B(n_642),
.Y(n_691)
);

A2O1A1O1Ixp25_ASAP7_75t_L g692 ( 
.A1(n_690),
.A2(n_679),
.B(n_686),
.C(n_680),
.D(n_662),
.Y(n_692)
);

AO21x1_ASAP7_75t_L g696 ( 
.A1(n_692),
.A2(n_693),
.B(n_694),
.Y(n_696)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_693),
.B(n_661),
.C(n_637),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_695),
.B(n_632),
.C(n_663),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_697),
.A2(n_696),
.B(n_637),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_698),
.B(n_646),
.Y(n_699)
);


endmodule