module fake_jpeg_10712_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.C(n_45),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_46),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_87),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_42),
.B1(n_51),
.B2(n_54),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_1),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_67),
.C(n_72),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_5),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_6),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_95),
.C(n_16),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_106),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_22),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_102),
.C(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_106),
.B(n_92),
.Y(n_112)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_105),
.Y(n_110)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_10),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_11),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_15),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_105),
.B1(n_101),
.B2(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_116),
.B1(n_113),
.B2(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_115),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_123),
.A2(n_120),
.B(n_117),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_122),
.A3(n_107),
.B1(n_123),
.B2(n_24),
.C1(n_26),
.C2(n_28),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_124),
.C(n_20),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_19),
.A3(n_21),
.B1(n_29),
.B2(n_30),
.C1(n_31),
.C2(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_35),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_36),
.Y(n_130)
);


endmodule