module real_jpeg_26501_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_0),
.A2(n_52),
.B(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_0),
.A2(n_26),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_26),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_41),
.B1(n_47),
.B2(n_107),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_21),
.Y(n_42)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_5),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_30),
.Y(n_107)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_22),
.A3(n_26),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_83),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_81),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_48),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_15),
.B(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_38),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_29),
.B2(n_31),
.Y(n_16)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_17),
.A2(n_18),
.B1(n_29),
.B2(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_25),
.Y(n_17)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_18),
.B(n_57),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_20),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_21),
.B(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_26),
.B(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_27),
.A2(n_52),
.A3(n_56),
.B1(n_59),
.B2(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_51),
.B1(n_58),
.B2(n_62),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_52),
.B(n_59),
.C(n_61),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_38),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_43),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_41),
.A2(n_45),
.B1(n_101),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_42),
.A2(n_46),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_97),
.B(n_116),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_104),
.B(n_115),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_103),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_114),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);


endmodule