module real_jpeg_4174_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_1),
.A2(n_43),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_43),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_43),
.B1(n_174),
.B2(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_21),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_5),
.Y(n_308)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_6),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_53),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_53),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_127),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_10),
.A2(n_250),
.B(n_253),
.C(n_257),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_10),
.B(n_28),
.C(n_63),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_10),
.B(n_81),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_10),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_10),
.B(n_69),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_134),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_11),
.A2(n_134),
.B1(n_264),
.B2(n_267),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_11),
.A2(n_71),
.B1(n_134),
.B2(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_217),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_215),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_192),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_16),
.B(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.C(n_176),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_17),
.B(n_176),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_18),
.B(n_110),
.C(n_139),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_45),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_19),
.B(n_45),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_36),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_20),
.A2(n_147),
.B(n_150),
.Y(n_146)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_25),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_31),
.B(n_40),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_31),
.A2(n_180),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_31),
.B(n_180),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_31),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_32),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g182 ( 
.A(n_33),
.Y(n_182)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_33),
.Y(n_287)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_36),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_36),
.B(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_39),
.Y(n_149)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_73),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_46),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_47),
.Y(n_242)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_51),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_51),
.Y(n_266)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_53),
.B(n_136),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_53),
.A2(n_113),
.B(n_159),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_53),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_56),
.B(n_74),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_56),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_56),
.B(n_263),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_59),
.Y(n_256)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_69),
.B(n_263),
.Y(n_278)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_71),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_73),
.A2(n_186),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_73),
.B(n_262),
.Y(n_289)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_76),
.Y(n_275)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_110),
.B1(n_139),
.B2(n_140),
.Y(n_79)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_93),
.B(n_105),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_81),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_81),
.B(n_169),
.Y(n_239)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_82),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_86),
.Y(n_252)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_93),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_93),
.B(n_105),
.Y(n_205)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_94),
.B(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_105),
.Y(n_167)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_106),
.Y(n_257)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_131),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_127),
.Y(n_143)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_118),
.B(n_200),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_127),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_131),
.B(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_141),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_164),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_142),
.B(n_164),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_145),
.B(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_146),
.B(n_151),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_155),
.A3(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_202),
.Y(n_224)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_184),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_178),
.B(n_281),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_183),
.B(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B(n_191),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_185),
.A2(n_212),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_185),
.B(n_242),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_191),
.B(n_278),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_192),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_206),
.CI(n_214),
.CON(n_192),
.SN(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_205),
.B(n_239),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_207),
.A2(n_213),
.B1(n_249),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_333),
.B(n_346),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_268),
.B(n_332),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_244),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_220),
.B(n_244),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_223),
.B(n_229),
.C(n_231),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_232),
.B(n_235),
.C(n_241),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_258),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_248),
.A2(n_258),
.B1(n_259),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_326),
.B(n_331),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_316),
.B(n_325),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_293),
.B(n_315),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_279),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_274),
.B1(n_277),
.B2(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_300),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_290),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_291),
.C(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_302),
.B(n_314),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_297),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_310),
.B(n_313),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_319),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.C(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_330),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_342),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_336),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_342),
.A2(n_347),
.B(n_348),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_345),
.Y(n_348)
);


endmodule