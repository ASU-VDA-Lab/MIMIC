module fake_jpeg_6343_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_20),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_23),
.B(n_20),
.C(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_55),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_65),
.B1(n_53),
.B2(n_19),
.Y(n_98)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_66),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_23),
.B(n_29),
.C(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_60),
.B1(n_52),
.B2(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_19),
.B1(n_17),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_73),
.B1(n_83),
.B2(n_7),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_22),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_22),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_18),
.B1(n_21),
.B2(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_18),
.B1(n_21),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_25),
.B1(n_22),
.B2(n_43),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_30),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_20),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_20),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_29),
.B1(n_19),
.B2(n_25),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_49),
.B1(n_53),
.B2(n_45),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_31),
.B(n_25),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_100),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_50),
.B1(n_57),
.B2(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_104),
.B1(n_85),
.B2(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_106),
.B1(n_111),
.B2(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_61),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_45),
.B1(n_53),
.B2(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_45),
.B1(n_20),
.B2(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_90),
.B1(n_94),
.B2(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_125),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_101),
.B1(n_114),
.B2(n_112),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_77),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_137),
.B(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_132),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_61),
.B(n_77),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_139),
.B(n_113),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_131),
.B1(n_133),
.B2(n_95),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_87),
.B1(n_69),
.B2(n_85),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_73),
.B1(n_72),
.B2(n_74),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_87),
.B1(n_69),
.B2(n_80),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_69),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_70),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_90),
.B1(n_104),
.B2(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_144),
.B1(n_152),
.B2(n_3),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_157),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_111),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_137),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_103),
.B1(n_95),
.B2(n_93),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_107),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_116),
.B1(n_115),
.B2(n_121),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_137),
.Y(n_176)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_168),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_171),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_63),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_93),
.C(n_9),
.Y(n_186)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_174),
.B(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_142),
.B1(n_131),
.B2(n_117),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_139),
.B(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_180),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_158),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_123),
.B1(n_125),
.B2(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_188),
.C(n_170),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_9),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

OR2x6_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_3),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_156),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_196),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_155),
.B1(n_156),
.B2(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_152),
.B1(n_143),
.B2(n_179),
.Y(n_219)
);

XNOR2x2_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_166),
.Y(n_198)
);

AOI321xp33_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_203),
.A3(n_206),
.B1(n_208),
.B2(n_210),
.C(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_213),
.C(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_164),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_147),
.C(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_157),
.C(n_161),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_191),
.B1(n_174),
.B2(n_192),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_217),
.B1(n_212),
.B2(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_197),
.B1(n_201),
.B2(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_150),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_233),
.B(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_229),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_213),
.C(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_231),
.C(n_210),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_175),
.C(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_151),
.B1(n_167),
.B2(n_189),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_183),
.B1(n_196),
.B2(n_189),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_241),
.B(n_15),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_238),
.B1(n_245),
.B2(n_4),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_242),
.C(n_244),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_224),
.B1(n_228),
.B2(n_148),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_212),
.B(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_206),
.C(n_208),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_243),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_215),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_144),
.B1(n_148),
.B2(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_248),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_230),
.C(n_231),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_218),
.B(n_225),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_254),
.B(n_8),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_229),
.C(n_171),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_15),
.B1(n_8),
.B2(n_11),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_237),
.B1(n_243),
.B2(n_239),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_237),
.B1(n_12),
.B2(n_7),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_262),
.B(n_11),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_8),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_253),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_267),
.B(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_262),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_13),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_272),
.B(n_273),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_13),
.B1(n_14),
.B2(n_5),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_269),
.B(n_5),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_5),
.B(n_6),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_5),
.Y(n_279)
);


endmodule