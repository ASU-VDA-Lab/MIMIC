module fake_jpeg_22020_n_244 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_19),
.B1(n_33),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_43),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.C(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_21),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_25),
.B1(n_23),
.B2(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_42),
.B1(n_19),
.B2(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_30),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_23),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_77),
.B1(n_51),
.B2(n_26),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_23),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_38),
.B1(n_19),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_72),
.B1(n_55),
.B2(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_28),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_73),
.B(n_22),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_43),
.B1(n_34),
.B2(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_21),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_95),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_63),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_40),
.B(n_58),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_75),
.B(n_64),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_29),
.A3(n_54),
.B1(n_18),
.B2(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_108),
.B1(n_91),
.B2(n_84),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_61),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_110),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_111),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_59),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_69),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_113),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_89),
.C(n_92),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_128),
.C(n_109),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_99),
.B1(n_86),
.B2(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_136),
.B1(n_107),
.B2(n_67),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_92),
.C(n_99),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_133),
.B1(n_135),
.B2(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_98),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_105),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_101),
.B1(n_113),
.B2(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_111),
.B(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_95),
.B1(n_88),
.B2(n_78),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_88),
.B1(n_78),
.B2(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_117),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_148),
.C(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_124),
.C(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_134),
.B1(n_70),
.B2(n_54),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_120),
.C(n_104),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_62),
.B(n_104),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_139),
.B(n_127),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_64),
.B(n_120),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_140),
.C(n_141),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_0),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_175),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_126),
.B(n_134),
.C(n_123),
.D(n_125),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_144),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_177),
.B1(n_14),
.B2(n_7),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_70),
.B1(n_18),
.B2(n_16),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_14),
.B(n_70),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_18),
.B(n_14),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_162),
.B1(n_151),
.B2(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_156),
.B1(n_149),
.B2(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_142),
.C(n_148),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_191),
.C(n_193),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_188),
.B(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_5),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_161),
.B(n_24),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_166),
.B(n_177),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_6),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_165),
.B1(n_167),
.B2(n_180),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_185),
.B1(n_181),
.B2(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_203),
.A2(n_199),
.B1(n_206),
.B2(n_205),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_172),
.C(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_163),
.C(n_180),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_5),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_7),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_7),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_213),
.C(n_4),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_0),
.C(n_1),
.Y(n_213)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_216),
.A2(n_201),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_4),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_202),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_11),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_218),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

AOI21x1_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_210),
.B(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_226),
.B(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_222),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_229),
.B(n_230),
.C(n_209),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_219),
.B(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_12),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_4),
.B1(n_10),
.B2(n_11),
.Y(n_238)
);

OAI311xp33_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.C1(n_2),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_242),
.A2(n_239),
.B(n_13),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_1),
.Y(n_244)
);


endmodule