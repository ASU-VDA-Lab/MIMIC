module real_jpeg_12517_n_16 (n_383, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_383;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_68),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_45),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_28),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_4),
.B(n_45),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_4),
.B(n_33),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_4),
.B(n_61),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_4),
.B(n_35),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_40),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_33),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_28),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_61),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_54),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_7),
.B(n_61),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_7),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_7),
.B(n_68),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_7),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_7),
.B(n_54),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_33),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_8),
.B(n_45),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_11),
.B(n_68),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_11),
.B(n_61),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_45),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_33),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_11),
.B(n_35),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_11),
.B(n_54),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_11),
.B(n_40),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_13),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_13),
.B(n_54),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_13),
.B(n_61),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_35),
.Y(n_165)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_15),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_15),
.B(n_28),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_45),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_147),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_97),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_21),
.B(n_81),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_23),
.B(n_49),
.C(n_57),
.Y(n_146)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.C(n_43),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_25),
.A2(n_26),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.C(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_27),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_120),
.C(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_27),
.A2(n_112),
.B1(n_120),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_27),
.A2(n_112),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_27),
.B(n_193),
.Y(n_209)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_28),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_29),
.A2(n_30),
.B1(n_67),
.B2(n_70),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_29),
.B(n_67),
.C(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_32),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_32),
.B(n_78),
.Y(n_319)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_34),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_34),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_34),
.A2(n_110),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_37),
.A2(n_43),
.B1(n_44),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_39),
.B(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_39),
.B(n_232),
.Y(n_303)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_66),
.C(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_43),
.A2(n_44),
.B1(n_122),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_43),
.A2(n_44),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_44),
.B(n_119),
.C(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_44),
.B(n_213),
.Y(n_267)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_46),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_46),
.B(n_232),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_51),
.B(n_53),
.C(n_55),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_54),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_72),
.C(n_79),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_59),
.A2(n_60),
.B1(n_106),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_106),
.C(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_66),
.C(n_67),
.Y(n_128)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_65),
.A2(n_66),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_66),
.B(n_253),
.C(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_67),
.A2(n_70),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx5_ASAP7_75t_SL g201 ( 
.A(n_68),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.C(n_76),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_74),
.B(n_191),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_77),
.B(n_189),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_80),
.A2(n_86),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_80),
.B(n_141),
.C(n_315),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.C(n_92),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_87),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_89),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_90),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_90),
.B(n_201),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_93),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_114),
.C(n_118),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_98),
.A2(n_99),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_101),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_106),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_107),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_120),
.A2(n_163),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_120),
.B(n_260),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_146),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_144),
.B2(n_145),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_140),
.A2(n_141),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_175),
.B(n_379),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_173),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_150),
.B(n_173),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_166),
.C(n_170),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_151),
.B(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_160),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_152),
.A2(n_153),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_157),
.B(n_160),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_161),
.B(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_164),
.A2(n_165),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_164),
.Y(n_352)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_165),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_166),
.B(n_170),
.Y(n_372)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI321xp33_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_359),
.A3(n_369),
.B1(n_373),
.B2(n_378),
.C(n_383),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_306),
.C(n_354),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_277),
.B(n_305),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_247),
.B(n_276),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_216),
.B(n_246),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_181),
.B(n_195),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_192),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_198),
.B1(n_199),
.B2(n_207),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_182),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_243),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.CI(n_185),
.CON(n_182),
.SN(n_182)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_186),
.A2(n_187),
.B1(n_192),
.B2(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_188),
.B(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_208),
.B2(n_215),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_207),
.C(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_203),
.C(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_205),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_213),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_213),
.A2(n_214),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_213),
.B(n_327),
.C(n_330),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_240),
.B(n_245),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_229),
.B(n_239),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_227),
.C(n_228),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_234),
.B(n_238),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_249),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_262),
.B2(n_263),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_264),
.C(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_274),
.B2(n_275),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_273),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_270),
.C(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_269),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_278),
.B(n_279),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_295),
.B2(n_304),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_294),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_294),
.C(n_304),
.Y(n_355)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_292),
.C(n_293),
.Y(n_323)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_286),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.CI(n_289),
.CON(n_286),
.SN(n_286)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_295),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.CI(n_301),
.CON(n_295),
.SN(n_295)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_297),
.C(n_301),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B(n_300),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_300),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g374 ( 
.A1(n_307),
.A2(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_336),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_308),
.B(n_336),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_324),
.C(n_335),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_323),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_316),
.C(n_323),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_320),
.C(n_322),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_325),
.B1(n_335),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_332),
.C(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_329),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_353),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_345),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_345),
.C(n_353),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_343),
.C(n_344),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_348),
.C(n_349),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_356),
.Y(n_375)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_360),
.A2(n_374),
.B(n_377),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_361),
.B(n_362),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_368),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.C(n_368),
.Y(n_370)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_371),
.Y(n_378)
);


endmodule