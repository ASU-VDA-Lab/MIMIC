module fake_netlist_1_2458_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g3 ( .A(n_2), .B(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
AND2x2_ASAP7_75t_L g5 ( .A(n_0), .B(n_1), .Y(n_5) );
INVx3_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_3), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx3_ASAP7_75t_SL g11 ( .A(n_8), .Y(n_11) );
NAND3xp33_ASAP7_75t_SL g12 ( .A(n_10), .B(n_3), .C(n_7), .Y(n_12) );
NAND4xp25_ASAP7_75t_SL g13 ( .A(n_11), .B(n_1), .C(n_6), .D(n_8), .Y(n_13) );
OAI21xp5_ASAP7_75t_SL g14 ( .A1(n_12), .A2(n_11), .B(n_6), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_13), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_14), .B(n_6), .Y(n_17) );
endmodule