module fake_jpeg_22895_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_22),
.Y(n_59)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_47),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_16),
.C(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_21),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_45),
.B1(n_36),
.B2(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_29),
.B1(n_17),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_45),
.B1(n_36),
.B2(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_16),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_44),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_61),
.C(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_81),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_66),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_82),
.B1(n_96),
.B2(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_34),
.Y(n_115)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_37),
.B1(n_35),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_91),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_97),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_106),
.B(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_107),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_67),
.B1(n_76),
.B2(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_61),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_36),
.B1(n_39),
.B2(n_67),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_43),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_123),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_66),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_53),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_53),
.B1(n_110),
.B2(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_137),
.B1(n_144),
.B2(n_146),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_140),
.Y(n_158)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_74),
.B1(n_92),
.B2(n_87),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_80),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_106),
.B1(n_107),
.B2(n_100),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_36),
.B1(n_45),
.B2(n_79),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_150),
.B1(n_119),
.B2(n_110),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_52),
.B(n_56),
.C(n_102),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_82),
.B1(n_86),
.B2(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_157),
.B(n_170),
.Y(n_187)
);

OR2x2_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_71),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_175),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_24),
.B(n_32),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_40),
.B(n_43),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_171),
.B(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_165),
.B1(n_166),
.B2(n_150),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_71),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_174),
.C(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_119),
.B1(n_97),
.B2(n_104),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_71),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_24),
.B(n_32),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_57),
.B(n_24),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_137),
.B(n_140),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_52),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_94),
.B1(n_91),
.B2(n_118),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_196),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_128),
.B1(n_149),
.B2(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_188),
.B1(n_203),
.B2(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_145),
.B1(n_135),
.B2(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_192),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_138),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_200),
.B1(n_32),
.B2(n_112),
.Y(n_219)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_139),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_111),
.B1(n_108),
.B2(n_130),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_154),
.B1(n_108),
.B2(n_153),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_130),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_130),
.B(n_175),
.C(n_156),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_111),
.B1(n_90),
.B2(n_91),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_207),
.B1(n_219),
.B2(n_179),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_205),
.A2(n_20),
.B(n_28),
.C(n_25),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_171),
.B(n_157),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_222),
.B(n_17),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_173),
.C(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_218),
.C(n_227),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_154),
.B1(n_159),
.B2(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_164),
.B1(n_136),
.B2(n_170),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_216),
.B1(n_200),
.B2(n_199),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_118),
.B1(n_125),
.B2(n_90),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_56),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_95),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_225),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_25),
.B(n_28),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_202),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_95),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_94),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_203),
.B1(n_197),
.B2(n_193),
.Y(n_234)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_235),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_183),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_182),
.C(n_185),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_194),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_251),
.B(n_252),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_214),
.B1(n_225),
.B2(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_247),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_183),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_27),
.B(n_18),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_210),
.B(n_195),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_248),
.B1(n_33),
.B2(n_30),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_186),
.C(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_20),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_125),
.C(n_77),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_204),
.B1(n_216),
.B2(n_209),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_260),
.B1(n_272),
.B2(n_0),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_205),
.B(n_223),
.Y(n_257)
);

OAI22x1_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_251),
.B1(n_232),
.B2(n_18),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_205),
.B1(n_219),
.B2(n_125),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_77),
.B1(n_25),
.B2(n_26),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_77),
.B1(n_26),
.B2(n_40),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_40),
.B1(n_33),
.B2(n_30),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_0),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_231),
.A2(n_0),
.B(n_1),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_239),
.C(n_263),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_SL g299 ( 
.A(n_273),
.B(n_278),
.C(n_266),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_269),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_248),
.C(n_242),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_282),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_245),
.C(n_242),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_281),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_232),
.B1(n_1),
.B2(n_2),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_287),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_15),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_268),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_267),
.C(n_254),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_292),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_270),
.C(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_294),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_298),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_14),
.B(n_13),
.C(n_12),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_256),
.C(n_271),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_304),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_271),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_280),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_311),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_283),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_11),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_310),
.B1(n_291),
.B2(n_303),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_11),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_3),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_3),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_4),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_301),
.C(n_4),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_325),
.C(n_308),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_324),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_11),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_9),
.C(n_6),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_314),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_328),
.B(n_5),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_331),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_318),
.C(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_307),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_310),
.B(n_6),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_326),
.C(n_332),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_5),
.B(n_6),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_9),
.C(n_7),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_7),
.C(n_8),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_7),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_8),
.B(n_326),
.Y(n_343)
);


endmodule