module fake_netlist_6_4376_n_1556 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1556);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1556;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_290),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_15),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_38),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_20),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_73),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_99),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_247),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_51),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_22),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_231),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_4),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_256),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_119),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_318),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_127),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_80),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_199),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_68),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_88),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_6),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_297),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_251),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_91),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_59),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_21),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_225),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_58),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_222),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_46),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_22),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_283),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_84),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_125),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_262),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_193),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_124),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_9),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_108),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_157),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_216),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_58),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_298),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_200),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_142),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_106),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_232),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_52),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_55),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_156),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_315),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_183),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_299),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_205),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_192),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_308),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_202),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_239),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_147),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_249),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_295),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_213),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_53),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_116),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_169),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_162),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_40),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_61),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_209),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_300),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_43),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_196),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_112),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_120),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_173),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_329),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_100),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_59),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_69),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_49),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_271),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_267),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_228),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_265),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_1),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_195),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_7),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_223),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_122),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_76),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_210),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_47),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_113),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_5),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_21),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_4),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_178),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_79),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_52),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_92),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_240),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_185),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_266),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_207),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_307),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_201),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_96),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_78),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_288),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_97),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_327),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_194),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_204),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_171),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_273),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_51),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_31),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_161),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_55),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_114),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_166),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_244),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_321),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_18),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_280),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_20),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_259),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_139),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_6),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_155),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_74),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_151),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_93),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_80),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_165),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_326),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_30),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_101),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_0),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_291),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_158),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_168),
.Y(n_484)
);

INVx4_ASAP7_75t_R g485 ( 
.A(n_148),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_160),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_163),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_3),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_257),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_164),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_83),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_190),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_174),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_40),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_14),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_292),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_261),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_184),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_24),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_129),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_203),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_226),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_126),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_144),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_121),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_179),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_272),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_237),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_15),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_322),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_238),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_0),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_320),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_313),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_277),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_242),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_63),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_149),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_135),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_74),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_117),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_317),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_304),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_110),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_8),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_45),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_104),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_217),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_154),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_182),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_314),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_90),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_268),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_10),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_34),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_49),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_72),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_330),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_234),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_293),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_76),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_19),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_105),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_64),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_109),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_309),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_319),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_218),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_279),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_316),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_310),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_269),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_62),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_191),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_197),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_145),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_70),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_306),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_393),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_378),
.B(n_552),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_342),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_404),
.B(n_1),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_378),
.B(n_2),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_393),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_342),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_2),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_393),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_404),
.B(n_3),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_393),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_342),
.B(n_7),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_355),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_342),
.B(n_8),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_499),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_342),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_396),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_342),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_499),
.B(n_10),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_342),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_396),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_436),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_461),
.B(n_11),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_388),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_436),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_334),
.B(n_11),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_12),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_436),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_539),
.B(n_12),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_334),
.B(n_13),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_340),
.B(n_13),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_340),
.B(n_14),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_381),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_388),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_396),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_541),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_394),
.B(n_16),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_396),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_333),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_348),
.B(n_16),
.Y(n_600)
);

BUFx8_ASAP7_75t_SL g601 ( 
.A(n_491),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_454),
.B(n_17),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_429),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_429),
.Y(n_604)
);

BUFx12f_ASAP7_75t_L g605 ( 
.A(n_388),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_429),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_360),
.B(n_17),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_348),
.B(n_18),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_472),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_339),
.B(n_458),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_394),
.B(n_23),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_406),
.B(n_23),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_472),
.B(n_85),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_336),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_392),
.B(n_24),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_525),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_472),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_338),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_398),
.B(n_443),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_398),
.B(n_25),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_345),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_472),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_338),
.Y(n_625)
);

BUFx12f_ASAP7_75t_L g626 ( 
.A(n_525),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_333),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_366),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_353),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_443),
.B(n_25),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_525),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_414),
.B(n_26),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_545),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_515),
.B(n_26),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_353),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_364),
.Y(n_636)
);

CKINVDCx11_ASAP7_75t_R g637 ( 
.A(n_338),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_515),
.B(n_27),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_422),
.B(n_27),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_451),
.B(n_28),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_545),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_494),
.B(n_28),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_29),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_377),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_494),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_389),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_354),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_383),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_383),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_419),
.Y(n_652)
);

BUFx12f_ASAP7_75t_L g653 ( 
.A(n_383),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_418),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_530),
.B(n_29),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_418),
.B(n_30),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_444),
.B(n_457),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_418),
.B(n_31),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_503),
.B(n_32),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_448),
.B(n_32),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_420),
.B(n_33),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_375),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_376),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_379),
.B(n_33),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_520),
.B(n_34),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_428),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_385),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_437),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_520),
.B(n_35),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_441),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_448),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_386),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_448),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_387),
.B(n_391),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_468),
.Y(n_675)
);

BUFx12f_ASAP7_75t_L g676 ( 
.A(n_337),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_347),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_399),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_471),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_488),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_401),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_517),
.Y(n_682)
);

INVx6_ASAP7_75t_L g683 ( 
.A(n_357),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_537),
.B(n_36),
.Y(n_684)
);

BUFx12f_ASAP7_75t_L g685 ( 
.A(n_361),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_489),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_528),
.B(n_36),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_403),
.B(n_86),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_331),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_405),
.B(n_37),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_410),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_482),
.B(n_37),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_362),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_526),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_535),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_485),
.Y(n_696)
);

BUFx8_ASAP7_75t_SL g697 ( 
.A(n_489),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_332),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_423),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_536),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_502),
.B(n_38),
.Y(n_701)
);

BUFx12f_ASAP7_75t_L g702 ( 
.A(n_367),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_427),
.B(n_39),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_368),
.B(n_39),
.Y(n_704)
);

BUFx12f_ASAP7_75t_L g705 ( 
.A(n_369),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_416),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_335),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_408),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_409),
.B(n_41),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_430),
.B(n_41),
.Y(n_710)
);

BUFx12f_ASAP7_75t_L g711 ( 
.A(n_412),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_442),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_453),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_462),
.B(n_42),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_654),
.B(n_555),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_587),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_588),
.A2(n_483),
.B1(n_486),
.B2(n_465),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_574),
.B(n_696),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_657),
.A2(n_508),
.B1(n_531),
.B2(n_504),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_696),
.B(n_657),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_642),
.A2(n_426),
.B1(n_432),
.B2(n_421),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_588),
.A2(n_501),
.B1(n_511),
.B2(n_498),
.Y(n_722)
);

XNOR2xp5_ASAP7_75t_L g723 ( 
.A(n_628),
.B(n_540),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_614),
.A2(n_549),
.B1(n_438),
.B2(n_440),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_600),
.A2(n_450),
.B1(n_459),
.B2(n_434),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_572),
.A2(n_473),
.B1(n_476),
.B2(n_466),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_696),
.B(n_341),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_686),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_676),
.B(n_513),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_656),
.A2(n_532),
.B1(n_533),
.B2(n_521),
.Y(n_730)
);

BUFx6f_ASAP7_75t_SL g731 ( 
.A(n_620),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_692),
.A2(n_481),
.B1(n_495),
.B2(n_479),
.Y(n_732)
);

INVx8_ASAP7_75t_L g733 ( 
.A(n_706),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_654),
.B(n_509),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_582),
.A2(n_534),
.B1(n_544),
.B2(n_512),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_696),
.B(n_343),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_677),
.B(n_344),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_658),
.A2(n_547),
.B1(n_44),
.B2(n_42),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_609),
.A2(n_557),
.B1(n_553),
.B2(n_349),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_578),
.A2(n_350),
.B1(n_351),
.B2(n_346),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_689),
.B(n_352),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_587),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_593),
.B(n_43),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_683),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_571),
.A2(n_358),
.B1(n_359),
.B2(n_356),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_617),
.A2(n_365),
.B1(n_370),
.B2(n_363),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_689),
.B(n_371),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_683),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_692),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_701),
.A2(n_382),
.B1(n_384),
.B2(n_380),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_660),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_584),
.Y(n_753)
);

OA22x2_ASAP7_75t_L g754 ( 
.A1(n_612),
.A2(n_395),
.B1(n_397),
.B2(n_390),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_SL g755 ( 
.A1(n_586),
.A2(n_402),
.B1(n_407),
.B2(n_400),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_701),
.A2(n_413),
.B1(n_415),
.B2(n_411),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_596),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_697),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_562),
.A2(n_424),
.B1(n_425),
.B2(n_417),
.Y(n_760)
);

BUFx10_ASAP7_75t_L g761 ( 
.A(n_560),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_617),
.A2(n_433),
.B1(n_435),
.B2(n_431),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_654),
.B(n_439),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_562),
.A2(n_446),
.B1(n_447),
.B2(n_445),
.Y(n_765)
);

AO22x2_ASAP7_75t_L g766 ( 
.A1(n_563),
.A2(n_566),
.B1(n_655),
.B2(n_640),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_563),
.A2(n_54),
.B1(n_48),
.B2(n_50),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_632),
.A2(n_452),
.B1(n_455),
.B2(n_449),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_SL g770 ( 
.A1(n_632),
.A2(n_558),
.B1(n_556),
.B2(n_554),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_566),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_708),
.A2(n_551),
.B1(n_550),
.B2(n_548),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_456),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_673),
.B(n_460),
.Y(n_774)
);

AO22x2_ASAP7_75t_L g775 ( 
.A1(n_640),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_673),
.B(n_463),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_SL g778 ( 
.A1(n_659),
.A2(n_546),
.B1(n_543),
.B2(n_538),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_687),
.A2(n_496),
.B1(n_527),
.B2(n_524),
.Y(n_779)
);

AND2x2_ASAP7_75t_SL g780 ( 
.A(n_684),
.B(n_56),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_559),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_568),
.A2(n_529),
.B1(n_523),
.B2(n_522),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_713),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_687),
.A2(n_519),
.B1(n_518),
.B2(n_514),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_SL g785 ( 
.A1(n_625),
.A2(n_650),
.B1(n_671),
.B2(n_651),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_568),
.A2(n_510),
.B1(n_507),
.B2(n_506),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_599),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_559),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_599),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_685),
.A2(n_505),
.B1(n_500),
.B2(n_497),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_639),
.A2(n_493),
.B1(n_492),
.B2(n_490),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_627),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_627),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_693),
.A2(n_487),
.B1(n_484),
.B2(n_480),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_702),
.A2(n_470),
.B1(n_477),
.B2(n_475),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_567),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_SL g797 ( 
.A1(n_639),
.A2(n_644),
.B1(n_661),
.B2(n_673),
.Y(n_797)
);

OA22x2_ASAP7_75t_L g798 ( 
.A1(n_670),
.A2(n_478),
.B1(n_474),
.B2(n_469),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_567),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_673),
.B(n_464),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_560),
.B(n_467),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_698),
.B(n_87),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_674),
.B(n_89),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_674),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_644),
.B(n_655),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_635),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_635),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_703),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_703),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_705),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_710),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_SL g812 ( 
.A1(n_602),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_647),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_787),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_783),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_718),
.B(n_704),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_781),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_781),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_788),
.Y(n_819)
);

XOR2xp5_ASAP7_75t_L g820 ( 
.A(n_723),
.B(n_601),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_796),
.Y(n_821)
);

INVxp33_ASAP7_75t_L g822 ( 
.A(n_805),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_720),
.B(n_709),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_799),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_748),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_742),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_761),
.B(n_637),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_748),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_761),
.B(n_762),
.Y(n_830)
);

XOR2xp5_ASAP7_75t_L g831 ( 
.A(n_719),
.B(n_94),
.Y(n_831)
);

XOR2xp5_ASAP7_75t_L g832 ( 
.A(n_728),
.B(n_759),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_753),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_716),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_797),
.B(n_607),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_757),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_789),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_716),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_801),
.B(n_664),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_792),
.B(n_698),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_744),
.B(n_664),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_769),
.Y(n_843)
);

BUFx5_ASAP7_75t_L g844 ( 
.A(n_803),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_746),
.B(n_698),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_758),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_793),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_733),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_806),
.Y(n_849)
);

XOR2xp5_ASAP7_75t_L g850 ( 
.A(n_790),
.B(n_95),
.Y(n_850)
);

XOR2xp5_ASAP7_75t_L g851 ( 
.A(n_794),
.B(n_98),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_807),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_813),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_737),
.B(n_647),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_754),
.A2(n_573),
.B(n_570),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_766),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_766),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_804),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_727),
.B(n_575),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_808),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_717),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_772),
.B(n_724),
.Y(n_863)
);

BUFx8_ASAP7_75t_L g864 ( 
.A(n_731),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_735),
.Y(n_865)
);

XNOR2x2_ASAP7_75t_L g866 ( 
.A(n_752),
.B(n_585),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_750),
.B(n_698),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_717),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_733),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_798),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_R g871 ( 
.A(n_743),
.B(n_690),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_756),
.B(n_707),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_722),
.Y(n_873)
);

NOR2x1_ASAP7_75t_L g874 ( 
.A(n_736),
.B(n_603),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_764),
.B(n_690),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_722),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_621),
.B(n_573),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_773),
.B(n_561),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_749),
.B(n_774),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_730),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_725),
.B(n_710),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_755),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_776),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_767),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_795),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_767),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_785),
.B(n_653),
.Y(n_887)
);

XOR2xp5_ASAP7_75t_L g888 ( 
.A(n_751),
.B(n_102),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_765),
.B(n_707),
.Y(n_889)
);

CKINVDCx16_ASAP7_75t_R g890 ( 
.A(n_800),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_771),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_741),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_771),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_802),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_780),
.B(n_621),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_786),
.B(n_707),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_775),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_809),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_715),
.B(n_616),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_745),
.B(n_707),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_763),
.B(n_564),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_770),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_775),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_778),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_738),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_768),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_854),
.B(n_738),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_857),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_822),
.B(n_823),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_822),
.B(n_752),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_815),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_875),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_856),
.B(n_688),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_833),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_836),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_870),
.B(n_688),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_855),
.B(n_670),
.Y(n_918)
);

AND2x2_ASAP7_75t_SL g919 ( 
.A(n_863),
.B(n_570),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_838),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_830),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_860),
.B(n_747),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_821),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_840),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_875),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_839),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_860),
.B(n_779),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_840),
.B(n_688),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_878),
.A2(n_740),
.B(n_739),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_875),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_846),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_878),
.A2(n_577),
.B(n_565),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_847),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_816),
.B(n_784),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_849),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_894),
.B(n_760),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_892),
.B(n_791),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_875),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_884),
.B(n_810),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_883),
.B(n_688),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_875),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_892),
.B(n_782),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_852),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_843),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_825),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_855),
.B(n_895),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_837),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_844),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_895),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_879),
.B(n_648),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_844),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_826),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_819),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_906),
.B(n_721),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_862),
.B(n_868),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_827),
.Y(n_956)
);

CKINVDCx8_ASAP7_75t_R g957 ( 
.A(n_890),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_814),
.B(n_729),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_853),
.B(n_726),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_835),
.A2(n_714),
.B(n_589),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_824),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_858),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_871),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_814),
.B(n_666),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_873),
.B(n_623),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_829),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_817),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_842),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_842),
.B(n_675),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_818),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_844),
.B(n_732),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_853),
.B(n_680),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_848),
.B(n_711),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_874),
.B(n_615),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_844),
.B(n_579),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_841),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_835),
.B(n_615),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_844),
.B(n_877),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_899),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_904),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_876),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_844),
.B(n_615),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_859),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_861),
.B(n_898),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_881),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_903),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_877),
.B(n_615),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_901),
.B(n_636),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_905),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_867),
.B(n_734),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_841),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_869),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_861),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_898),
.B(n_682),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_828),
.B(n_729),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_886),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_891),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_897),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_893),
.B(n_679),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_889),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_924),
.B(n_845),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_963),
.B(n_865),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_919),
.B(n_887),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_993),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_980),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_SL g1007 ( 
.A(n_930),
.B(n_902),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_987),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_924),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_914),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_909),
.B(n_900),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_924),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_930),
.B(n_882),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_986),
.B(n_885),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_914),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_985),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_909),
.B(n_900),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_L g1018 ( 
.A(n_986),
.B(n_850),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_987),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_964),
.B(n_831),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_922),
.B(n_867),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_924),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_1001),
.B(n_872),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_993),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_930),
.B(n_872),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_919),
.B(n_889),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_937),
.B(n_1001),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_956),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_921),
.B(n_866),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_994),
.B(n_832),
.Y(n_1030)
);

BUFx4f_ASAP7_75t_L g1031 ( 
.A(n_981),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_981),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_985),
.B(n_896),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_964),
.B(n_896),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_997),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_996),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_938),
.B(n_585),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_956),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_960),
.B(n_918),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_L g1040 ( 
.A(n_938),
.B(n_851),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_946),
.Y(n_1041)
);

BUFx8_ASAP7_75t_SL g1042 ( 
.A(n_942),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_965),
.B(n_646),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_965),
.B(n_652),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_915),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_938),
.B(n_567),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_918),
.B(n_811),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_910),
.B(n_820),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_995),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_965),
.B(n_668),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_910),
.B(n_888),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_955),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_957),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_955),
.B(n_694),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_927),
.B(n_583),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_956),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_944),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_947),
.B(n_594),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_946),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_995),
.B(n_714),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_944),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_998),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_911),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_978),
.B(n_999),
.Y(n_1064)
);

AND2x2_ASAP7_75t_SL g1065 ( 
.A(n_973),
.B(n_589),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_926),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_999),
.B(n_591),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_933),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_939),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_917),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_912),
.B(n_812),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_949),
.B(n_605),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_977),
.B(n_591),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_935),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_950),
.B(n_972),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_917),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_950),
.B(n_618),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_962),
.B(n_626),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_972),
.B(n_631),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_1000),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_976),
.B(n_592),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_962),
.B(n_665),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_957),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_907),
.B(n_665),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_1032),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1032),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_1069),
.B(n_938),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1039),
.A2(n_959),
.B1(n_939),
.B2(n_929),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_1024),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1005),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_1032),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_1012),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1006),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_1006),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_1053),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1077),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_1036),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1012),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_1012),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1010),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_1037),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1033),
.B(n_1027),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1008),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_1031),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_1016),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1021),
.B(n_934),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_SL g1108 ( 
.A(n_1078),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1031),
.B(n_941),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1039),
.A2(n_959),
.B1(n_939),
.B2(n_954),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1059),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_1009),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_1036),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1052),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1002),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1015),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1019),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_907),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1054),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1002),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1016),
.B(n_991),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1052),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_1083),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1042),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1035),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_1049),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1014),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_1048),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1051),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1062),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_1009),
.B(n_941),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1022),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_1049),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1022),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1082),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1021),
.B(n_992),
.Y(n_1137)
);

BUFx2_ASAP7_75t_SL g1138 ( 
.A(n_1075),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1054),
.Y(n_1139)
);

INVx8_ASAP7_75t_L g1140 ( 
.A(n_1037),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1043),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1028),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1028),
.Y(n_1143)
);

BUFx2_ASAP7_75t_R g1144 ( 
.A(n_1026),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1038),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1026),
.A2(n_951),
.B1(n_948),
.B2(n_981),
.Y(n_1146)
);

CKINVDCx8_ASAP7_75t_R g1147 ( 
.A(n_1078),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1079),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1066),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1068),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_1072),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1038),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1074),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1043),
.Y(n_1154)
);

BUFx10_ASAP7_75t_L g1155 ( 
.A(n_1058),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1080),
.B(n_1044),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1044),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1050),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1127),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1128),
.A2(n_1030),
.B1(n_1003),
.B2(n_1018),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1111),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1101),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1132),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1127),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1134),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1101),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1089),
.A2(n_1060),
.B1(n_1047),
.B2(n_1034),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1134),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1125),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1149),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1116),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1103),
.A2(n_1071),
.B1(n_1047),
.B2(n_1013),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1118),
.B(n_1011),
.Y(n_1174)
);

INVx8_ASAP7_75t_L g1175 ( 
.A(n_1093),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1116),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1107),
.B(n_1060),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1132),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1150),
.Y(n_1179)
);

CKINVDCx6p67_ASAP7_75t_R g1180 ( 
.A(n_1123),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1153),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1104),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1117),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1088),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1133),
.Y(n_1185)
);

INVx6_ASAP7_75t_L g1186 ( 
.A(n_1093),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1106),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1146),
.A2(n_932),
.B(n_1064),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1138),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1115),
.B(n_955),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1133),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1106),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1093),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1091),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_1096),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1135),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1089),
.A2(n_1004),
.B1(n_1017),
.B2(n_1071),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1110),
.A2(n_1081),
.B1(n_1041),
.B2(n_1064),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_1108),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1156),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1121),
.A2(n_1073),
.B(n_1023),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1093),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1100),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1121),
.A2(n_1081),
.B1(n_1029),
.B2(n_1025),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1156),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1100),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1088),
.A2(n_1025),
.B1(n_1067),
.B2(n_1084),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1108),
.A2(n_1013),
.B1(n_1065),
.B2(n_1007),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1123),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1099),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1136),
.A2(n_1073),
.B1(n_954),
.B2(n_936),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1099),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1100),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1088),
.B(n_1067),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1135),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1099),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1130),
.A2(n_1007),
.B1(n_1040),
.B2(n_1055),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1142),
.B(n_1057),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1099),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1142),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1142),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1141),
.A2(n_939),
.B1(n_1082),
.B2(n_936),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1090),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1094),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1102),
.A2(n_951),
.B(n_948),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1147),
.A2(n_1082),
.B1(n_1151),
.B2(n_971),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1141),
.A2(n_939),
.B1(n_958),
.B2(n_971),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1124),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1087),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1100),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1094),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1229),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1179),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1227),
.A2(n_1155),
.B1(n_1151),
.B2(n_1129),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1170),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1209),
.A2(n_984),
.B1(n_1148),
.B2(n_1097),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1171),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1175),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1174),
.B(n_1119),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1173),
.A2(n_622),
.B1(n_613),
.B2(n_597),
.C(n_638),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1162),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1162),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1177),
.B(n_1126),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1181),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1182),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1161),
.A2(n_871),
.B1(n_1157),
.B2(n_1154),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1183),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1163),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1205),
.A2(n_1095),
.B1(n_1113),
.B2(n_1098),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1195),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1218),
.A2(n_1209),
.B1(n_1189),
.B2(n_1198),
.Y(n_1252)
);

AOI222xp33_ASAP7_75t_L g1253 ( 
.A1(n_1173),
.A2(n_669),
.B1(n_1085),
.B2(n_613),
.C1(n_622),
.C2(n_592),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1189),
.A2(n_1144),
.B1(n_1105),
.B2(n_1131),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1194),
.B(n_1126),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1205),
.A2(n_1157),
.B1(n_1159),
.B2(n_1158),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1212),
.A2(n_1105),
.B1(n_1131),
.B2(n_1158),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1206),
.B(n_1159),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1196),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1175),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1172),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1176),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1168),
.A2(n_1139),
.B1(n_1072),
.B2(n_1113),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1180),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1160),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1165),
.Y(n_1268)
);

NOR2x1_ASAP7_75t_SL g1269 ( 
.A(n_1166),
.B(n_1102),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1168),
.A2(n_1120),
.B1(n_1115),
.B2(n_1037),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1202),
.B(n_1212),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1223),
.A2(n_1120),
.B1(n_1037),
.B2(n_989),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1202),
.B(n_968),
.Y(n_1273)
);

BUFx5_ASAP7_75t_L g1274 ( 
.A(n_1169),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1199),
.A2(n_988),
.B(n_931),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_SL g1276 ( 
.A1(n_1228),
.A2(n_989),
.B(n_969),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1187),
.B(n_969),
.Y(n_1277)
);

INVx4_ASAP7_75t_SL g1278 ( 
.A(n_1186),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1190),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1232),
.B(n_1114),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1199),
.A2(n_1208),
.B(n_1215),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1208),
.A2(n_1215),
.B1(n_1184),
.B2(n_1061),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1184),
.A2(n_1076),
.B1(n_1070),
.B2(n_920),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1210),
.B(n_1114),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1192),
.A2(n_630),
.B1(n_634),
.B2(n_597),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1219),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1200),
.A2(n_920),
.B1(n_953),
.B2(n_961),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1219),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1186),
.A2(n_1109),
.B1(n_1102),
.B2(n_1114),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_SL g1290 ( 
.A(n_1224),
.B(n_864),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1211),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1185),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1175),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1225),
.A2(n_961),
.B1(n_967),
.B2(n_970),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1213),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1191),
.B(n_979),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1197),
.B(n_1122),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1217),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1237),
.A2(n_630),
.B1(n_638),
.B2(n_634),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1258),
.B(n_1221),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1237),
.A2(n_1247),
.B1(n_1252),
.B2(n_1253),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1255),
.B(n_1221),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1285),
.A2(n_1254),
.B1(n_1271),
.B2(n_1281),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1286),
.B(n_1230),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1235),
.A2(n_1109),
.B1(n_1203),
.B2(n_1186),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1267),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1285),
.A2(n_1140),
.B1(n_1207),
.B2(n_1203),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1241),
.A2(n_669),
.B1(n_1140),
.B2(n_967),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1250),
.A2(n_1140),
.B1(n_928),
.B2(n_1216),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1268),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1244),
.B(n_1222),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1265),
.A2(n_679),
.B1(n_695),
.B2(n_700),
.C(n_1000),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1256),
.A2(n_928),
.B1(n_952),
.B2(n_1122),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1272),
.A2(n_928),
.B1(n_1122),
.B2(n_700),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1270),
.A2(n_1122),
.B1(n_695),
.B2(n_1045),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1240),
.A2(n_1273),
.B1(n_1257),
.B2(n_1242),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1274),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1288),
.B(n_1222),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1282),
.A2(n_1164),
.B1(n_1178),
.B2(n_940),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1236),
.B(n_1188),
.Y(n_1320)
);

AOI222xp33_ASAP7_75t_L g1321 ( 
.A1(n_1276),
.A2(n_629),
.B1(n_983),
.B2(n_981),
.C1(n_940),
.C2(n_916),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1279),
.A2(n_940),
.B1(n_923),
.B2(n_956),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1238),
.B(n_1220),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1294),
.B(n_662),
.C(n_649),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1243),
.A2(n_923),
.B1(n_966),
.B2(n_941),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1259),
.A2(n_923),
.B1(n_966),
.B2(n_941),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1287),
.A2(n_966),
.B1(n_916),
.B2(n_1152),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1277),
.A2(n_1275),
.B1(n_1234),
.B2(n_1284),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1290),
.A2(n_1207),
.B1(n_1214),
.B2(n_1231),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1266),
.A2(n_912),
.B1(n_925),
.B2(n_1112),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1274),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1280),
.A2(n_966),
.B1(n_916),
.B2(n_1145),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1297),
.A2(n_1274),
.B1(n_1251),
.B2(n_1246),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1274),
.A2(n_1152),
.B1(n_1142),
.B2(n_1143),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1274),
.A2(n_1152),
.B1(n_1143),
.B2(n_1145),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1233),
.A2(n_1296),
.B1(n_1260),
.B2(n_1245),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1263),
.B(n_1220),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1248),
.A2(n_1292),
.B1(n_1283),
.B2(n_1249),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1291),
.B(n_1143),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1261),
.A2(n_1145),
.B1(n_1152),
.B2(n_1143),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1264),
.A2(n_1145),
.B1(n_945),
.B2(n_913),
.Y(n_1341)
);

AOI222xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1298),
.A2(n_629),
.B1(n_72),
.B2(n_73),
.C1(n_75),
.C2(n_77),
.Y(n_1342)
);

OAI222xp33_ASAP7_75t_L g1343 ( 
.A1(n_1295),
.A2(n_1204),
.B1(n_1193),
.B2(n_1056),
.C1(n_945),
.C2(n_913),
.Y(n_1343)
);

AOI222xp33_ASAP7_75t_L g1344 ( 
.A1(n_1278),
.A2(n_913),
.B1(n_649),
.B2(n_662),
.C1(n_663),
.C2(n_667),
.Y(n_1344)
);

OAI221xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1262),
.A2(n_990),
.B1(n_974),
.B2(n_77),
.C(n_78),
.Y(n_1345)
);

AOI221xp5_ASAP7_75t_L g1346 ( 
.A1(n_1289),
.A2(n_691),
.B1(n_712),
.B2(n_699),
.C(n_681),
.Y(n_1346)
);

OAI222xp33_ASAP7_75t_L g1347 ( 
.A1(n_1262),
.A2(n_1204),
.B1(n_1193),
.B2(n_1056),
.C1(n_945),
.C2(n_990),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1278),
.B(n_982),
.C(n_925),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1269),
.B(n_1087),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1239),
.A2(n_925),
.B1(n_912),
.B2(n_663),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1239),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1239),
.A2(n_662),
.B1(n_672),
.B2(n_678),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1293),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1293),
.A2(n_649),
.B1(n_678),
.B2(n_681),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1252),
.A2(n_1086),
.B1(n_1092),
.B2(n_908),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1252),
.B(n_1092),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1258),
.B(n_1092),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1235),
.A2(n_908),
.B1(n_975),
.B2(n_663),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1237),
.A2(n_672),
.B1(n_691),
.B2(n_699),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1281),
.A2(n_932),
.B(n_1226),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1235),
.A2(n_1086),
.B1(n_908),
.B2(n_1046),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1258),
.B(n_667),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1235),
.A2(n_951),
.B1(n_948),
.B2(n_975),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1323),
.B(n_71),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1306),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1301),
.A2(n_75),
.B1(n_79),
.B2(n_81),
.C(n_82),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_R g1367 ( 
.A(n_1351),
.B(n_103),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1311),
.B(n_82),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1303),
.A2(n_712),
.B1(n_681),
.B2(n_678),
.Y(n_1369)
);

OAI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1299),
.A2(n_672),
.B1(n_667),
.B2(n_624),
.C(n_604),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1302),
.B(n_83),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1306),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1300),
.B(n_569),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1310),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_645),
.B1(n_569),
.B2(n_641),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1304),
.B(n_569),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1345),
.A2(n_645),
.B1(n_576),
.B2(n_641),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1328),
.B(n_645),
.C(n_576),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_576),
.C(n_641),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1304),
.B(n_595),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1318),
.B(n_595),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1318),
.B(n_598),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1356),
.B(n_1362),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1339),
.B(n_107),
.Y(n_1384)
);

OAI221xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1359),
.A2(n_111),
.B1(n_115),
.B2(n_118),
.C(n_123),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1336),
.A2(n_1329),
.B(n_1307),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1339),
.B(n_128),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1358),
.A2(n_1308),
.B(n_1324),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1357),
.B(n_598),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1338),
.B(n_598),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1333),
.B(n_130),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1312),
.B(n_610),
.C(n_633),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1355),
.B(n_610),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1337),
.B(n_619),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1320),
.B(n_619),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1321),
.B(n_643),
.C(n_611),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1361),
.B(n_564),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1320),
.A2(n_131),
.B(n_132),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1351),
.B(n_133),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1353),
.B(n_134),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1309),
.A2(n_643),
.B1(n_611),
.B2(n_606),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1313),
.A2(n_136),
.B(n_137),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1353),
.B(n_138),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1317),
.A2(n_140),
.B(n_141),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1319),
.B(n_643),
.C(n_611),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1317),
.B(n_143),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1344),
.B(n_606),
.C(n_580),
.Y(n_1407)
);

AOI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1305),
.A2(n_146),
.B(n_150),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1331),
.B(n_152),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1331),
.B(n_153),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1349),
.B(n_159),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1315),
.B(n_167),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1314),
.A2(n_170),
.B1(n_172),
.B2(n_175),
.C(n_177),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1395),
.Y(n_1414)
);

NAND4xp75_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1330),
.C(n_1346),
.D(n_1360),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1383),
.B(n_1360),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1372),
.B(n_1360),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1372),
.Y(n_1419)
);

OA211x2_ASAP7_75t_L g1420 ( 
.A1(n_1397),
.A2(n_1369),
.B(n_1393),
.C(n_1378),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1369),
.B(n_1352),
.C(n_1354),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1397),
.A2(n_1347),
.B(n_1343),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1366),
.B(n_1340),
.C(n_1332),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1374),
.B(n_1334),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1371),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1364),
.B(n_1335),
.Y(n_1426)
);

NOR3xp33_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_1408),
.C(n_1385),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1402),
.A2(n_1327),
.B1(n_1322),
.B2(n_1348),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1365),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1368),
.B(n_1326),
.C(n_1325),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1398),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1396),
.A2(n_1341),
.B1(n_1363),
.B2(n_1350),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1398),
.B(n_1404),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1411),
.B(n_580),
.C(n_564),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1379),
.B(n_580),
.C(n_564),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1404),
.B(n_180),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1406),
.A2(n_181),
.B(n_186),
.Y(n_1438)
);

AOI211xp5_ASAP7_75t_L g1439 ( 
.A1(n_1413),
.A2(n_187),
.B(n_188),
.C(n_189),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1380),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1381),
.B(n_198),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1384),
.B(n_206),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1370),
.A2(n_1375),
.B1(n_1407),
.B2(n_1405),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1373),
.B(n_208),
.C(n_211),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1387),
.B(n_212),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1389),
.B(n_214),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1382),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1394),
.B(n_215),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1416),
.B(n_1391),
.Y(n_1449)
);

NAND4xp75_ASAP7_75t_L g1450 ( 
.A(n_1420),
.B(n_1399),
.C(n_1400),
.D(n_1403),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1419),
.B(n_1367),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1417),
.B(n_1434),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1414),
.B(n_1447),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1433),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1409),
.Y(n_1457)
);

INVxp33_ASAP7_75t_SL g1458 ( 
.A(n_1418),
.Y(n_1458)
);

XOR2x2_ASAP7_75t_L g1459 ( 
.A(n_1439),
.B(n_1412),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1447),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1431),
.B(n_1390),
.Y(n_1461)
);

AND4x1_ASAP7_75t_L g1462 ( 
.A(n_1427),
.B(n_1392),
.C(n_1410),
.D(n_1401),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_219),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1425),
.B(n_220),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_221),
.Y(n_1465)
);

XNOR2x1_ASAP7_75t_L g1466 ( 
.A(n_1426),
.B(n_224),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1424),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1422),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1422),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1453),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1453),
.Y(n_1471)
);

XNOR2x1_ASAP7_75t_L g1472 ( 
.A(n_1466),
.B(n_1415),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1460),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1456),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1452),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1452),
.Y(n_1476)
);

XNOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1466),
.B(n_1423),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1454),
.Y(n_1478)
);

XOR2x2_ASAP7_75t_L g1479 ( 
.A(n_1458),
.B(n_1430),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1455),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1454),
.Y(n_1481)
);

XOR2x2_ASAP7_75t_L g1482 ( 
.A(n_1459),
.B(n_1442),
.Y(n_1482)
);

XOR2x1_ASAP7_75t_L g1483 ( 
.A(n_1469),
.B(n_1468),
.Y(n_1483)
);

XOR2x2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1442),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1467),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1469),
.B(n_1435),
.Y(n_1486)
);

XOR2x2_ASAP7_75t_L g1487 ( 
.A(n_1450),
.B(n_1445),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1474),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1485),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1476),
.B(n_1451),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.Y(n_1491)
);

AO22x2_ASAP7_75t_L g1492 ( 
.A1(n_1477),
.A2(n_1461),
.B1(n_1449),
.B2(n_1457),
.Y(n_1492)
);

AOI22x1_ASAP7_75t_L g1493 ( 
.A1(n_1472),
.A2(n_1479),
.B1(n_1475),
.B2(n_1482),
.Y(n_1493)
);

AO22x2_ASAP7_75t_L g1494 ( 
.A1(n_1486),
.A2(n_1461),
.B1(n_1457),
.B2(n_1465),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1480),
.Y(n_1495)
);

OA22x2_ASAP7_75t_L g1496 ( 
.A1(n_1473),
.A2(n_1464),
.B1(n_1463),
.B2(n_1465),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1484),
.A2(n_1487),
.B1(n_1486),
.B2(n_1438),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1478),
.A2(n_1438),
.B1(n_1443),
.B2(n_1421),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1478),
.Y(n_1500)
);

OAI22x1_ASAP7_75t_L g1501 ( 
.A1(n_1481),
.A2(n_1462),
.B1(n_1444),
.B2(n_1441),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1488),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1489),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1500),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1491),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1497),
.Y(n_1506)
);

XOR2x2_ASAP7_75t_L g1507 ( 
.A(n_1498),
.B(n_1443),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1495),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1494),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1494),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1505),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1505),
.Y(n_1512)
);

OA22x2_ASAP7_75t_L g1513 ( 
.A1(n_1509),
.A2(n_1499),
.B1(n_1501),
.B2(n_1493),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1506),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1504),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1508),
.A2(n_1492),
.B1(n_1483),
.B2(n_1490),
.C(n_1428),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1510),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1502),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1511),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1517),
.B(n_1507),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1513),
.A2(n_1492),
.B1(n_1509),
.B2(n_1496),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1516),
.A2(n_1503),
.B1(n_1504),
.B2(n_1428),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1523)
);

OAI22x1_ASAP7_75t_L g1524 ( 
.A1(n_1518),
.A2(n_1436),
.B1(n_1448),
.B2(n_1446),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1515),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1514),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1519),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1525),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1526),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1523),
.Y(n_1530)
);

OA22x2_ASAP7_75t_L g1531 ( 
.A1(n_1521),
.A2(n_1432),
.B1(n_230),
.B2(n_233),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1520),
.A2(n_1522),
.B1(n_1524),
.B2(n_1432),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1527),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1531),
.A2(n_229),
.B1(n_235),
.B2(n_236),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1530),
.A2(n_1532),
.B1(n_1528),
.B2(n_1529),
.Y(n_1535)
);

AO22x2_ASAP7_75t_L g1536 ( 
.A1(n_1533),
.A2(n_241),
.B1(n_243),
.B2(n_245),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1535),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_1534),
.B1(n_248),
.B2(n_250),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1536),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1536),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1538),
.A2(n_246),
.B1(n_252),
.B2(n_253),
.Y(n_1541)
);

OAI22x1_ASAP7_75t_L g1542 ( 
.A1(n_1540),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1539),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1543),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1542),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1541),
.Y(n_1546)
);

AOI22x1_ASAP7_75t_SL g1547 ( 
.A1(n_1544),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1545),
.A2(n_270),
.B1(n_274),
.B2(n_275),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1547),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1548),
.Y(n_1550)
);

AO22x2_ASAP7_75t_L g1551 ( 
.A1(n_1549),
.A2(n_1546),
.B1(n_278),
.B2(n_281),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1550),
.A2(n_276),
.B1(n_282),
.B2(n_284),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1551),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1552),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1553),
.A2(n_289),
.B1(n_294),
.B2(n_296),
.C(n_301),
.Y(n_1555)
);

AOI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1555),
.A2(n_1554),
.B(n_302),
.C(n_303),
.Y(n_1556)
);


endmodule