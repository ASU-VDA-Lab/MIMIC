module fake_netlist_1_636_n_16 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_16);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_9;
wire n_14;
wire n_10;
wire n_15;
wire n_7;
wire n_8;
AOI22xp33_ASAP7_75t_L g7 ( .A1(n_0), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_7) );
AOI22xp5_ASAP7_75t_L g8 ( .A1(n_1), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_3), .B(n_2), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_1), .B(n_0), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
OAI21xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_12), .B(n_7), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_14), .B1(n_12), .B2(n_2), .Y(n_16) );
endmodule