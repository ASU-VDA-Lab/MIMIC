module fake_jpeg_8042_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_18),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_20),
.B(n_16),
.C(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_54),
.B1(n_61),
.B2(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_29),
.B1(n_25),
.B2(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_31),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_79),
.B(n_32),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_19),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_71),
.Y(n_104)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_78),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_75),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_30),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_29),
.B(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_89),
.B1(n_28),
.B2(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_48),
.B(n_37),
.C(n_38),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_88),
.B(n_69),
.C(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_62),
.B1(n_51),
.B2(n_52),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_101),
.B1(n_114),
.B2(n_116),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_95),
.B(n_94),
.C(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_26),
.B(n_24),
.C(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_48),
.B1(n_53),
.B2(n_16),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_71),
.B1(n_68),
.B2(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_94),
.B(n_103),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_84),
.B1(n_71),
.B2(n_67),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_37),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_66),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_131),
.C(n_143),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_126),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_123),
.B1(n_140),
.B2(n_14),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_86),
.B1(n_79),
.B2(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_132),
.B1(n_145),
.B2(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_75),
.B1(n_60),
.B2(n_85),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_133),
.B(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_31),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_83),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_141),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_115),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_108),
.B1(n_100),
.B2(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_0),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_31),
.Y(n_143)
);

AOI22x1_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_106),
.B1(n_92),
.B2(n_91),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_81),
.B1(n_70),
.B2(n_60),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_109),
.B1(n_111),
.B2(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_149),
.B(n_153),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_40),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_168),
.C(n_169),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_171),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_159),
.B(n_173),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_0),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_13),
.B(n_10),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_40),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_60),
.B1(n_56),
.B2(n_93),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_153),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_38),
.B1(n_16),
.B2(n_64),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_123),
.B1(n_136),
.B2(n_128),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_64),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_0),
.C(n_1),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_176),
.C(n_177),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_15),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_13),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_8),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_175),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_121),
.A2(n_120),
.B1(n_133),
.B2(n_129),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_14),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_13),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_0),
.C(n_1),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_2),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_176),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_132),
.B(n_134),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_201),
.B(n_202),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_132),
.B(n_14),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_151),
.B1(n_157),
.B2(n_154),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_178),
.B1(n_166),
.B2(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_2),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_10),
.B(n_9),
.C(n_4),
.D(n_5),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_223),
.B1(n_226),
.B2(n_201),
.Y(n_239)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_198),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_152),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_165),
.C(n_168),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_165),
.C(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_6),
.C(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_6),
.B1(n_9),
.B2(n_185),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_184),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_208),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_182),
.C(n_194),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_186),
.C(n_183),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_225),
.C(n_217),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_180),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_228),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_191),
.B(n_202),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_215),
.B(n_191),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_251),
.C(n_253),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_243),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_191),
.A3(n_195),
.B1(n_215),
.B2(n_216),
.C(n_214),
.Y(n_257)
);

NOR2x1_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_245),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_206),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_231),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_259),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_212),
.B1(n_208),
.B2(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_229),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_270),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_273),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_232),
.B(n_237),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_249),
.B(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_180),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_231),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_209),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_278),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_255),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_271),
.B(n_217),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_248),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_212),
.B1(n_258),
.B2(n_242),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_256),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_267),
.B(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_267),
.C(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_221),
.B(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

OAI21x1_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_251),
.B(n_224),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_296),
.B(n_284),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_282),
.C(n_281),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_298),
.B(n_292),
.Y(n_299)
);

OAI211xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_295),
.B(n_281),
.C(n_219),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_222),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_192),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_9),
.Y(n_303)
);


endmodule