module fake_jpeg_2465_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_70),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_51),
.B1(n_46),
.B2(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_0),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_61),
.B1(n_44),
.B2(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_75),
.B1(n_82),
.B2(n_68),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_61),
.B1(n_56),
.B2(n_49),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_79),
.B(n_67),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_57),
.C(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_54),
.C(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_44),
.B1(n_53),
.B2(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_57),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_69),
.B1(n_63),
.B2(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_92),
.B1(n_100),
.B2(n_81),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_77),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_97),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_2),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_1),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_56),
.B1(n_52),
.B2(n_66),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_108),
.B1(n_112),
.B2(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_52),
.B1(n_60),
.B2(n_46),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_77),
.B(n_4),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_116),
.B(n_96),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_77),
.B1(n_8),
.B2(n_9),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_23),
.B1(n_41),
.B2(n_40),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_8),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_11),
.CON(n_133),
.SN(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_117),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_128),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_10),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_100),
.B1(n_27),
.B2(n_28),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_135),
.B1(n_12),
.B2(n_13),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_11),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_13),
.B(n_14),
.Y(n_150)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_25),
.B1(n_39),
.B2(n_38),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_22),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_43),
.B(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_12),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_150),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_31),
.B(n_32),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_141),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_15),
.B(n_16),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_15),
.B1(n_18),
.B2(n_131),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_125),
.B1(n_135),
.B2(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_125),
.C(n_133),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_146),
.C(n_144),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_152),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.C(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_155),
.Y(n_170)
);

OAI31xp33_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_160),
.A3(n_166),
.B(n_153),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_158),
.B(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_164),
.C(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_149),
.Y(n_179)
);


endmodule