module fake_jpeg_22594_n_310 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_34),
.B1(n_26),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_33),
.B1(n_17),
.B2(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_32),
.B1(n_21),
.B2(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_79),
.B1(n_89),
.B2(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_49),
.B1(n_25),
.B2(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_85),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_39),
.B(n_23),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_91),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_59),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_27),
.B1(n_20),
.B2(n_19),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_17),
.C(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_58),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_45),
.C(n_15),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_47),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_83),
.B(n_80),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_89),
.B(n_84),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_110),
.Y(n_142)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_67),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_52),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_118),
.Y(n_148)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_48),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_90),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_81),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_131),
.B(n_107),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_136),
.C(n_85),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_79),
.B1(n_76),
.B2(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_72),
.B(n_74),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_146),
.B(n_98),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_140),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_84),
.C(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_88),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_94),
.B(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_120),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_78),
.B1(n_46),
.B2(n_63),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_157),
.B(n_159),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_102),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_175),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_103),
.B(n_110),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_96),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_179),
.C(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_171),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_120),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_121),
.B(n_109),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_147),
.B1(n_144),
.B2(n_124),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_0),
.Y(n_181)
);

XNOR2x2_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_112),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_152),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_136),
.B1(n_137),
.B2(n_128),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_185),
.B1(n_187),
.B2(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_197),
.C(n_205),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_129),
.B(n_143),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_140),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_169),
.B(n_138),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_204),
.B(n_157),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_201),
.B1(n_163),
.B2(n_160),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_158),
.B1(n_167),
.B2(n_155),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_156),
.B1(n_168),
.B2(n_173),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_133),
.C(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_171),
.C(n_165),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_178),
.C(n_154),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_153),
.C(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_163),
.B1(n_153),
.B2(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_180),
.C(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_172),
.B1(n_180),
.B2(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_161),
.C(n_172),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_184),
.C(n_187),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_181),
.C(n_169),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_185),
.B1(n_198),
.B2(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_52),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_189),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_231),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_249),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_111),
.B(n_2),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_247),
.B1(n_251),
.B2(n_66),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_203),
.B1(n_204),
.B2(n_198),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_189),
.B1(n_52),
.B2(n_59),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_255),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_228),
.B(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_256),
.B1(n_251),
.B2(n_245),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_211),
.B(n_222),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_212),
.B1(n_217),
.B2(n_225),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_216),
.C(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.C(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_210),
.C(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_111),
.C(n_93),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_237),
.B(n_0),
.CI(n_1),
.CON(n_263),
.SN(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_61),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_248),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_243),
.B1(n_241),
.B2(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_233),
.B1(n_249),
.B2(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_258),
.C(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_246),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_7),
.B(n_16),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_259),
.B(n_261),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_7),
.B(n_16),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_263),
.C(n_11),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_276),
.C(n_278),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_66),
.B1(n_61),
.B2(n_57),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_276),
.B1(n_270),
.B2(n_273),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_292),
.C(n_295),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_9),
.B(n_16),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_293),
.A2(n_286),
.B(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_297),
.B(n_3),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_57),
.C(n_66),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_303),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_279),
.A3(n_282),
.B1(n_281),
.B2(n_287),
.C1(n_5),
.C2(n_6),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_305)
);

A2O1A1O1Ixp25_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_5),
.B(n_12),
.C(n_14),
.D(n_4),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_5),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_2),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_4),
.B1(n_297),
.B2(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_307),
.Y(n_310)
);


endmodule