module fake_jpeg_29935_n_433 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_433);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_49),
.Y(n_149)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_8),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_56),
.Y(n_107)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_10),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_83),
.Y(n_101)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_63),
.Y(n_120)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_10),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_22),
.A2(n_6),
.B1(n_13),
.B2(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_39),
.B1(n_44),
.B2(n_27),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_34),
.B(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_84),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_46),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_11),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_91),
.Y(n_127)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_29),
.C(n_33),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_45),
.B1(n_76),
.B2(n_88),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_32),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_18),
.B1(n_22),
.B2(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_123),
.B1(n_142),
.B2(n_53),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_44),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_126),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_22),
.B1(n_33),
.B2(n_37),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_36),
.B(n_32),
.C(n_27),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_19),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_37),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_37),
.B1(n_45),
.B2(n_38),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_37),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_38),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_150),
.Y(n_208)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_155),
.Y(n_232)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_158),
.A2(n_140),
.B1(n_120),
.B2(n_98),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_159),
.A2(n_170),
.B1(n_175),
.B2(n_184),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_89),
.B1(n_77),
.B2(n_92),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_91),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_168),
.Y(n_204)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_24),
.Y(n_217)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_96),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_67),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_100),
.A2(n_72),
.B1(n_82),
.B2(n_81),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_42),
.CI(n_90),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_80),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_179),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_38),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_185),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_64),
.B1(n_74),
.B2(n_71),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_101),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_75),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_68),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_183),
.Y(n_206)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_95),
.A2(n_24),
.B(n_38),
.C(n_31),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_182),
.B(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_48),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_112),
.A2(n_61),
.B1(n_57),
.B2(n_37),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_47),
.B1(n_14),
.B2(n_2),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_107),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_187),
.Y(n_198)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_122),
.B(n_31),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_31),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_134),
.Y(n_214)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_38),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_24),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_168),
.C(n_171),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_179),
.C(n_174),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_217),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_145),
.B1(n_136),
.B2(n_148),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_123),
.B1(n_150),
.B2(n_143),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_210),
.A2(n_212),
.B1(n_155),
.B2(n_166),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_98),
.B1(n_116),
.B2(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_206),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_120),
.B(n_107),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_141),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_231),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_105),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_154),
.B(n_131),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_184),
.B1(n_174),
.B2(n_195),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_234),
.A2(n_240),
.B1(n_244),
.B2(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_239),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_264),
.C(n_223),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_195),
.B1(n_170),
.B2(n_159),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_188),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_206),
.B(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_252),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_136),
.B1(n_145),
.B2(n_178),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_245),
.A2(n_265),
.B(n_223),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_182),
.B1(n_161),
.B2(n_152),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_185),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_211),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_204),
.B(n_157),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_251),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_156),
.C(n_176),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_205),
.A2(n_146),
.B1(n_114),
.B2(n_115),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_146),
.B1(n_114),
.B2(n_143),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_117),
.B1(n_208),
.B2(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_261),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_194),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_225),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_205),
.A2(n_117),
.B1(n_148),
.B2(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_181),
.C(n_151),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_106),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_198),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_245),
.B(n_227),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_270),
.A2(n_281),
.B(n_220),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_202),
.C(n_228),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_271),
.B(n_272),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_237),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_279),
.C(n_286),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_214),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_247),
.A2(n_226),
.B(n_211),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_285),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_198),
.C(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_249),
.B(n_230),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_258),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_250),
.B1(n_261),
.B2(n_252),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_218),
.C(n_197),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_197),
.C(n_221),
.Y(n_292)
);

XOR2x2_ASAP7_75t_SL g293 ( 
.A(n_246),
.B(n_216),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_294),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_254),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_236),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_311),
.Y(n_335)
);

OAI22x1_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_260),
.B1(n_240),
.B2(n_234),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_303),
.B1(n_309),
.B2(n_312),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_301),
.B(n_313),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_272),
.C(n_238),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_305),
.B(n_270),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_266),
.B1(n_235),
.B2(n_247),
.Y(n_306)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_235),
.B1(n_264),
.B2(n_248),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_277),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_283),
.A2(n_255),
.B1(n_256),
.B2(n_262),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_263),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_243),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_317),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_321),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_269),
.A2(n_243),
.B1(n_253),
.B2(n_225),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_290),
.B1(n_285),
.B2(n_284),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_320),
.A2(n_275),
.B(n_289),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_221),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_196),
.B1(n_200),
.B2(n_220),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_323),
.A2(n_275),
.B1(n_200),
.B2(n_295),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_296),
.C(n_271),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_331),
.C(n_334),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_271),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_339),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_330),
.A2(n_347),
.B1(n_312),
.B2(n_323),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_279),
.C(n_286),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_291),
.C(n_292),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_320),
.B(n_300),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_341),
.B(n_315),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_282),
.C(n_268),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_342),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_340),
.B1(n_190),
.B2(n_108),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_277),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_309),
.A2(n_269),
.B1(n_268),
.B2(n_287),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_287),
.C(n_289),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_284),
.C(n_196),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_229),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_208),
.B1(n_193),
.B2(n_219),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_324),
.B(n_308),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_329),
.C(n_339),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_349),
.A2(n_367),
.B(n_119),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_346),
.A2(n_308),
.B1(n_303),
.B2(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_328),
.A2(n_307),
.B1(n_318),
.B2(n_316),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_351),
.A2(n_352),
.B1(n_337),
.B2(n_333),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_358),
.Y(n_376)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_359),
.Y(n_372)
);

A2O1A1O1Ixp25_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_313),
.B(n_321),
.C(n_302),
.D(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_0),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_361),
.B(n_362),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_363),
.A2(n_338),
.B1(n_341),
.B2(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_364),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_368),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_330),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_366),
.B(n_325),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_229),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_187),
.C(n_173),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_384),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_343),
.C(n_342),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_378),
.C(n_381),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_374),
.A2(n_380),
.B1(n_367),
.B2(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_331),
.C(n_334),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_327),
.C(n_164),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_108),
.C(n_119),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_368),
.C(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_382),
.B(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_389),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_379),
.A2(n_352),
.B1(n_364),
.B2(n_349),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_387),
.A2(n_392),
.B1(n_13),
.B2(n_14),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_382),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_373),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_355),
.B1(n_361),
.B2(n_348),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_395),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_371),
.B(n_359),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_360),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_381),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_378),
.C(n_370),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_380),
.B(n_384),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_403),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_373),
.B(n_376),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_385),
.C(n_403),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_407),
.C(n_23),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_385),
.A2(n_376),
.B(n_358),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_404),
.B(n_399),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_31),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_5),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_413),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_402),
.A2(n_391),
.B1(n_392),
.B2(n_388),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g411 ( 
.A1(n_398),
.A2(n_13),
.B(n_14),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_411),
.B(n_12),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_416),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_401),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_23),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_412),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_420),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_421),
.B(n_0),
.Y(n_425)
);

A2O1A1O1Ixp25_ASAP7_75t_L g428 ( 
.A1(n_425),
.A2(n_426),
.B(n_427),
.C(n_411),
.D(n_423),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_400),
.C(n_417),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_405),
.C(n_415),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_429),
.C(n_0),
.Y(n_430)
);

AOI321xp33_ASAP7_75t_L g429 ( 
.A1(n_424),
.A2(n_407),
.A3(n_12),
.B1(n_13),
.B2(n_23),
.C(n_31),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_1),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_1),
.B(n_23),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_1),
.B1(n_382),
.B2(n_308),
.Y(n_433)
);


endmodule