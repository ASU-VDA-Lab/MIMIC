module fake_jpeg_28768_n_408 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_79),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_27),
.B(n_2),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_72),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_73),
.B(n_75),
.Y(n_142)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_77),
.B(n_81),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_2),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_41),
.B1(n_34),
.B2(n_22),
.Y(n_105)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_14),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_12),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_80),
.Y(n_140)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_17),
.B(n_12),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_37),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_33),
.B1(n_40),
.B2(n_43),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_118),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_21),
.B1(n_43),
.B2(n_17),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_47),
.B1(n_77),
.B2(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_26),
.B1(n_34),
.B2(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_68),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_122),
.B1(n_67),
.B2(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_46),
.A2(n_28),
.B1(n_11),
.B2(n_10),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_116),
.B1(n_129),
.B2(n_132),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_50),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_94),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_65),
.B1(n_64),
.B2(n_78),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_8),
.B1(n_9),
.B2(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_114),
.B1(n_119),
.B2(n_96),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_69),
.A2(n_61),
.B1(n_56),
.B2(n_57),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_8),
.B1(n_80),
.B2(n_81),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_58),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_60),
.A2(n_81),
.B1(n_48),
.B2(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_48),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_146),
.A2(n_151),
.B1(n_164),
.B2(n_93),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_98),
.B(n_55),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_148),
.B(n_188),
.Y(n_204)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_162),
.Y(n_196)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_156),
.Y(n_190)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_119),
.Y(n_157)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_58),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_159),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_54),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_98),
.B(n_66),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_179),
.Y(n_202)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_110),
.A2(n_140),
.B(n_108),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_183),
.B(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_92),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_113),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_102),
.B1(n_128),
.B2(n_165),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_111),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_137),
.B1(n_118),
.B2(n_139),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_180),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_104),
.B(n_124),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_106),
.B(n_101),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_144),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_134),
.B1(n_141),
.B2(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_141),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_224),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_123),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_216),
.B(n_153),
.C(n_151),
.D(n_164),
.Y(n_244)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_159),
.B(n_138),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_127),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_221),
.Y(n_230)
);

AOI22x1_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_127),
.B1(n_93),
.B2(n_143),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_179),
.B(n_121),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_171),
.B(n_121),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_154),
.A2(n_128),
.B1(n_145),
.B2(n_164),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_155),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_226),
.B(n_231),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_220),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_220),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_154),
.B1(n_175),
.B2(n_183),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_237),
.B1(n_240),
.B2(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_152),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_246),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_162),
.B1(n_177),
.B2(n_166),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_216),
.B1(n_192),
.B2(n_221),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_248),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_148),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_256),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_244),
.A2(n_189),
.B(n_190),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_180),
.B1(n_167),
.B2(n_145),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_225),
.B1(n_211),
.B2(n_214),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_152),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_206),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_197),
.A2(n_180),
.B1(n_167),
.B2(n_145),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_156),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_207),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_161),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_157),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_205),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_208),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_211),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_281),
.C(n_239),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_283),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_192),
.B(n_200),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_228),
.B(n_238),
.Y(n_303)
);

AOI221xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_198),
.B1(n_219),
.B2(n_199),
.C(n_210),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_237),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_189),
.B(n_205),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_280),
.B(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_199),
.B1(n_185),
.B2(n_190),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_282),
.B1(n_284),
.B2(n_257),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_252),
.Y(n_292)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_193),
.A3(n_217),
.B1(n_209),
.B2(n_150),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_228),
.Y(n_297)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_189),
.B(n_193),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_203),
.C(n_209),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_217),
.B1(n_184),
.B2(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_229),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_242),
.A2(n_203),
.B1(n_157),
.B2(n_212),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_227),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_295),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_297),
.B1(n_261),
.B2(n_267),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_293),
.B(n_248),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_298),
.B1(n_282),
.B2(n_262),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_246),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_236),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_254),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_307),
.C(n_258),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_239),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_301),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_306),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_305),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_266),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_231),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_278),
.A2(n_253),
.A3(n_255),
.B1(n_243),
.B2(n_244),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_258),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_270),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_268),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_261),
.B1(n_278),
.B2(n_285),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_312),
.A2(n_301),
.B1(n_298),
.B2(n_294),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_313),
.B(n_324),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_277),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_317),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_281),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_276),
.C(n_272),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_330),
.C(n_331),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_309),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_321),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_331),
.B(n_330),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_326),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_272),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_278),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_271),
.C(n_280),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_289),
.C(n_303),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_318),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_312),
.A2(n_301),
.B1(n_316),
.B2(n_313),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_340),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_344),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_349),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_308),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_284),
.B(n_310),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_348),
.A2(n_338),
.B(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_320),
.A2(n_310),
.B(n_315),
.Y(n_350)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_288),
.B(n_249),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_327),
.B1(n_328),
.B2(n_290),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_351),
.A2(n_288),
.B1(n_234),
.B2(n_279),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_329),
.C(n_327),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_355),
.C(n_360),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_287),
.C(n_283),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_345),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_302),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_344),
.B(n_251),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_362),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_335),
.B1(n_349),
.B2(n_351),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_334),
.C(n_347),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_346),
.B(n_287),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_365),
.Y(n_369)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_370),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_361),
.A2(n_348),
.B1(n_337),
.B2(n_333),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_373),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_352),
.A2(n_334),
.B1(n_343),
.B2(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_366),
.Y(n_385)
);

OAI211xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_234),
.B(n_319),
.C(n_208),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_376),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_354),
.A2(n_319),
.B(n_273),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_273),
.C(n_247),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_372),
.C(n_363),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

NOR2x1p5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_365),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_386),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_386),
.C(n_383),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_360),
.C(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_388),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_223),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_381),
.A2(n_373),
.B(n_378),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_389),
.A2(n_395),
.B(n_383),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_393),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_371),
.C(n_369),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_380),
.A2(n_376),
.B(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_384),
.A2(n_176),
.B(n_212),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_392),
.Y(n_402)
);

AOI311xp33_ASAP7_75t_SL g399 ( 
.A1(n_393),
.A2(n_208),
.A3(n_213),
.B(n_223),
.C(n_201),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_213),
.A3(n_201),
.B1(n_163),
.B2(n_187),
.C1(n_149),
.C2(n_169),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_213),
.B(n_223),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_201),
.A3(n_163),
.B1(n_391),
.B2(n_176),
.C1(n_182),
.C2(n_170),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_401),
.B(n_397),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_404),
.C(n_150),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_406),
.B(n_178),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_178),
.Y(n_408)
);


endmodule