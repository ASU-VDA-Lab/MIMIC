module fake_netlist_6_4020_n_904 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_904);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_904;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_683;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_811;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_817;
wire n_701;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_SL g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_89),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_54),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_104),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_125),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_22),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_60),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_80),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_121),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_65),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_186),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_128),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_91),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_120),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_130),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_188),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_10),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_189),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_199),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_17),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_18),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_82),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_145),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_117),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_51),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_44),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_138),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_99),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_72),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_170),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_144),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_166),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_50),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_2),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

INVxp33_ASAP7_75t_SL g285 ( 
.A(n_216),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_203),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_205),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_213),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_224),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_209),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_211),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_207),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_207),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_206),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_206),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_260),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_210),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_226),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_R g326 ( 
.A(n_229),
.B(n_28),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_230),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_202),
.B1(n_212),
.B2(n_273),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_314),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_277),
.B(n_214),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_265),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_201),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_325),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_282),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_280),
.B(n_315),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

AND3x1_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_263),
.C(n_247),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_214),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_277),
.B(n_214),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_315),
.B(n_247),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_324),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_291),
.B(n_293),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_286),
.B(n_267),
.Y(n_363)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_263),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_244),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_319),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_319),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_287),
.A2(n_269),
.B(n_257),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_269),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_288),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_285),
.A2(n_261),
.B1(n_262),
.B2(n_266),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_244),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_294),
.B(n_244),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_298),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_R g385 ( 
.A(n_342),
.B(n_299),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_342),
.B(n_296),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g390 ( 
.A1(n_330),
.A2(n_316),
.B1(n_287),
.B2(n_303),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_368),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_249),
.Y(n_392)
);

AND3x2_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_381),
.C(n_374),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_337),
.B(n_259),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

OAI221xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_357),
.B1(n_343),
.B2(n_340),
.C(n_339),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_383),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_337),
.B(n_350),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_379),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_299),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_303),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_316),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_371),
.A2(n_275),
.B1(n_272),
.B2(n_268),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_350),
.B(n_270),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_231),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_370),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_380),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_276),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_362),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_367),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_234),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_235),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_367),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_383),
.B(n_237),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_318),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_364),
.B(n_238),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_344),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_369),
.B(n_322),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_376),
.B(n_29),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_334),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_367),
.B(n_240),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_242),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_339),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_242),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_347),
.A2(n_262),
.B1(n_266),
.B2(n_271),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_383),
.B(n_243),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_380),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_338),
.B(n_248),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_338),
.B(n_251),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_341),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g453 ( 
.A1(n_373),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_358),
.B(n_252),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_373),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_420),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_369),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_369),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_403),
.A2(n_369),
.B1(n_382),
.B2(n_336),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_385),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_385),
.Y(n_466)
);

AO22x2_ASAP7_75t_L g467 ( 
.A1(n_415),
.A2(n_403),
.B1(n_453),
.B2(n_391),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_397),
.B(n_358),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

OAI221xp5_ASAP7_75t_L g473 ( 
.A1(n_400),
.A2(n_341),
.B1(n_343),
.B2(n_375),
.C(n_366),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

OR2x2_ASAP7_75t_SL g475 ( 
.A(n_410),
.B(n_289),
.Y(n_475)
);

AO22x2_ASAP7_75t_L g476 ( 
.A1(n_415),
.A2(n_453),
.B1(n_413),
.B2(n_355),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_418),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_384),
.B(n_380),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_345),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

OAI221xp5_ASAP7_75t_L g482 ( 
.A1(n_451),
.A2(n_405),
.B1(n_411),
.B2(n_408),
.C(n_449),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_431),
.A2(n_412),
.B1(n_418),
.B2(n_444),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_453),
.A2(n_338),
.B1(n_365),
.B2(n_366),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_423),
.A2(n_365),
.B(n_348),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_429),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_392),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_392),
.B(n_358),
.Y(n_494)
);

BUFx8_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g497 ( 
.A1(n_440),
.A2(n_365),
.B1(n_6),
.B2(n_7),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_392),
.A2(n_365),
.B1(n_274),
.B2(n_345),
.Y(n_498)
);

AO22x2_ASAP7_75t_L g499 ( 
.A1(n_417),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_499)
);

NOR4xp25_ASAP7_75t_SL g500 ( 
.A(n_423),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_395),
.A2(n_345),
.B1(n_346),
.B2(n_358),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

AO22x2_ASAP7_75t_L g503 ( 
.A1(n_432),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

AO22x2_ASAP7_75t_L g506 ( 
.A1(n_432),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_429),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_422),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_452),
.A2(n_346),
.B1(n_359),
.B2(n_361),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_359),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_414),
.A2(n_346),
.B1(n_352),
.B2(n_349),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_433),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_429),
.Y(n_513)
);

AO22x2_ASAP7_75t_L g514 ( 
.A1(n_422),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_427),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_427),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_419),
.B(n_359),
.Y(n_519)
);

AOI22x1_ASAP7_75t_L g520 ( 
.A1(n_450),
.A2(n_447),
.B1(n_446),
.B2(n_426),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_393),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_450),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_452),
.A2(n_361),
.B1(n_359),
.B2(n_352),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

AO22x2_ASAP7_75t_L g527 ( 
.A1(n_443),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_464),
.B(n_443),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_457),
.B(n_401),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_461),
.B(n_401),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_468),
.B(n_419),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_456),
.B(n_419),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_493),
.B(n_390),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_455),
.B(n_419),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_SL g535 ( 
.A(n_466),
.B(n_446),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_493),
.B(n_390),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g537 ( 
.A(n_477),
.B(n_447),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_458),
.B(n_419),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_458),
.B(n_414),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_486),
.B(n_416),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_459),
.B(n_430),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_507),
.B(n_454),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_460),
.B(n_441),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_502),
.B(n_437),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_434),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_513),
.B(n_393),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_479),
.B(n_421),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_480),
.B(n_495),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_495),
.B(n_434),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_485),
.B(n_492),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_510),
.B(n_421),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_463),
.B(n_434),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_465),
.B(n_470),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_500),
.B(n_421),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_474),
.B(n_421),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_484),
.B(n_434),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_487),
.B(n_335),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_498),
.B(n_335),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_494),
.B(n_348),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_501),
.B(n_434),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_496),
.B(n_359),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_520),
.B(n_349),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_520),
.B(n_361),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_524),
.B(n_361),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_521),
.B(n_497),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_509),
.B(n_361),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_496),
.B(n_23),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_483),
.B(n_31),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_483),
.B(n_32),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_481),
.B(n_33),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_490),
.B(n_34),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_24),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_504),
.B(n_36),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_505),
.B(n_37),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_491),
.B(n_25),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_512),
.B(n_38),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_516),
.B(n_518),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_522),
.B(n_25),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_519),
.B(n_26),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_511),
.B(n_40),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_41),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_482),
.B(n_42),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_526),
.B(n_43),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_523),
.B(n_46),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_525),
.B(n_47),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_469),
.B(n_48),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_471),
.B(n_472),
.Y(n_587)
);

O2A1O1Ixp5_ASAP7_75t_SL g588 ( 
.A1(n_562),
.A2(n_527),
.B(n_517),
.C(n_515),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_548),
.B(n_478),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_539),
.A2(n_473),
.B(n_467),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_584),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_584),
.Y(n_592)
);

AO31x2_ASAP7_75t_L g593 ( 
.A1(n_532),
.A2(n_467),
.A3(n_476),
.B(n_488),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_582),
.A2(n_503),
.B1(n_506),
.B2(n_475),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_541),
.B(n_476),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_538),
.A2(n_488),
.B(n_497),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

AOI31xp67_ASAP7_75t_L g598 ( 
.A1(n_563),
.A2(n_527),
.A3(n_517),
.B(n_515),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_533),
.B(n_26),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_539),
.A2(n_534),
.B1(n_530),
.B2(n_560),
.Y(n_601)
);

AO31x2_ASAP7_75t_L g602 ( 
.A1(n_531),
.A2(n_506),
.A3(n_503),
.B(n_514),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_540),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_R g604 ( 
.A(n_560),
.B(n_49),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_536),
.A2(n_514),
.B(n_508),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

O2A1O1Ixp5_ASAP7_75t_L g607 ( 
.A1(n_529),
.A2(n_508),
.B(n_499),
.C(n_55),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_116),
.B(n_52),
.Y(n_608)
);

AOI221xp5_ASAP7_75t_SL g609 ( 
.A1(n_572),
.A2(n_499),
.B1(n_27),
.B2(n_57),
.C(n_58),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_551),
.A2(n_118),
.B(n_56),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_553),
.B(n_27),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_545),
.A2(n_59),
.B(n_61),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_581),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_550),
.B(n_586),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_543),
.B(n_62),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_578),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

OAI22x1_ASAP7_75t_L g620 ( 
.A1(n_580),
.A2(n_558),
.B1(n_586),
.B2(n_555),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_556),
.A2(n_63),
.B(n_66),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_575),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_549),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_67),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_564),
.A2(n_68),
.B(n_69),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_568),
.B(n_70),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_566),
.A2(n_71),
.B(n_74),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_554),
.A2(n_75),
.B(n_76),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_569),
.A2(n_77),
.B(n_78),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_573),
.A2(n_79),
.B(n_81),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_528),
.B(n_542),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_579),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_585),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_537),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_615),
.B(n_574),
.Y(n_636)
);

OA21x2_ASAP7_75t_L g637 ( 
.A1(n_590),
.A2(n_576),
.B(n_571),
.Y(n_637)
);

OAI21x1_ASAP7_75t_SL g638 ( 
.A1(n_629),
.A2(n_547),
.B(n_570),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_620),
.A2(n_535),
.B(n_546),
.Y(n_639)
);

BUFx2_ASAP7_75t_SL g640 ( 
.A(n_624),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_609),
.A2(n_83),
.B(n_85),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_618),
.B(n_86),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_600),
.B(n_87),
.C(n_88),
.Y(n_643)
);

OAI21x1_ASAP7_75t_SL g644 ( 
.A1(n_617),
.A2(n_90),
.B(n_92),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_618),
.B(n_93),
.Y(n_645)
);

AO221x2_ASAP7_75t_L g646 ( 
.A1(n_594),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_646)
);

NAND2x1p5_ASAP7_75t_L g647 ( 
.A(n_624),
.B(n_100),
.Y(n_647)
);

AOI21xp33_ASAP7_75t_L g648 ( 
.A1(n_603),
.A2(n_101),
.B(n_102),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_626),
.A2(n_105),
.B(n_106),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_624),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_605),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_628),
.A2(n_110),
.B(n_111),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_606),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_616),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_599),
.Y(n_656)
);

OAI21x1_ASAP7_75t_SL g657 ( 
.A1(n_595),
.A2(n_115),
.B(n_119),
.Y(n_657)
);

CKINVDCx11_ASAP7_75t_R g658 ( 
.A(n_597),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_610),
.A2(n_122),
.B(n_123),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_630),
.A2(n_124),
.B(n_126),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_605),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.C(n_132),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_604),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_592),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_614),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_592),
.B(n_139),
.Y(n_665)
);

OAI21xp33_ASAP7_75t_L g666 ( 
.A1(n_611),
.A2(n_140),
.B(n_141),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_632),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_147),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_619),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_613),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_608),
.A2(n_148),
.B(n_151),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_631),
.A2(n_152),
.B(n_153),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_635),
.Y(n_674)
);

AOI21xp33_ASAP7_75t_L g675 ( 
.A1(n_601),
.A2(n_633),
.B(n_623),
.Y(n_675)
);

AOI221xp5_ASAP7_75t_SL g676 ( 
.A1(n_635),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.C(n_159),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_613),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_596),
.A2(n_160),
.B(n_161),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_612),
.A2(n_163),
.B(n_167),
.Y(n_679)
);

OAI21x1_ASAP7_75t_SL g680 ( 
.A1(n_622),
.A2(n_171),
.B(n_172),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_650),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_641),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_641),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_655),
.Y(n_685)
);

AO21x2_ASAP7_75t_L g686 ( 
.A1(n_638),
.A2(n_627),
.B(n_634),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_669),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_664),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_656),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_674),
.B(n_589),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_678),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_659),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_646),
.B(n_602),
.Y(n_693)
);

AO31x2_ASAP7_75t_L g694 ( 
.A1(n_652),
.A2(n_598),
.A3(n_588),
.B(n_609),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_651),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_651),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_678),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_646),
.B(n_602),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_646),
.A2(n_625),
.B1(n_592),
.B2(n_627),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_672),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_675),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_660),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_639),
.A2(n_607),
.B(n_625),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_673),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_680),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_637),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_637),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_637),
.B(n_593),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_636),
.B(n_602),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_679),
.A2(n_593),
.B(n_174),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_677),
.Y(n_713)
);

OA21x2_ASAP7_75t_L g714 ( 
.A1(n_676),
.A2(n_593),
.B(n_176),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_657),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_642),
.B(n_173),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_644),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_662),
.A2(n_178),
.B1(n_180),
.B2(n_183),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_652),
.B(n_184),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_665),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_670),
.B(n_198),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_665),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_658),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_665),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_663),
.B(n_185),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_643),
.A2(n_193),
.B(n_194),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_647),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_647),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_SL g730 ( 
.A(n_700),
.B(n_651),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_702),
.B(n_642),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_711),
.B(n_645),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_R g733 ( 
.A(n_723),
.B(n_663),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_720),
.B(n_671),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_720),
.B(n_671),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_722),
.B(n_677),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_722),
.B(n_668),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_R g738 ( 
.A(n_719),
.B(n_640),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_690),
.B(n_658),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_R g740 ( 
.A(n_719),
.B(n_196),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_713),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_726),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_713),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_685),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_R g745 ( 
.A(n_721),
.B(n_662),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_724),
.B(n_667),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_685),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_711),
.B(n_667),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_697),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_713),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_724),
.B(n_654),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_724),
.B(n_654),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_697),
.B(n_661),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_688),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_R g755 ( 
.A(n_721),
.B(n_648),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_726),
.B(n_666),
.Y(n_756)
);

XOR2xp5_ASAP7_75t_L g757 ( 
.A(n_716),
.B(n_725),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_702),
.B(n_689),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_R g759 ( 
.A(n_697),
.B(n_695),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_697),
.B(n_695),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_688),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_728),
.B(n_729),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_697),
.B(n_729),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_728),
.B(n_697),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_R g765 ( 
.A(n_725),
.B(n_715),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_687),
.B(n_689),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_687),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_687),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_689),
.Y(n_769)
);

CKINVDCx12_ASAP7_75t_R g770 ( 
.A(n_707),
.Y(n_770)
);

INVx5_ASAP7_75t_SL g771 ( 
.A(n_751),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_732),
.B(n_693),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_731),
.B(n_699),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_766),
.B(n_693),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_766),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_768),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_758),
.B(n_708),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_747),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_769),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_762),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_757),
.B(n_699),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_754),
.B(n_708),
.Y(n_783)
);

NOR2x1_ASAP7_75t_SL g784 ( 
.A(n_761),
.B(n_686),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_767),
.B(n_709),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_742),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_762),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_748),
.B(n_710),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_764),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_737),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_765),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_764),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_743),
.B(n_709),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_737),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_749),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_734),
.B(n_709),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_734),
.B(n_709),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_746),
.B(n_710),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_746),
.B(n_710),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_751),
.B(n_698),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_752),
.B(n_698),
.Y(n_801)
);

NAND5xp2_ASAP7_75t_L g802 ( 
.A(n_782),
.B(n_704),
.C(n_727),
.D(n_739),
.E(n_715),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_781),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_778),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_794),
.B(n_750),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_776),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_794),
.B(n_736),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_778),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_791),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_794),
.B(n_736),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_786),
.B(n_752),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_779),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_773),
.B(n_741),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_790),
.A2(n_740),
.B1(n_738),
.B2(n_730),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_787),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_795),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_787),
.B(n_735),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_784),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_783),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_774),
.B(n_735),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_781),
.B(n_753),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_819),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_806),
.B(n_774),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_819),
.B(n_788),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_804),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_816),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_815),
.B(n_811),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_808),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_805),
.B(n_775),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_809),
.B(n_788),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_809),
.B(n_798),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_812),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_827),
.B(n_814),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_823),
.A2(n_821),
.B1(n_745),
.B2(n_755),
.Y(n_834)
);

AO221x2_ASAP7_75t_L g835 ( 
.A1(n_825),
.A2(n_813),
.B1(n_802),
.B2(n_821),
.C(n_792),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_830),
.B(n_763),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_827),
.B(n_816),
.Y(n_837)
);

AO221x2_ASAP7_75t_L g838 ( 
.A1(n_832),
.A2(n_789),
.B1(n_792),
.B2(n_779),
.C(n_775),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_838),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_833),
.B(n_822),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_837),
.B(n_824),
.Y(n_841)
);

CKINVDCx16_ASAP7_75t_R g842 ( 
.A(n_834),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_835),
.B(n_829),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_L g844 ( 
.A1(n_839),
.A2(n_818),
.B(n_823),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_842),
.A2(n_836),
.B1(n_840),
.B2(n_843),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_840),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_841),
.A2(n_826),
.B1(n_807),
.B2(n_803),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_839),
.A2(n_817),
.B(n_831),
.C(n_830),
.Y(n_848)
);

NOR2x1_ASAP7_75t_L g849 ( 
.A(n_846),
.B(n_831),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_845),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_849),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_850),
.B(n_848),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_849),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_852),
.B(n_844),
.C(n_847),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_851),
.A2(n_817),
.B(n_828),
.C(n_824),
.Y(n_855)
);

NAND4xp25_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_733),
.C(n_717),
.D(n_810),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_L g857 ( 
.A(n_852),
.B(n_718),
.C(n_717),
.Y(n_857)
);

NOR4xp25_ASAP7_75t_L g858 ( 
.A(n_852),
.B(n_828),
.C(n_795),
.D(n_789),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_852),
.B(n_707),
.C(n_712),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

OA211x2_ASAP7_75t_L g861 ( 
.A1(n_857),
.A2(n_770),
.B(n_759),
.C(n_760),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_858),
.B(n_820),
.Y(n_862)
);

AOI222xp33_ASAP7_75t_L g863 ( 
.A1(n_855),
.A2(n_784),
.B1(n_810),
.B2(n_756),
.C1(n_772),
.C2(n_771),
.Y(n_863)
);

OAI211xp5_ASAP7_75t_SL g864 ( 
.A1(n_854),
.A2(n_793),
.B(n_682),
.C(n_681),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_859),
.B(n_810),
.Y(n_865)
);

OAI211xp5_ASAP7_75t_L g866 ( 
.A1(n_860),
.A2(n_714),
.B(n_793),
.C(n_712),
.Y(n_866)
);

XNOR2x1_ASAP7_75t_L g867 ( 
.A(n_861),
.B(n_756),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_864),
.B(n_797),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_SL g869 ( 
.A(n_865),
.B(n_714),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_862),
.B(n_681),
.C(n_682),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_863),
.B(n_780),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_868),
.B(n_772),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_R g873 ( 
.A(n_867),
.B(n_801),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_870),
.B(n_714),
.C(n_777),
.Y(n_874)
);

XNOR2xp5_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_686),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_866),
.B(n_869),
.C(n_714),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_870),
.B(n_800),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_R g878 ( 
.A(n_868),
.B(n_801),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_870),
.B(n_800),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_870),
.B(n_797),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_SL g881 ( 
.A(n_870),
.B(n_777),
.C(n_705),
.Y(n_881)
);

XOR2xp5_ASAP7_75t_L g882 ( 
.A(n_875),
.B(n_797),
.Y(n_882)
);

OAI221xp5_ASAP7_75t_L g883 ( 
.A1(n_876),
.A2(n_705),
.B1(n_703),
.B2(n_701),
.C(n_692),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_880),
.A2(n_686),
.B1(n_797),
.B2(n_796),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_877),
.A2(n_796),
.B1(n_798),
.B2(n_799),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_873),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_879),
.Y(n_887)
);

OAI221xp5_ASAP7_75t_L g888 ( 
.A1(n_874),
.A2(n_703),
.B1(n_701),
.B2(n_692),
.C(n_706),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_881),
.B(n_771),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_872),
.A2(n_691),
.B1(n_796),
.B2(n_780),
.C(n_799),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_886),
.A2(n_878),
.B1(n_796),
.B2(n_771),
.Y(n_891)
);

OR5x1_ASAP7_75t_L g892 ( 
.A(n_887),
.B(n_771),
.C(n_694),
.D(n_691),
.E(n_696),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_889),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_882),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_884),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_890),
.A2(n_780),
.B(n_691),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_894),
.A2(n_883),
.B1(n_888),
.B2(n_885),
.C(n_701),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_891),
.A2(n_771),
.B1(n_783),
.B2(n_785),
.Y(n_898)
);

AOI31xp33_ASAP7_75t_L g899 ( 
.A1(n_897),
.A2(n_895),
.A3(n_893),
.B(n_892),
.Y(n_899)
);

OR3x1_ASAP7_75t_L g900 ( 
.A(n_899),
.B(n_898),
.C(n_896),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_SL g901 ( 
.A1(n_900),
.A2(n_696),
.B1(n_706),
.B2(n_785),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_901),
.Y(n_902)
);

OAI221xp5_ASAP7_75t_L g903 ( 
.A1(n_902),
.A2(n_706),
.B1(n_696),
.B2(n_684),
.C(n_683),
.Y(n_903)
);

AOI211xp5_ASAP7_75t_L g904 ( 
.A1(n_903),
.A2(n_696),
.B(n_683),
.C(n_684),
.Y(n_904)
);


endmodule