module fake_jpeg_15922_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_15),
.B1(n_36),
.B2(n_23),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_24),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_23),
.B1(n_15),
.B2(n_17),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_25),
.B1(n_28),
.B2(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_35),
.B(n_37),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_19),
.C(n_26),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_66),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_37),
.B1(n_35),
.B2(n_18),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_73),
.B1(n_53),
.B2(n_41),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_34),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_34),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_78),
.Y(n_86)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_58),
.B1(n_53),
.B2(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_68),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_87),
.B(n_98),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_92),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_90),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_30),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_53),
.B1(n_41),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_74),
.B1(n_60),
.B2(n_89),
.Y(n_106)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_34),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_59),
.B1(n_73),
.B2(n_61),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_68),
.B1(n_59),
.B2(n_35),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_79),
.B1(n_93),
.B2(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_34),
.C(n_39),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_34),
.C(n_38),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_32),
.B1(n_43),
.B2(n_56),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_126),
.C(n_131),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_121),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_83),
.B(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_114),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_32),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_26),
.CON(n_127),
.SN(n_127)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_26),
.B(n_77),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_32),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_100),
.B(n_111),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_109),
.C(n_117),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_81),
.B1(n_95),
.B2(n_43),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_81),
.B1(n_38),
.B2(n_30),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_39),
.C(n_50),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_141),
.C(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_140),
.B(n_143),
.Y(n_159)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_121),
.B(n_122),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_126),
.Y(n_141)
);

INVxp33_ASAP7_75t_SL g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_146),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_21),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_1),
.B(n_2),
.Y(n_158)
);

OAI322xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_127),
.A3(n_128),
.B1(n_118),
.B2(n_119),
.C1(n_21),
.C2(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_151),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_128),
.A3(n_21),
.B1(n_10),
.B2(n_12),
.C1(n_9),
.C2(n_13),
.Y(n_151)
);

OA21x2_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_13),
.B(n_12),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_158),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.C(n_147),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_38),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_142),
.B1(n_137),
.B2(n_135),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_156),
.A2(n_139),
.B1(n_136),
.B2(n_11),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_156),
.B1(n_159),
.B2(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_159),
.B(n_162),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_169),
.B(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_183),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_176),
.B(n_3),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_2),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_187),
.C(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_4),
.C(n_5),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_11),
.Y(n_190)
);


endmodule