module fake_jpeg_21916_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_28),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_35),
.B1(n_40),
.B2(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_29),
.B1(n_16),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_62),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_24),
.B2(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_56),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_23),
.B1(n_25),
.B2(n_31),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_19),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_57),
.B1(n_28),
.B2(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_86),
.B1(n_87),
.B2(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_72),
.B1(n_54),
.B2(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_25),
.B1(n_28),
.B2(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_35),
.C(n_39),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_43),
.C(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_31),
.B(n_26),
.C(n_32),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_80),
.C(n_81),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_12),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_12),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_22),
.B1(n_33),
.B2(n_19),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_43),
.A2(n_22),
.B1(n_33),
.B2(n_17),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_70),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_105),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_99),
.C(n_81),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_102),
.B1(n_107),
.B2(n_78),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_14),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_58),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_68),
.B1(n_67),
.B2(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_63),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_66),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_96),
.C(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_26),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_67),
.B1(n_85),
.B2(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_93),
.B1(n_89),
.B2(n_111),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_78),
.B1(n_80),
.B2(n_53),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_129),
.B(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_140),
.B1(n_91),
.B2(n_109),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_84),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_61),
.B1(n_66),
.B2(n_73),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_59),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_167),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_165),
.C(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_155),
.B1(n_138),
.B2(n_143),
.Y(n_180)
);

XNOR2x2_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_98),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_154),
.B(n_159),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_99),
.B(n_110),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_91),
.B1(n_99),
.B2(n_97),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_166),
.B1(n_172),
.B2(n_140),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_93),
.A3(n_112),
.B1(n_114),
.B2(n_17),
.C1(n_27),
.C2(n_26),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_160),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_27),
.B(n_26),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_126),
.B(n_122),
.C(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_133),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_32),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_114),
.B1(n_32),
.B2(n_92),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_7),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_3),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_1),
.C(n_2),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_1),
.C(n_3),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_136),
.C(n_11),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_137),
.B1(n_130),
.B2(n_127),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_160),
.B1(n_169),
.B2(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_150),
.B1(n_167),
.B2(n_144),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_122),
.B(n_126),
.C(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_186),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_119),
.B1(n_117),
.B2(n_121),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_171),
.B(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_194),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_132),
.B1(n_141),
.B2(n_136),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_193),
.B1(n_172),
.B2(n_153),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_168),
.C(n_162),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_141),
.B1(n_133),
.B2(n_6),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_171),
.B1(n_153),
.B2(n_154),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_165),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_193),
.B(n_187),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_175),
.C(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_183),
.C(n_182),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_162),
.B1(n_141),
.B2(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_9),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_186),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_179),
.B(n_192),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_224),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_197),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_217),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_195),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_184),
.C(n_178),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_231),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_230),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_207),
.B(n_218),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_191),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_5),
.C(n_7),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_233),
.A2(n_201),
.B1(n_223),
.B2(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_240),
.B1(n_213),
.B2(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_211),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_202),
.B(n_204),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_239),
.Y(n_254)
);

OAI21x1_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_219),
.B(n_202),
.Y(n_246)
);

AOI21x1_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_249),
.B(n_198),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_208),
.B(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_220),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_254),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_198),
.B1(n_211),
.B2(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_241),
.B1(n_247),
.B2(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_220),
.C(n_221),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_256),
.C(n_259),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_258),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_237),
.B(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_8),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_247),
.B1(n_210),
.B2(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_259),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_258),
.B(n_251),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_262),
.C(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_8),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_269),
.A3(n_261),
.B1(n_264),
.B2(n_263),
.C1(n_250),
.C2(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_8),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_269),
.B(n_253),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_278),
.A3(n_279),
.B1(n_273),
.B2(n_270),
.C1(n_14),
.C2(n_15),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_280),
.Y(n_282)
);

AOI221xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_10),
.B1(n_12),
.B2(n_281),
.C(n_279),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_283),
.Y(n_284)
);


endmodule