module fake_jpeg_3448_n_533 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_533);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_63),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_0),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_62),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_0),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_81),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_22),
.B(n_2),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_28),
.C(n_32),
.Y(n_159)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_17),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_86),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_87),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_93),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_3),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_107),
.Y(n_134)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_29),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_110),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_36),
.B(n_4),
.C(n_5),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_37),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_36),
.B(n_4),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_112),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

CKINVDCx11_ASAP7_75t_R g171 ( 
.A(n_113),
.Y(n_171)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_38),
.B(n_5),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_118),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_21),
.B1(n_46),
.B2(n_43),
.Y(n_156)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_121),
.Y(n_184)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_57),
.B1(n_56),
.B2(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_139),
.A2(n_146),
.B1(n_156),
.B2(n_158),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_63),
.B(n_32),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_144),
.B(n_147),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_56),
.B1(n_45),
.B2(n_40),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_43),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_28),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_153),
.B(n_182),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_70),
.A2(n_71),
.B1(n_122),
.B2(n_82),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_137),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_77),
.A2(n_49),
.B(n_46),
.C(n_33),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_161),
.A2(n_137),
.B(n_155),
.C(n_171),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_69),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_162),
.B(n_167),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_67),
.A2(n_49),
.B1(n_33),
.B2(n_42),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_164),
.A2(n_179),
.B1(n_191),
.B2(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_94),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_108),
.A2(n_42),
.B1(n_35),
.B2(n_26),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_172),
.A2(n_178),
.B1(n_194),
.B2(n_191),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_174),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_87),
.B(n_5),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_6),
.B(n_7),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_100),
.B(n_51),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_73),
.A2(n_83),
.B1(n_90),
.B2(n_99),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_70),
.A2(n_42),
.B1(n_54),
.B2(n_26),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_89),
.B(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_62),
.B(n_8),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_186),
.A2(n_198),
.B(n_131),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_102),
.A2(n_42),
.B1(n_26),
.B2(n_51),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_74),
.B(n_9),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_195),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_113),
.A2(n_26),
.B1(n_51),
.B2(n_54),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_71),
.B(n_9),
.Y(n_195)
);

CKINVDCx11_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_104),
.B(n_14),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_85),
.B(n_14),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_86),
.B(n_15),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_97),
.B1(n_103),
.B2(n_119),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_207),
.B(n_221),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_104),
.B(n_16),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_209),
.A2(n_247),
.B(n_189),
.C(n_231),
.Y(n_281)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_210),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_211),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_212),
.B(n_224),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_214),
.A2(n_240),
.B1(n_206),
.B2(n_232),
.Y(n_305)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_215),
.Y(n_317)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_217),
.Y(n_322)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_218),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_185),
.A2(n_15),
.B1(n_132),
.B2(n_125),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_125),
.A2(n_145),
.B1(n_170),
.B2(n_142),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_220),
.A2(n_260),
.B1(n_270),
.B2(n_210),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_166),
.A2(n_134),
.B1(n_152),
.B2(n_129),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_149),
.A2(n_150),
.B1(n_178),
.B2(n_155),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_234),
.Y(n_295)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_223),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_225),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_221),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_156),
.A2(n_179),
.B1(n_130),
.B2(n_160),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_244),
.B1(n_255),
.B2(n_207),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_124),
.A2(n_141),
.B1(n_180),
.B2(n_168),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_140),
.Y(n_235)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_127),
.B(n_157),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_242),
.Y(n_287)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_146),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_243),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_139),
.B(n_143),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_261),
.Y(n_319)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_246),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_136),
.A2(n_158),
.B(n_190),
.C(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_148),
.Y(n_248)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_249),
.B(n_262),
.Y(n_285)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_256),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_130),
.A2(n_160),
.B1(n_192),
.B2(n_183),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_165),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_263),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_142),
.A2(n_131),
.B1(n_188),
.B2(n_133),
.Y(n_260)
);

AO22x1_ASAP7_75t_SL g261 ( 
.A1(n_183),
.A2(n_200),
.B1(n_192),
.B2(n_126),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_200),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_154),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_265),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_267),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_154),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_269),
.Y(n_294)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_126),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_276),
.A2(n_308),
.B1(n_256),
.B2(n_211),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_163),
.B1(n_133),
.B2(n_189),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_293),
.B1(n_320),
.B2(n_254),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_133),
.B1(n_189),
.B2(n_135),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_279),
.A2(n_305),
.B1(n_277),
.B2(n_320),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_282),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_310),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_229),
.A2(n_238),
.B1(n_205),
.B2(n_244),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_206),
.C(n_240),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_306),
.C(n_309),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_230),
.C(n_227),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_250),
.A2(n_232),
.B1(n_233),
.B2(n_209),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_264),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_222),
.A2(n_237),
.B1(n_209),
.B2(n_234),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_237),
.C(n_216),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_252),
.C(n_248),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_218),
.A2(n_236),
.B1(n_217),
.B2(n_247),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_315),
.A2(n_283),
.B1(n_321),
.B2(n_290),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_261),
.B1(n_223),
.B2(n_203),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_293),
.A2(n_261),
.B1(n_215),
.B2(n_235),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_346),
.B1(n_353),
.B2(n_354),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_300),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_333),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_213),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_326),
.B(n_329),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_328),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_272),
.B(n_253),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_311),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_339),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_332),
.A2(n_291),
.B1(n_322),
.B2(n_313),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_266),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_290),
.A2(n_241),
.B1(n_268),
.B2(n_270),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_340),
.B(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_269),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_208),
.B(n_251),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_226),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_343),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_342),
.A2(n_344),
.B1(n_284),
.B2(n_316),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_246),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_276),
.A2(n_319),
.B1(n_307),
.B2(n_289),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_295),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_356),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_325),
.B1(n_328),
.B2(n_346),
.Y(n_390)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

INVx2_ASAP7_75t_R g351 ( 
.A(n_281),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_351),
.B(n_301),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_319),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_295),
.A2(n_305),
.B1(n_275),
.B2(n_273),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_283),
.A2(n_286),
.B1(n_310),
.B2(n_304),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_298),
.A2(n_304),
.B1(n_292),
.B2(n_299),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_355),
.A2(n_359),
.B1(n_361),
.B2(n_345),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_302),
.B(n_303),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_303),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_358),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_271),
.B(n_280),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_298),
.A2(n_317),
.B1(n_296),
.B2(n_316),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_297),
.A2(n_294),
.B(n_314),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_360),
.A2(n_288),
.B(n_318),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_296),
.A2(n_312),
.B1(n_291),
.B2(n_314),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_312),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_297),
.C(n_278),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_370),
.C(n_384),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_357),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_368),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_288),
.C(n_313),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_323),
.B1(n_355),
.B2(n_327),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_329),
.B(n_322),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_374),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_373),
.A2(n_379),
.B(n_367),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_322),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_318),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_382),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_356),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_333),
.B(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_395),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_390),
.A2(n_328),
.B1(n_332),
.B2(n_337),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_380),
.B1(n_374),
.B2(n_389),
.Y(n_419)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_347),
.C(n_354),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_353),
.C(n_362),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_325),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_401),
.B1(n_411),
.B2(n_422),
.Y(n_433)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_335),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_404),
.C(n_420),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_387),
.A2(n_337),
.B1(n_351),
.B2(n_341),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_417),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_340),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_385),
.Y(n_426)
);

FAx1_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_351),
.CI(n_336),
.CON(n_406),
.SN(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_409),
.B(n_371),
.C(n_391),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_360),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_381),
.Y(n_438)
);

XNOR2x2_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_361),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_359),
.B1(n_342),
.B2(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_367),
.A2(n_342),
.B(n_331),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_413),
.A2(n_415),
.B(n_373),
.Y(n_424)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_372),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_419),
.A2(n_386),
.B1(n_388),
.B2(n_392),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_369),
.C(n_365),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_387),
.A2(n_380),
.B1(n_381),
.B2(n_369),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_424),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_393),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_425),
.B(n_428),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_431),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_393),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_399),
.B(n_385),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_423),
.B(n_363),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_437),
.Y(n_454)
);

BUFx12f_ASAP7_75t_SL g435 ( 
.A(n_406),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_SL g467 ( 
.A(n_435),
.B(n_438),
.C(n_427),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_415),
.A2(n_381),
.B(n_379),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_436),
.B(n_413),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_363),
.C(n_375),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_405),
.C(n_408),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_375),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_443),
.Y(n_453)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_377),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_417),
.B(n_377),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_448),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_445),
.A2(n_444),
.B1(n_397),
.B2(n_437),
.Y(n_450)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_451),
.B(n_460),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_401),
.B1(n_396),
.B2(n_406),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_452),
.A2(n_456),
.B1(n_427),
.B2(n_441),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_402),
.B1(n_414),
.B2(n_407),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_433),
.A2(n_406),
.B1(n_421),
.B2(n_398),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_458),
.A2(n_461),
.B1(n_465),
.B2(n_445),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_383),
.Y(n_459)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_383),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_409),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_469),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_433),
.A2(n_421),
.B1(n_398),
.B2(n_409),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_426),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_410),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_465),
.B1(n_458),
.B2(n_466),
.Y(n_493)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_467),
.B1(n_430),
.B2(n_447),
.Y(n_498)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_455),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_483),
.B1(n_485),
.B2(n_468),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_463),
.A2(n_435),
.B(n_436),
.C(n_424),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_478),
.B(n_462),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_432),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_440),
.C(n_431),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_451),
.Y(n_489)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_455),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_411),
.B(n_446),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_484),
.A2(n_452),
.B(n_463),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_448),
.Y(n_485)
);

NOR3xp33_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_466),
.C(n_457),
.Y(n_486)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_457),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_490),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_489),
.B(n_496),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_493),
.A2(n_475),
.B1(n_472),
.B2(n_476),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_477),
.B(n_483),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_484),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_468),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_485),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_472),
.B1(n_430),
.B2(n_446),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_481),
.C(n_453),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_507),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_508),
.B(n_504),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_480),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_493),
.C(n_480),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_479),
.C(n_482),
.Y(n_507)
);

AOI31xp67_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_486),
.A3(n_495),
.B(n_492),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_470),
.C(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_516),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_501),
.A2(n_488),
.B(n_497),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_502),
.B(n_449),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_517),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_507),
.B(n_386),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_499),
.C(n_505),
.Y(n_519)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_519),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_521),
.A2(n_510),
.B(n_518),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_506),
.C(n_508),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_524),
.B(n_517),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_523),
.A2(n_520),
.B1(n_522),
.B2(n_519),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_525),
.B(n_526),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_528),
.A2(n_449),
.B(n_410),
.C(n_412),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_525),
.A3(n_527),
.B1(n_416),
.B2(n_364),
.C1(n_442),
.C2(n_418),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_442),
.C(n_364),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_532),
.B(n_530),
.Y(n_533)
);


endmodule