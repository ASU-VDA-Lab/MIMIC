module fake_jpeg_19529_n_319 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_11),
.B1(n_12),
.B2(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_26),
.B1(n_11),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_52),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_33),
.C(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_23),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_31),
.C(n_16),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_26),
.B1(n_11),
.B2(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_11),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_26),
.B1(n_11),
.B2(n_13),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_59)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_35),
.B1(n_43),
.B2(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_45),
.B1(n_35),
.B2(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_79),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_46),
.B1(n_53),
.B2(n_60),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_61),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_35),
.B1(n_37),
.B2(n_45),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_47),
.B1(n_56),
.B2(n_55),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_60),
.B1(n_46),
.B2(n_49),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_17),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_88),
.B1(n_95),
.B2(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_73),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_61),
.B(n_52),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_73),
.B(n_70),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_59),
.B1(n_52),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_68),
.B1(n_76),
.B2(n_70),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_97),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_52),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_75),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_110),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_62),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_75),
.C(n_65),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_111),
.C(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_114),
.B1(n_116),
.B2(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_118),
.B(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_108),
.B1(n_115),
.B2(n_113),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_74),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_73),
.C(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_70),
.B1(n_77),
.B2(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_95),
.B1(n_98),
.B2(n_89),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_70),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_94),
.B1(n_62),
.B2(n_40),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_132),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_130),
.B1(n_141),
.B2(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_135),
.B(n_109),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_90),
.B1(n_82),
.B2(n_70),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_118),
.B(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_85),
.C(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_149),
.C(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_40),
.B1(n_28),
.B2(n_25),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_82),
.B1(n_97),
.B2(n_66),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_148),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_82),
.C(n_32),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_129),
.B1(n_136),
.B2(n_133),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_17),
.B(n_22),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_117),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_16),
.B1(n_14),
.B2(n_22),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_20),
.B1(n_19),
.B2(n_13),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_177),
.C(n_149),
.Y(n_197)
);

AND3x1_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_142),
.C(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_104),
.B1(n_102),
.B2(n_0),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_174),
.B1(n_142),
.B2(n_131),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_171),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_172),
.B1(n_180),
.B2(n_182),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_14),
.B1(n_22),
.B2(n_16),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_0),
.B1(n_14),
.B2(n_2),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_176),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_32),
.C(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_154),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_19),
.B1(n_20),
.B2(n_94),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_117),
.B1(n_18),
.B2(n_62),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_185),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_18),
.B1(n_62),
.B2(n_28),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_30),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_171),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_128),
.B(n_141),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_208),
.B1(n_174),
.B2(n_165),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_181),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_192),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_195),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_187),
.B(n_161),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_203),
.C(n_207),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_153),
.C(n_152),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_180),
.B(n_166),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_144),
.C(n_31),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_50),
.C(n_25),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_0),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_25),
.B1(n_50),
.B2(n_31),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_169),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_223),
.B1(n_232),
.B2(n_205),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_189),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_165),
.B1(n_184),
.B2(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_177),
.B1(n_166),
.B2(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_30),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_50),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_50),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_207),
.B(n_18),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_205),
.C(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_229),
.B1(n_231),
.B2(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_202),
.B1(n_209),
.B2(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_247),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_225),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_199),
.B1(n_190),
.B2(n_50),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_50),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_217),
.C(n_220),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_245),
.C(n_239),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_221),
.B(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_217),
.B(n_222),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_242),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_215),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_263),
.B1(n_34),
.B2(n_5),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_264),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_252),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_256),
.B(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_260),
.B1(n_266),
.B2(n_270),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_262),
.B1(n_268),
.B2(n_7),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_279),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_255),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_284),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_18),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_258),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_34),
.C(n_5),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_4),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_290),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_301)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_297),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_6),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_6),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_34),
.B(n_7),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_6),
.B(n_7),
.Y(n_298)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_299),
.A3(n_306),
.B1(n_285),
.B2(n_288),
.C(n_287),
.Y(n_308)
);

HAxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_283),
.CON(n_299),
.SN(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_8),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_296),
.C(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_8),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_309),
.B(n_299),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_293),
.B(n_285),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_310),
.C(n_311),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_9),
.B(n_10),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.C(n_10),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_9),
.Y(n_319)
);


endmodule