module real_jpeg_23393_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_34),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_20),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_27),
.B1(n_46),
.B2(n_66),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_30),
.B1(n_54),
.B2(n_55),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_6),
.B(n_20),
.C(n_23),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_38),
.C(n_40),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_52),
.C(n_55),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_44),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_6),
.B(n_120),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_74),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_70),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_70),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_60),
.C(n_62),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_15),
.A2(n_16),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_31),
.C(n_47),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_17),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_17),
.A2(n_83),
.B1(n_99),
.B2(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_17),
.B(n_116),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_17),
.A2(n_83),
.B1(n_115),
.B2(n_116),
.Y(n_138)
);

AOI211xp5_ASAP7_75t_L g160 ( 
.A1(n_17),
.A2(n_129),
.B(n_132),
.C(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_17),
.A2(n_83),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_17),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_17),
.A2(n_83),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_17),
.A2(n_97),
.B(n_100),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_19),
.A2(n_25),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_19),
.A2(n_25),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_19),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_20),
.A2(n_24),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_20),
.B(n_192),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_31),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_32)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_36),
.A2(n_37),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_40),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_47),
.A2(n_48),
.B1(n_86),
.B2(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_83),
.C(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_57),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_55),
.B(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_61),
.B(n_88),
.Y(n_116)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_90),
.B(n_269),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_76),
.B(n_79),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_85),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_115),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_85),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI31xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_250),
.A3(n_261),
.B(n_266),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_151),
.B(n_249),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_134),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_93),
.B(n_134),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_123),
.B1(n_124),
.B2(n_133),
.Y(n_93)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_113),
.B2(n_114),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_96),
.B(n_113),
.C(n_123),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_111),
.B2(n_112),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_100),
.B1(n_107),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_104),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_127),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_117),
.B(n_122),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_117),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_159),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_116),
.B1(n_129),
.B2(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_115),
.A2(n_116),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_164),
.C(n_179),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_116),
.A2(n_129),
.B(n_161),
.C(n_224),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_122),
.A2(n_255),
.B1(n_259),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_130),
.B(n_131),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_126),
.A2(n_129),
.B1(n_159),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_145),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_129),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_129),
.A2(n_159),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_129),
.A2(n_159),
.B1(n_201),
.B2(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_129),
.A2(n_159),
.B1(n_189),
.B2(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_130),
.A2(n_131),
.B(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_143),
.B(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.C(n_142),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_138),
.B1(n_163),
.B2(n_170),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_144),
.Y(n_238)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_142),
.B(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_243),
.B(n_248),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_182),
.B(n_234),
.C(n_242),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_172),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_154),
.B(n_172),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_162),
.B2(n_171),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_157),
.B(n_160),
.C(n_171),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_186),
.C(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_165),
.C(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_165),
.B1(n_179),
.B2(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_165),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_164),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_164),
.A2(n_165),
.B1(n_190),
.B2(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_165),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_165),
.B(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_174),
.A2(n_175),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_233),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_196),
.B(n_232),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_185),
.B(n_193),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_226),
.B(n_231),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_220),
.B(n_225),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_209),
.B(n_219),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_204),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_236),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_263),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_265),
.Y(n_267)
);


endmodule