module real_aes_835_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g241 ( .A(n_0), .B(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_1), .A2(n_71), .B1(n_385), .B2(n_409), .Y(n_593) );
AO22x2_ASAP7_75t_L g258 ( .A1(n_2), .A2(n_165), .B1(n_248), .B2(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g629 ( .A(n_2), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_3), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_4), .A2(n_13), .B1(n_341), .B2(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_5), .A2(n_61), .B1(n_508), .B2(n_614), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_6), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_7), .A2(n_151), .B1(n_343), .B2(n_481), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_8), .A2(n_52), .B1(n_460), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_9), .A2(n_103), .B1(n_387), .B2(n_388), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_10), .A2(n_199), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_11), .A2(n_121), .B1(n_299), .B2(n_503), .Y(n_502) );
AOI22x1_ASAP7_75t_L g411 ( .A1(n_12), .A2(n_96), .B1(n_387), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_14), .A2(n_192), .B1(n_377), .B2(n_378), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_15), .A2(n_92), .B1(n_489), .B2(n_490), .Y(n_488) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_16), .A2(n_47), .B1(n_248), .B2(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_16), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_17), .A2(n_139), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_18), .A2(n_204), .B1(n_380), .B2(n_381), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_19), .A2(n_160), .B1(n_319), .B2(n_481), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_20), .A2(n_223), .B(n_231), .C(n_631), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_21), .B(n_577), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g389 ( .A(n_22), .B(n_390), .Y(n_389) );
XNOR2xp5_ASAP7_75t_L g415 ( .A(n_22), .B(n_390), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_23), .A2(n_182), .B1(n_299), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_24), .A2(n_25), .B1(n_387), .B2(n_388), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g513 ( .A1(n_26), .A2(n_141), .B1(n_191), .B2(n_275), .C1(n_329), .C2(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_27), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_28), .A2(n_177), .B1(n_284), .B2(n_334), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_29), .A2(n_206), .B1(n_370), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_30), .A2(n_82), .B1(n_385), .B2(n_409), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_31), .B(n_242), .Y(n_474) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_32), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_32), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_33), .A2(n_112), .B1(n_221), .B2(n_261), .C1(n_329), .C2(n_477), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_34), .A2(n_155), .B1(n_369), .B2(n_370), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_35), .A2(n_98), .B1(n_280), .B2(n_284), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_36), .A2(n_62), .B1(n_307), .B2(n_310), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_37), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_38), .A2(n_215), .B1(n_334), .B2(n_470), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_39), .A2(n_216), .B1(n_537), .B2(n_539), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_40), .A2(n_209), .B1(n_275), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_41), .A2(n_175), .B1(n_399), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_42), .A2(n_123), .B1(n_503), .B2(n_587), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_43), .A2(n_633), .B1(n_644), .B2(n_645), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_43), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_44), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_45), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_46), .A2(n_145), .B1(n_319), .B2(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_48), .A2(n_76), .B1(n_372), .B2(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_49), .A2(n_107), .B1(n_291), .B2(n_354), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_50), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_51), .A2(n_110), .B1(n_349), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_53), .A2(n_211), .B1(n_271), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_54), .A2(n_189), .B1(n_377), .B2(n_378), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_55), .A2(n_113), .B1(n_349), .B2(n_454), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_56), .A2(n_97), .B1(n_372), .B2(n_373), .Y(n_424) );
INVx3_ASAP7_75t_L g248 ( .A(n_57), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_58), .A2(n_138), .B1(n_261), .B2(n_337), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_59), .A2(n_166), .B1(n_352), .B2(n_354), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_60), .A2(n_161), .B1(n_486), .B2(n_487), .Y(n_485) );
XOR2x2_ASAP7_75t_L g238 ( .A(n_63), .B(n_239), .Y(n_238) );
AO222x2_ASAP7_75t_L g363 ( .A1(n_64), .A2(n_119), .B1(n_144), .B2(n_364), .C1(n_365), .C2(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g516 ( .A(n_65), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_66), .A2(n_153), .B1(n_378), .B2(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_67), .A2(n_125), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_68), .A2(n_205), .B1(n_271), .B2(n_457), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_69), .A2(n_101), .B1(n_261), .B2(n_512), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_70), .Y(n_547) );
INVx1_ASAP7_75t_SL g249 ( .A(n_72), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_72), .B(n_105), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_73), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_74), .Y(n_395) );
INVx2_ASAP7_75t_L g230 ( .A(n_75), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_77), .A2(n_147), .B1(n_314), .B2(n_318), .Y(n_313) );
OA22x2_ASAP7_75t_L g442 ( .A1(n_78), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_78), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_79), .A2(n_124), .B1(n_346), .B2(n_354), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_80), .A2(n_188), .B1(n_294), .B2(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_81), .A2(n_200), .B1(n_384), .B2(n_385), .Y(n_383) );
OA22x2_ASAP7_75t_L g463 ( .A1(n_83), .A2(n_464), .B1(n_492), .B2(n_493), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_83), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_84), .A2(n_91), .B1(n_280), .B2(n_470), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_85), .A2(n_217), .B1(n_349), .B2(n_350), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_86), .A2(n_134), .B1(n_280), .B2(n_470), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_87), .A2(n_162), .B1(n_486), .B2(n_508), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_88), .A2(n_120), .B1(n_531), .B2(n_533), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_89), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_90), .A2(n_164), .B1(n_452), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_93), .A2(n_181), .B1(n_412), .B2(n_614), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_94), .A2(n_116), .B1(n_280), .B2(n_335), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_95), .A2(n_195), .B1(n_305), .B2(n_489), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_99), .A2(n_115), .B1(n_291), .B2(n_294), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_100), .A2(n_190), .B1(n_588), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_102), .A2(n_201), .B1(n_337), .B2(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_104), .A2(n_196), .B1(n_280), .B2(n_335), .Y(n_461) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_105), .A2(n_172), .B1(n_248), .B2(n_252), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_106), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_108), .A2(n_186), .B1(n_508), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_109), .A2(n_130), .B1(n_334), .B2(n_335), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_111), .A2(n_198), .B1(n_299), .B2(n_302), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_114), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_117), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_118), .A2(n_137), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_122), .A2(n_133), .B1(n_343), .B2(n_452), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_126), .A2(n_179), .B1(n_261), .B2(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g250 ( .A(n_127), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_128), .A2(n_185), .B1(n_365), .B2(n_366), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_129), .A2(n_158), .B1(n_294), .B2(n_299), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_131), .B(n_329), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_132), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_135), .A2(n_148), .B1(n_380), .B2(n_381), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_136), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_140), .A2(n_174), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_142), .A2(n_170), .B1(n_452), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_143), .A2(n_176), .B1(n_261), .B2(n_266), .Y(n_260) );
INVx1_ASAP7_75t_L g597 ( .A(n_146), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_149), .A2(n_167), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_150), .A2(n_159), .B1(n_448), .B2(n_449), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_152), .A2(n_208), .B1(n_299), .B2(n_304), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_154), .A2(n_210), .B1(n_261), .B2(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_156), .A2(n_169), .B1(n_271), .B2(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_157), .B(n_579), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_163), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_168), .A2(n_180), .B1(n_380), .B2(n_388), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_171), .A2(n_218), .B1(n_304), .B2(n_592), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_173), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_178), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g625 ( .A(n_178), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_183), .A2(n_214), .B1(n_512), .B2(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
AND2x2_ASAP7_75t_R g647 ( .A(n_184), .B(n_625), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_187), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_193), .A2(n_220), .B1(n_271), .B2(n_275), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_194), .A2(n_212), .B1(n_271), .B2(n_275), .Y(n_331) );
INVxp67_ASAP7_75t_L g228 ( .A(n_197), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_202), .A2(n_219), .B1(n_385), .B2(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_203), .B(n_364), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_207), .B(n_275), .Y(n_665) );
XNOR2x1_ASAP7_75t_L g324 ( .A(n_213), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_SL g223 ( .A(n_224), .B(n_227), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g673 ( .A(n_225), .B(n_227), .Y(n_673) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_226), .B(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_518), .B1(n_620), .B2(n_621), .C(n_622), .Y(n_231) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_232), .Y(n_620) );
OAI22xp5_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_234), .B1(n_439), .B2(n_517), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B1(n_356), .B2(n_438), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_321), .B1(n_322), .B2(n_355), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g355 ( .A(n_238), .Y(n_355) );
NOR2xp67_ASAP7_75t_L g239 ( .A(n_240), .B(n_289), .Y(n_239) );
NAND4xp25_ASAP7_75t_SL g240 ( .A(n_241), .B(n_260), .C(n_270), .D(n_279), .Y(n_240) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx4_ASAP7_75t_SL g329 ( .A(n_243), .Y(n_329) );
INVx3_ASAP7_75t_SL g528 ( .A(n_243), .Y(n_528) );
INVx3_ASAP7_75t_L g579 ( .A(n_243), .Y(n_579) );
INVx6_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_253), .Y(n_244) );
AND2x4_ASAP7_75t_L g268 ( .A(n_245), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g286 ( .A(n_245), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g364 ( .A(n_245), .B(n_253), .Y(n_364) );
AND2x2_ASAP7_75t_L g370 ( .A(n_245), .B(n_269), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_245), .B(n_287), .Y(n_373) );
AND2x2_ASAP7_75t_L g404 ( .A(n_245), .B(n_287), .Y(n_404) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_251), .Y(n_245) );
INVx2_ASAP7_75t_L g265 ( .A(n_246), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_246), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_246), .Y(n_278) );
OAI22x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B1(n_249), .B2(n_250), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g252 ( .A(n_248), .Y(n_252) );
INVx2_ASAP7_75t_L g256 ( .A(n_248), .Y(n_256) );
INVx1_ASAP7_75t_L g259 ( .A(n_248), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g274 ( .A(n_251), .Y(n_274) );
BUFx2_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
AND2x2_ASAP7_75t_L g293 ( .A(n_253), .B(n_264), .Y(n_293) );
AND2x4_ASAP7_75t_L g301 ( .A(n_253), .B(n_297), .Y(n_301) );
AND2x4_ASAP7_75t_L g309 ( .A(n_253), .B(n_273), .Y(n_309) );
AND2x2_ASAP7_75t_L g380 ( .A(n_253), .B(n_297), .Y(n_380) );
AND2x2_ASAP7_75t_L g384 ( .A(n_253), .B(n_273), .Y(n_384) );
AND2x6_ASAP7_75t_L g387 ( .A(n_253), .B(n_264), .Y(n_387) );
AND2x2_ASAP7_75t_L g409 ( .A(n_253), .B(n_273), .Y(n_409) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g263 ( .A(n_255), .B(n_257), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_255), .B(n_258), .Y(n_277) );
INVx1_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
INVxp67_ASAP7_75t_L g269 ( .A(n_257), .Y(n_269) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g282 ( .A(n_258), .B(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g460 ( .A(n_262), .Y(n_460) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_262), .Y(n_543) );
BUFx2_ASAP7_75t_L g607 ( .A(n_262), .Y(n_607) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g305 ( .A(n_263), .B(n_297), .Y(n_305) );
AND2x4_ASAP7_75t_L g366 ( .A(n_263), .B(n_273), .Y(n_366) );
AND2x2_ASAP7_75t_L g369 ( .A(n_263), .B(n_264), .Y(n_369) );
AND2x2_ASAP7_75t_L g381 ( .A(n_263), .B(n_297), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_263), .B(n_264), .Y(n_402) );
AND2x2_ASAP7_75t_L g317 ( .A(n_264), .B(n_282), .Y(n_317) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_264), .B(n_282), .Y(n_377) );
AND2x2_ASAP7_75t_L g429 ( .A(n_264), .B(n_282), .Y(n_429) );
AND2x4_ASAP7_75t_L g297 ( .A(n_265), .B(n_274), .Y(n_297) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g337 ( .A(n_267), .Y(n_337) );
INVx2_ASAP7_75t_SL g477 ( .A(n_267), .Y(n_477) );
INVx2_ASAP7_75t_L g512 ( .A(n_267), .Y(n_512) );
INVx2_ASAP7_75t_L g583 ( .A(n_267), .Y(n_583) );
INVx2_ASAP7_75t_L g608 ( .A(n_267), .Y(n_608) );
INVx6_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx5_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g515 ( .A(n_272), .Y(n_515) );
BUFx3_ASAP7_75t_L g534 ( .A(n_272), .Y(n_534) );
AND2x2_ASAP7_75t_L g281 ( .A(n_273), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g372 ( .A(n_273), .B(n_282), .Y(n_372) );
BUFx12f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g458 ( .A(n_276), .Y(n_458) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x4_ASAP7_75t_L g312 ( .A(n_277), .B(n_297), .Y(n_312) );
AND2x4_ASAP7_75t_L g319 ( .A(n_277), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_277), .B(n_278), .Y(n_365) );
AND2x4_ASAP7_75t_L g378 ( .A(n_277), .B(n_320), .Y(n_378) );
AND2x4_ASAP7_75t_L g385 ( .A(n_277), .B(n_297), .Y(n_385) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_277), .B(n_278), .Y(n_399) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_281), .Y(n_334) );
INVx3_ASAP7_75t_L g472 ( .A(n_281), .Y(n_472) );
AND2x4_ASAP7_75t_L g296 ( .A(n_282), .B(n_297), .Y(n_296) );
AND2x6_ASAP7_75t_L g388 ( .A(n_282), .B(n_297), .Y(n_388) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
BUFx6f_ASAP7_75t_SL g470 ( .A(n_286), .Y(n_470) );
BUFx3_ASAP7_75t_L g540 ( .A(n_286), .Y(n_540) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND4xp25_ASAP7_75t_L g289 ( .A(n_290), .B(n_298), .C(n_306), .D(n_313), .Y(n_289) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_SL g346 ( .A(n_292), .Y(n_346) );
INVx2_ASAP7_75t_SL g448 ( .A(n_292), .Y(n_448) );
INVx2_ASAP7_75t_L g489 ( .A(n_292), .Y(n_489) );
INVx3_ASAP7_75t_L g587 ( .A(n_292), .Y(n_587) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g449 ( .A(n_295), .Y(n_449) );
INVx2_ASAP7_75t_L g483 ( .A(n_295), .Y(n_483) );
INVx2_ASAP7_75t_L g503 ( .A(n_295), .Y(n_503) );
INVx2_ASAP7_75t_L g562 ( .A(n_295), .Y(n_562) );
INVx2_ASAP7_75t_SL g588 ( .A(n_295), .Y(n_588) );
INVx8_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
INVx2_ASAP7_75t_SL g553 ( .A(n_300), .Y(n_553) );
INVx2_ASAP7_75t_L g592 ( .A(n_300), .Y(n_592) );
INVx3_ASAP7_75t_SL g618 ( .A(n_300), .Y(n_618) );
INVx3_ASAP7_75t_L g660 ( .A(n_300), .Y(n_660) );
INVx8_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g354 ( .A(n_305), .Y(n_354) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_305), .Y(n_412) );
INVx2_ASAP7_75t_L g491 ( .A(n_305), .Y(n_491) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g349 ( .A(n_308), .Y(n_349) );
INVx2_ASAP7_75t_L g486 ( .A(n_308), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_308), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_545) );
INVx6_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g614 ( .A(n_309), .Y(n_614) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g454 ( .A(n_311), .Y(n_454) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_SL g350 ( .A(n_312), .Y(n_350) );
BUFx3_ASAP7_75t_L g487 ( .A(n_312), .Y(n_487) );
BUFx3_ASAP7_75t_L g508 ( .A(n_312), .Y(n_508) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g655 ( .A(n_316), .Y(n_655) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_317), .Y(n_452) );
BUFx3_ASAP7_75t_L g481 ( .A(n_317), .Y(n_481) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx5_ASAP7_75t_SL g344 ( .A(n_319), .Y(n_344) );
BUFx2_ASAP7_75t_L g612 ( .A(n_319), .Y(n_612) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_338), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_327), .B(n_332), .Y(n_326) );
OAI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_330), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
NOR2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_347), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g566 ( .A(n_342), .Y(n_566) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g506 ( .A(n_344), .Y(n_506) );
OAI22xp33_ASAP7_75t_SL g564 ( .A1(n_344), .A2(n_565), .B1(n_567), .B2(n_568), .Y(n_564) );
INVx2_ASAP7_75t_L g656 ( .A(n_344), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g555 ( .A(n_350), .Y(n_555) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g438 ( .A(n_356), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_416), .B1(n_435), .B2(n_437), .Y(n_356) );
INVxp67_ASAP7_75t_L g437 ( .A(n_357), .Y(n_437) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_389), .B(n_414), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_359), .B(n_415), .Y(n_414) );
XNOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_374), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
INVx2_ASAP7_75t_SL g394 ( .A(n_364), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_366), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_382), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_379), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_391), .B(n_405), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_400), .Y(n_391) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_395), .B2(n_396), .C1(n_397), .C2(n_398), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g600 ( .A1(n_394), .A2(n_601), .B(n_602), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_394), .A2(n_663), .B(n_664), .C(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g603 ( .A(n_396), .Y(n_603) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
NOR2x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx2_ASAP7_75t_L g548 ( .A(n_412), .Y(n_548) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g436 ( .A(n_417), .Y(n_436) );
XOR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_434), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .Y(n_418) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_431), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g517 ( .A(n_439), .Y(n_517) );
OA22x2_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_497), .B2(n_498), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_463), .B1(n_495), .B2(n_496), .Y(n_441) );
INVx1_ASAP7_75t_L g495 ( .A(n_442), .Y(n_495) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_450), .C(n_451), .D(n_453), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .C(n_461), .D(n_462), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g468 ( .A(n_458), .Y(n_468) );
INVx3_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
INVx2_ASAP7_75t_L g496 ( .A(n_463), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_478), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_473), .C(n_475), .Y(n_465) );
NOR4xp25_ASAP7_75t_L g493 ( .A(n_466), .B(n_479), .C(n_484), .D(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g538 ( .A(n_472), .Y(n_538) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_474), .B(n_476), .Y(n_494) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_484), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .Y(n_484) );
BUFx2_ASAP7_75t_L g559 ( .A(n_489), .Y(n_559) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_516), .Y(n_498) );
NAND4xp75_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .C(n_509), .D(n_513), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g577 ( .A(n_515), .Y(n_577) );
INVx1_ASAP7_75t_L g621 ( .A(n_518), .Y(n_621) );
OAI22xp33_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_569), .B1(n_570), .B2(n_619), .Y(n_518) );
INVx1_ASAP7_75t_L g619 ( .A(n_519), .Y(n_619) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND3x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_544), .C(n_556), .Y(n_523) );
NOR2xp67_ASAP7_75t_SL g524 ( .A(n_525), .B(n_535), .Y(n_524) );
OAI21xp5_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_529), .B(n_530), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_541), .Y(n_535) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_554), .B2(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_564), .Y(n_556) );
OAI22xp33_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_560), .B1(n_561), .B2(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OA22x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_595), .B2(n_596), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_594), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_584), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
XNOR2x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_609), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_624), .B(n_627), .Y(n_672) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
OAI222xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_646), .B1(n_648), .B2(n_669), .C1(n_670), .C2(n_673), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_633), .Y(n_645) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .C(n_638), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .C(n_642), .D(n_643), .Y(n_639) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_669), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_661), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_657), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
CKINVDCx6p67_ASAP7_75t_R g671 ( .A(n_672), .Y(n_671) );
endmodule