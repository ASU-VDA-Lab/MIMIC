module fake_jpeg_10903_n_17 (n_3, n_2, n_1, n_0, n_4, n_17);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_17;

wire n_13;
wire n_11;
wire n_14;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

BUFx12f_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_7),
.B(n_1),
.Y(n_11)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_2),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_13),
.B(n_6),
.Y(n_14)
);

OAI32xp33_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_2),
.A3(n_8),
.B1(n_5),
.B2(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_12),
.Y(n_16)
);

AOI321xp33_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_5),
.A3(n_9),
.B1(n_15),
.B2(n_10),
.C(n_7),
.Y(n_17)
);


endmodule