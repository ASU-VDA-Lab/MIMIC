module real_jpeg_11472_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_229, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_229;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_35),
.B1(n_38),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_2),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_43),
.B1(n_61),
.B2(n_63),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_43),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_7),
.B(n_51),
.C(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_70),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_2),
.B(n_22),
.C(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_2),
.B(n_48),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_2),
.B(n_52),
.C(n_66),
.Y(n_189)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_35),
.B1(n_38),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_22),
.B1(n_28),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_9),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_116)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_41),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_11),
.A2(n_22),
.B1(n_28),
.B2(n_41),
.Y(n_141)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_16),
.B(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_73),
.C(n_83),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_17),
.B(n_73),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_44),
.B2(n_45),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_18),
.B(n_46),
.C(n_72),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_20),
.A2(n_32),
.B1(n_147),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_20),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_21),
.A2(n_25),
.B1(n_89),
.B2(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_25),
.A2(n_27),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_25),
.A2(n_87),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_25),
.B(n_43),
.Y(n_168)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_28),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_32),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_32),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_32),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_32),
.B(n_157),
.C(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_32),
.B(n_134),
.C(n_146),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_33),
.A2(n_39),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_33),
.Y(n_195)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_35),
.B(n_153),
.Y(n_152)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_38),
.A2(n_43),
.B(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_42),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_43),
.B(n_79),
.Y(n_170)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_46),
.A2(n_71),
.B1(n_90),
.B2(n_91),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_46),
.A2(n_71),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_46),
.B(n_96),
.C(n_194),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_54),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_47),
.A2(n_50),
.B1(n_94),
.B2(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B(n_52),
.C(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_58),
.A2(n_72),
.B1(n_117),
.B2(n_118),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_58),
.B(n_117),
.C(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_68),
.B(n_98),
.Y(n_97)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_63),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_70),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_91),
.C(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_82),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_81),
.B(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_79),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_83),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.C(n_96),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_84),
.A2(n_85),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_86),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_90),
.A2(n_91),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_91),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_96),
.A2(n_97),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_120),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B(n_119),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_117),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_118),
.B1(n_136),
.B2(n_142),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_118),
.B(n_137),
.C(n_140),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_222),
.B(n_226),
.Y(n_122)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_198),
.A3(n_217),
.B1(n_220),
.B2(n_221),
.C(n_229),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_181),
.B(n_197),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_148),
.B(n_180),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_127),
.B(n_133),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_128),
.A2(n_129),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_143),
.B2(n_144),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_174),
.B(n_179),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_161),
.B(n_173),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_159),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_170),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_187),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B(n_172),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_169),
.B(n_171),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_182),
.B(n_183),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.C(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_206),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_203),
.CI(n_205),
.CON(n_219),
.SN(n_219)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_214),
.C(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_225),
.Y(n_226)
);


endmodule