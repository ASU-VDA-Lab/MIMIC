module real_aes_10084_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g196 ( .A(n_0), .Y(n_196) );
INVx1_ASAP7_75t_L g599 ( .A(n_1), .Y(n_599) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_1), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_2), .A2(n_12), .B1(n_544), .B2(n_546), .Y(n_543) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_2), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_3), .B(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_4), .Y(n_204) );
INVx2_ASAP7_75t_L g487 ( .A(n_5), .Y(n_487) );
INVxp33_ASAP7_75t_SL g524 ( .A(n_6), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_6), .A2(n_50), .B1(n_571), .B2(n_579), .Y(n_570) );
BUFx2_ASAP7_75t_L g534 ( .A(n_7), .Y(n_534) );
BUFx2_ASAP7_75t_L g552 ( .A(n_7), .Y(n_552) );
INVx1_ASAP7_75t_L g595 ( .A(n_7), .Y(n_595) );
INVx1_ASAP7_75t_L g659 ( .A(n_8), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_9), .A2(n_72), .B1(n_538), .B2(n_541), .Y(n_537) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_9), .Y(n_617) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_10), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_10), .A2(n_47), .B1(n_624), .B2(n_628), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_11), .A2(n_70), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_11), .A2(n_70), .B1(n_571), .B2(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_12), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_13), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_14), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_15), .A2(n_16), .B1(n_541), .B2(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_15), .A2(n_16), .B1(n_588), .B2(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_17), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_18), .B(n_145), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_19), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_20), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_21), .B(n_112), .Y(n_186) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_23), .B(n_127), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_24), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_25), .B(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_26), .Y(n_92) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_27), .A2(n_94), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g532 ( .A(n_28), .Y(n_532) );
INVx1_ASAP7_75t_L g695 ( .A(n_28), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_29), .B(n_112), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_30), .Y(n_231) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_31), .A2(n_52), .B(n_120), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_32), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_33), .B(n_112), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_34), .Y(n_113) );
AND2x6_ASAP7_75t_L g84 ( .A(n_35), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_35), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_35), .B(n_678), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_36), .A2(n_64), .B1(n_147), .B2(n_184), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_37), .B(n_155), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_38), .Y(n_224) );
INVx1_ASAP7_75t_L g85 ( .A(n_39), .Y(n_85) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_39), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_40), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_41), .B(n_184), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_42), .B(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_43), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_44), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_45), .B(n_131), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_46), .B(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_46), .Y(n_669) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_47), .Y(n_518) );
INVx2_ASAP7_75t_L g205 ( .A(n_48), .Y(n_205) );
INVx1_ASAP7_75t_L g522 ( .A(n_49), .Y(n_522) );
INVxp33_ASAP7_75t_SL g496 ( .A(n_50), .Y(n_496) );
INVx2_ASAP7_75t_L g578 ( .A(n_51), .Y(n_578) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_53), .Y(n_663) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_54), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_55), .B(n_124), .Y(n_246) );
INVx1_ASAP7_75t_L g199 ( .A(n_56), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_57), .A2(n_479), .B1(n_480), .B2(n_698), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_57), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_58), .Y(n_129) );
BUFx10_ASAP7_75t_L g689 ( .A(n_59), .Y(n_689) );
INVx2_ASAP7_75t_L g598 ( .A(n_60), .Y(n_598) );
INVx1_ASAP7_75t_L g614 ( .A(n_60), .Y(n_614) );
INVx1_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_62), .B(n_124), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_63), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_65), .B(n_155), .Y(n_188) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_66), .Y(n_665) );
INVx1_ASAP7_75t_L g207 ( .A(n_67), .Y(n_207) );
INVxp33_ASAP7_75t_SL g495 ( .A(n_68), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_68), .A2(n_74), .B1(n_585), .B2(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g120 ( .A(n_69), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g290 ( .A(n_71), .B(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_71), .Y(n_670) );
INVxp67_ASAP7_75t_SL g632 ( .A(n_72), .Y(n_632) );
INVx2_ASAP7_75t_L g575 ( .A(n_73), .Y(n_575) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_74), .Y(n_507) );
BUFx3_ASAP7_75t_L g492 ( .A(n_75), .Y(n_492) );
INVx1_ASAP7_75t_L g528 ( .A(n_75), .Y(n_528) );
BUFx3_ASAP7_75t_L g494 ( .A(n_76), .Y(n_494) );
INVx1_ASAP7_75t_L g501 ( .A(n_76), .Y(n_501) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_77), .B(n_155), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_96), .B(n_477), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_83), .A2(n_131), .B(n_132), .Y(n_130) );
INVx8_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
INVx2_ASAP7_75t_SL g248 ( .A(n_83), .Y(n_248) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g173 ( .A(n_84), .Y(n_173) );
AOI21xp33_ASAP7_75t_L g208 ( .A1(n_84), .A2(n_117), .B(n_206), .Y(n_208) );
INVx1_ASAP7_75t_L g228 ( .A(n_84), .Y(n_228) );
INVxp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g711 ( .A1(n_87), .A2(n_712), .B(n_713), .Y(n_711) );
NAND2xp33_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g184 ( .A(n_91), .Y(n_184) );
INVx2_ASAP7_75t_L g203 ( .A(n_91), .Y(n_203) );
INVx2_ASAP7_75t_L g292 ( .A(n_91), .Y(n_292) );
INVx2_ASAP7_75t_L g294 ( .A(n_91), .Y(n_294) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g110 ( .A(n_92), .Y(n_110) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_92), .Y(n_112) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_92), .Y(n_128) );
INVx2_ASAP7_75t_L g148 ( .A(n_92), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_93), .A2(n_195), .B(n_198), .Y(n_194) );
BUFx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_94), .Y(n_114) );
INVx3_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_94), .B(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_94), .A2(n_290), .B1(n_293), .B2(n_295), .Y(n_289) );
BUFx12f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx5_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
INVx5_ASAP7_75t_L g163 ( .A(n_95), .Y(n_163) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND3x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_361), .C(n_434), .Y(n_97) );
NOR2xp67_ASAP7_75t_L g98 ( .A(n_99), .B(n_269), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_100), .B(n_250), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_189), .B(n_209), .C(n_235), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_133), .Y(n_101) );
INVx1_ASAP7_75t_L g211 ( .A(n_102), .Y(n_211) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g216 ( .A(n_104), .Y(n_216) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g254 ( .A(n_105), .Y(n_254) );
INVx1_ASAP7_75t_L g279 ( .A(n_105), .Y(n_279) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_121), .B(n_130), .Y(n_105) );
AO21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_114), .B(n_115), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_109), .B1(n_111), .B2(n_113), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g197 ( .A(n_111), .Y(n_197) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
AOI21x1_ASAP7_75t_L g121 ( .A1(n_114), .A2(n_122), .B(n_125), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_114), .A2(n_201), .B(n_206), .Y(n_200) );
INVxp67_ASAP7_75t_L g132 ( .A(n_115), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx3_ASAP7_75t_L g131 ( .A(n_117), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_117), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_123), .A2(n_479), .B1(n_480), .B2(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_123), .Y(n_705) );
INVx5_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVxp67_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_127), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g225 ( .A(n_128), .Y(n_225) );
INVx1_ASAP7_75t_L g714 ( .A(n_129), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_133), .A2(n_447), .B1(n_449), .B2(n_451), .Y(n_446) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_157), .Y(n_133) );
AND2x4_ASAP7_75t_L g320 ( .A(n_134), .B(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g212 ( .A(n_135), .B(n_174), .Y(n_212) );
INVx2_ASAP7_75t_L g336 ( .A(n_135), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_135), .B(n_268), .Y(n_355) );
AND2x2_ASAP7_75t_L g371 ( .A(n_135), .B(n_158), .Y(n_371) );
AND2x2_ASAP7_75t_L g467 ( .A(n_135), .B(n_279), .Y(n_467) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
OAI21x1_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_152), .B(n_154), .Y(n_136) );
OAI21x1_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_143), .B(n_151), .Y(n_137) );
AOI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_142), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_149), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_147), .B1(n_165), .B2(n_166), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_145), .A2(n_202), .B1(n_204), .B2(n_205), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_147), .A2(n_224), .B1(n_225), .B2(n_226), .Y(n_223) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx1_ASAP7_75t_L g232 ( .A(n_148), .Y(n_232) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_150), .A2(n_186), .B(n_187), .Y(n_185) );
OAI21xp33_ASAP7_75t_L g222 ( .A1(n_150), .A2(n_223), .B(n_227), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_151), .A2(n_180), .B(n_185), .Y(n_179) );
AO31x2_ASAP7_75t_L g287 ( .A1(n_151), .A2(n_288), .A3(n_289), .B(n_296), .Y(n_287) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_152), .A2(n_240), .B(n_249), .Y(n_239) );
BUFx4f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_153), .B(n_228), .Y(n_227) );
NOR2x1p5_ASAP7_75t_SL g172 ( .A(n_155), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g288 ( .A(n_155), .Y(n_288) );
BUFx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g298 ( .A(n_156), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_157), .B(n_278), .Y(n_406) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_174), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_158), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g283 ( .A(n_158), .Y(n_283) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g257 ( .A(n_159), .Y(n_257) );
HB1xp67_ASAP7_75t_SL g281 ( .A(n_159), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_159), .B(n_279), .Y(n_310) );
AND2x2_ASAP7_75t_L g325 ( .A(n_159), .B(n_258), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_159), .B(n_268), .Y(n_326) );
INVx1_ASAP7_75t_L g354 ( .A(n_159), .Y(n_354) );
AND2x2_ASAP7_75t_L g377 ( .A(n_159), .B(n_216), .Y(n_377) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_167), .C(n_172), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_162), .A2(n_181), .B(n_183), .Y(n_180) );
CKINVDCx6p67_ASAP7_75t_R g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_SL g171 ( .A(n_163), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_163), .A2(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_SL g247 ( .A(n_163), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_171), .Y(n_167) );
BUFx2_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
AND2x4_ASAP7_75t_L g335 ( .A(n_174), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g370 ( .A(n_174), .Y(n_370) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x4_ASAP7_75t_L g321 ( .A(n_175), .B(n_254), .Y(n_321) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
OAI21x1_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_179), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_189), .B(n_286), .Y(n_452) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g372 ( .A(n_190), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_190), .B(n_360), .Y(n_448) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_191), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g418 ( .A(n_191), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_191), .B(n_419), .Y(n_445) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g260 ( .A(n_192), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g384 ( .A(n_192), .B(n_253), .Y(n_384) );
AND2x2_ASAP7_75t_L g393 ( .A(n_192), .B(n_317), .Y(n_393) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g220 ( .A(n_193), .Y(n_220) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_200), .B(n_208), .Y(n_193) );
NOR2x1_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21xp33_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_213), .B(n_217), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_212), .A2(n_275), .B(n_280), .C(n_282), .Y(n_274) );
AND2x2_ASAP7_75t_L g376 ( .A(n_212), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_212), .B(n_281), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_212), .B(n_430), .Y(n_429) );
OAI222xp33_ASAP7_75t_L g471 ( .A1(n_213), .A2(n_272), .B1(n_389), .B2(n_472), .C1(n_473), .C2(n_476), .Y(n_471) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x4_ASAP7_75t_L g255 ( .A(n_214), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g282 ( .A(n_214), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g414 ( .A(n_214), .Y(n_414) );
INVx2_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_217), .A2(n_400), .B(n_402), .C(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_218), .A2(n_251), .B1(n_259), .B2(n_262), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_218), .A2(n_410), .B1(n_411), .B2(n_412), .Y(n_409) );
AND2x2_ASAP7_75t_L g455 ( .A(n_218), .B(n_286), .Y(n_455) );
BUFx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g390 ( .A(n_219), .B(n_360), .Y(n_390) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
OR2x2_ASAP7_75t_L g300 ( .A(n_220), .B(n_221), .Y(n_300) );
INVx2_ASAP7_75t_L g306 ( .A(n_220), .Y(n_306) );
INVx2_ASAP7_75t_SL g261 ( .A(n_221), .Y(n_261) );
AND2x2_ASAP7_75t_L g305 ( .A(n_221), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g345 ( .A(n_221), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_221), .Y(n_358) );
INVx1_ASAP7_75t_L g374 ( .A(n_221), .Y(n_374) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_229), .B(n_234), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_225), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g259 ( .A(n_237), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
OR2x2_ASAP7_75t_L g395 ( .A(n_237), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_237), .B(n_343), .Y(n_470) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x4_ASAP7_75t_L g286 ( .A(n_238), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g379 ( .A(n_238), .B(n_331), .Y(n_379) );
BUFx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B(n_248), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_247), .Y(n_244) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
AND2x2_ASAP7_75t_L g273 ( .A(n_252), .B(n_256), .Y(n_273) );
OR2x2_ASAP7_75t_L g368 ( .A(n_252), .B(n_324), .Y(n_368) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_252), .Y(n_442) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_255), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g462 ( .A(n_255), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g265 ( .A(n_256), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g383 ( .A(n_256), .B(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g388 ( .A(n_256), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_256), .B(n_321), .Y(n_450) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_258), .B(n_268), .Y(n_349) );
INVx2_ASAP7_75t_L g339 ( .A(n_260), .Y(n_339) );
AND2x4_ASAP7_75t_SL g378 ( .A(n_260), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g425 ( .A(n_260), .B(n_304), .Y(n_425) );
AND2x2_ASAP7_75t_L g329 ( .A(n_261), .B(n_317), .Y(n_329) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g333 ( .A(n_264), .B(n_326), .Y(n_333) );
INVx2_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g308 ( .A(n_267), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g423 ( .A(n_267), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g428 ( .A(n_267), .B(n_353), .Y(n_428) );
AND2x2_ASAP7_75t_L g433 ( .A(n_267), .B(n_325), .Y(n_433) );
AND2x2_ASAP7_75t_L g454 ( .A(n_267), .B(n_377), .Y(n_454) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_307), .C(n_340), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_301), .Y(n_270) );
AOI21xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_274), .B(n_284), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
BUFx2_ASAP7_75t_L g422 ( .A(n_277), .Y(n_422) );
INVx1_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g353 ( .A(n_279), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_283), .B(n_355), .Y(n_382) );
AND2x4_ASAP7_75t_SL g466 ( .A(n_283), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_285), .A2(n_341), .B1(n_343), .B2(n_347), .C(n_350), .Y(n_340) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_299), .Y(n_285) );
INVx2_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g401 ( .A(n_286), .Y(n_401) );
AND2x2_ASAP7_75t_L g432 ( .A(n_286), .B(n_305), .Y(n_432) );
INVx1_ASAP7_75t_L g315 ( .A(n_287), .Y(n_315) );
INVx2_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
INVx2_ASAP7_75t_SL g346 ( .A(n_287), .Y(n_346) );
AND2x2_ASAP7_75t_L g360 ( .A(n_287), .B(n_317), .Y(n_360) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g380 ( .A(n_299), .B(n_313), .Y(n_380) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g404 ( .A(n_300), .Y(n_404) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g476 ( .A(n_303), .Y(n_476) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g463 ( .A(n_304), .B(n_373), .Y(n_463) );
AND2x4_ASAP7_75t_L g330 ( .A(n_306), .B(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_306), .Y(n_344) );
AOI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_311), .B(n_318), .C(n_332), .Y(n_307) );
INVx1_ASAP7_75t_L g363 ( .A(n_308), .Y(n_363) );
AND2x2_ASAP7_75t_L g347 ( .A(n_309), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g415 ( .A(n_310), .Y(n_415) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_314), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_314), .Y(n_408) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g373 ( .A(n_315), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g440 ( .A(n_317), .Y(n_440) );
AOI31xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .A3(n_326), .B(n_327), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_320), .A2(n_392), .B1(n_394), .B2(n_397), .Y(n_391) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g417 ( .A(n_329), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_329), .B(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_337), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_333), .A2(n_351), .B(n_356), .Y(n_350) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_335), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
OR2x6_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVxp67_ASAP7_75t_L g385 ( .A(n_338), .Y(n_385) );
OR2x6_ASAP7_75t_L g458 ( .A(n_342), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g475 ( .A(n_344), .Y(n_475) );
AND2x2_ASAP7_75t_L g392 ( .A(n_345), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g396 ( .A(n_345), .Y(n_396) );
AND2x2_ASAP7_75t_L g474 ( .A(n_345), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g419 ( .A(n_346), .Y(n_419) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g424 ( .A(n_353), .Y(n_424) );
AND2x2_ASAP7_75t_L g411 ( .A(n_355), .B(n_377), .Y(n_411) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_386), .C(n_407), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_375), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_372), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_369), .A2(n_437), .B1(n_441), .B2(n_443), .Y(n_436) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx2_ASAP7_75t_L g459 ( .A(n_371), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_380), .B2(n_381), .C1(n_383), .C2(n_385), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_391), .C(n_399), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_388), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g457 ( .A(n_392), .Y(n_457) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_395), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g438 ( .A(n_396), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_403), .A2(n_430), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g410 ( .A(n_404), .Y(n_410) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI211xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_409), .B(n_416), .C(n_431), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B1(n_425), .B2(n_426), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_417), .A2(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_460), .C(n_471), .Y(n_434) );
NAND3xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_446), .C(n_453), .Y(n_435) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI21xp33_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_455), .B(n_456), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_468), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g472 ( .A(n_467), .Y(n_472) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_674), .B1(n_697), .B2(n_699), .C(n_703), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_650), .B2(n_651), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_535), .C(n_615), .Y(n_481) );
AOI31xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_506), .A3(n_521), .B(n_529), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_495), .B1(n_496), .B2(n_497), .C(n_502), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .Y(n_484) );
AND2x6_ASAP7_75t_L g525 ( .A(n_485), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g499 ( .A(n_487), .Y(n_499) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
INVx2_ASAP7_75t_L g554 ( .A(n_487), .Y(n_554) );
AND2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_532), .Y(n_567) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g540 ( .A(n_489), .Y(n_540) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_489), .Y(n_558) );
INVx6_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g523 ( .A(n_490), .B(n_513), .Y(n_523) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g520 ( .A(n_491), .Y(n_520) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g500 ( .A(n_492), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g505 ( .A(n_492), .B(n_494), .Y(n_505) );
INVx1_ASAP7_75t_L g517 ( .A(n_493), .Y(n_517) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g527 ( .A(n_494), .B(n_528), .Y(n_527) );
AND2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g503 ( .A(n_498), .Y(n_503) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x6_ASAP7_75t_L g519 ( .A(n_499), .B(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_500), .Y(n_545) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_504), .Y(n_542) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_505), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_511), .B2(n_512), .C1(n_518), .C2(n_519), .Y(n_506) );
BUFx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_SL g512 ( .A(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g687 ( .A(n_517), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_522), .A2(n_632), .B1(n_633), .B2(n_637), .Y(n_631) );
INVx1_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g553 ( .A(n_532), .B(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g568 ( .A(n_534), .Y(n_568) );
NAND4xp25_ASAP7_75t_L g535 ( .A(n_536), .B(n_555), .C(n_569), .D(n_600), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .C(n_550), .Y(n_536) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OR2x6_ASAP7_75t_L g648 ( .A(n_552), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g693 ( .A(n_554), .B(n_694), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .C(n_564), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx4f_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_565), .Y(n_564) );
OR2x6_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_SL g683 ( .A(n_567), .Y(n_683) );
AND2x4_ASAP7_75t_L g610 ( .A(n_568), .B(n_611), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_584), .C(n_592), .Y(n_569) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g642 ( .A(n_573), .B(n_639), .Y(n_642) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g582 ( .A(n_575), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g587 ( .A(n_575), .B(n_578), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_575), .Y(n_591) );
INVx1_ASAP7_75t_L g630 ( .A(n_575), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_575), .B(n_578), .Y(n_636) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g583 ( .A(n_578), .Y(n_583) );
INVx1_ASAP7_75t_L g627 ( .A(n_578), .Y(n_627) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g605 ( .A(n_582), .Y(n_605) );
INVx1_ASAP7_75t_L g646 ( .A(n_582), .Y(n_646) );
AND2x4_ASAP7_75t_L g590 ( .A(n_583), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g609 ( .A(n_586), .Y(n_609) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx3_ASAP7_75t_L g619 ( .A(n_590), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_590), .B(n_621), .Y(n_620) );
INVx5_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x6_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g640 ( .A(n_598), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .C(n_610), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_612), .Y(n_649) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_SL g626 ( .A(n_614), .Y(n_626) );
OR2x2_ASAP7_75t_L g628 ( .A(n_614), .B(n_629), .Y(n_628) );
AOI31xp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_631), .A3(n_641), .B(n_648), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_620), .C(n_623), .Y(n_616) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
OR2x6_ASAP7_75t_L g634 ( .A(n_626), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx8_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x6_ASAP7_75t_L g638 ( .A(n_635), .B(n_639), .Y(n_638) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx4_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g644 ( .A(n_639), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_647), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_661), .B1(n_672), .B2(n_673), .Y(n_651) );
INVx1_ASAP7_75t_L g672 ( .A(n_652), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g660 ( .A(n_653), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_653) );
INVx4_ASAP7_75t_L g657 ( .A(n_654), .Y(n_657) );
INVx1_ASAP7_75t_L g656 ( .A(n_655), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g673 ( .A(n_661), .Y(n_673) );
XOR2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_667), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_663), .Y(n_666) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_670), .Y(n_671) );
INVx8_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x6_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
OR2x4_ASAP7_75t_L g709 ( .A(n_677), .B(n_681), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_678), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g712 ( .A(n_678), .Y(n_712) );
INVx1_ASAP7_75t_L g702 ( .A(n_679), .Y(n_702) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .A3(n_688), .B(n_690), .Y(n_681) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g696 ( .A(n_687), .Y(n_696) );
INVx6_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B1(n_710), .B2(n_714), .Y(n_703) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx8_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
endmodule