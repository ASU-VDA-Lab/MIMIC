module fake_jpeg_15336_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_63),
.B1(n_64),
.B2(n_29),
.Y(n_67)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_21),
.B(n_34),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_34),
.B1(n_17),
.B2(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_45),
.B1(n_29),
.B2(n_19),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_34),
.B1(n_17),
.B2(n_20),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_86),
.B1(n_88),
.B2(n_98),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_42),
.Y(n_81)
);

NOR2x1_ASAP7_75t_R g108 ( 
.A(n_82),
.B(n_16),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_35),
.B1(n_40),
.B2(n_45),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_40),
.B1(n_45),
.B2(n_38),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_25),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_56),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_40),
.B1(n_32),
.B2(n_18),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_38),
.Y(n_101)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_33),
.B(n_30),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_44),
.C(n_37),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_86),
.C(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_32),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_30),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_37),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_133),
.C(n_139),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_67),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_101),
.B1(n_90),
.B2(n_73),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_134),
.A2(n_116),
.B1(n_23),
.B2(n_24),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_68),
.B1(n_77),
.B2(n_73),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_147),
.B1(n_154),
.B2(n_162),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_109),
.B(n_131),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_68),
.B1(n_80),
.B2(n_74),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_158),
.B1(n_110),
.B2(n_106),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_100),
.C(n_96),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_74),
.B(n_30),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_119),
.B(n_104),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_75),
.B1(n_85),
.B2(n_70),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_89),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_157),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_75),
.B1(n_23),
.B2(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_28),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_14),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_94),
.B1(n_72),
.B2(n_26),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_124),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_23),
.B1(n_28),
.B2(n_24),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_112),
.CI(n_125),
.CON(n_166),
.SN(n_166)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_170),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_124),
.B(n_104),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_173),
.B(n_178),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_184),
.B1(n_87),
.B2(n_24),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

XNOR2x2_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_126),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_181),
.C(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_117),
.C(n_102),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_105),
.C(n_44),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_39),
.B(n_16),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_44),
.C(n_123),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_188),
.C(n_39),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_87),
.C(n_131),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_130),
.B1(n_116),
.B2(n_28),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_0),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_194),
.B(n_16),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_142),
.B(n_136),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_72),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_137),
.B1(n_150),
.B2(n_138),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_204),
.B1(n_207),
.B2(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_150),
.B1(n_144),
.B2(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_174),
.B1(n_177),
.B2(n_181),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_208),
.B(n_179),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_166),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_143),
.B1(n_140),
.B2(n_26),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_87),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_223),
.C(n_180),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_169),
.B1(n_190),
.B2(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_173),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_193),
.B1(n_176),
.B2(n_169),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_164),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_222),
.B1(n_163),
.B2(n_167),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_39),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_1),
.B(n_2),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_194),
.B(n_2),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_195),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_247),
.C(n_205),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_243),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_225),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_1),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_208),
.B(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_240),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_245),
.B(n_201),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_204),
.B1(n_229),
.B2(n_203),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_182),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_202),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_175),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_196),
.B1(n_26),
.B2(n_4),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_250),
.A2(n_224),
.B1(n_217),
.B2(n_211),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_211),
.B1(n_201),
.B2(n_199),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_262),
.C(n_265),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_218),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_263),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_245),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_214),
.C(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_199),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_197),
.B1(n_207),
.B2(n_209),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_213),
.C(n_226),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_226),
.B1(n_11),
.B2(n_12),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_232),
.B1(n_266),
.B2(n_255),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_3),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_237),
.B(n_240),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_283),
.B(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_243),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_236),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.C(n_251),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_261),
.B(n_254),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_262),
.C(n_265),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_293),
.C(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_230),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_295),
.C(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_270),
.C(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_232),
.C(n_257),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_260),
.B(n_250),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_39),
.C(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_39),
.C(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_3),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_271),
.B(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_291),
.A2(n_272),
.B1(n_278),
.B2(n_279),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_309),
.C(n_292),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_286),
.B(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_11),
.B(n_6),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_9),
.B(n_6),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_6),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_295),
.B(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_7),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_315),
.C(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_325),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_303),
.B(n_307),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_316),
.B(n_8),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_328),
.C(n_323),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_7),
.B(n_8),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_327),
.B(n_13),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_7),
.C(n_13),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_14),
.C(n_15),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_15),
.C(n_39),
.Y(n_333)
);


endmodule