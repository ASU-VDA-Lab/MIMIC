module fake_jpeg_20364_n_210 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_1),
.B(n_3),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_24),
.Y(n_93)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2x1_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_18),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_29),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_24),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_45),
.B1(n_26),
.B2(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_20),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_16),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_30),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_76),
.B1(n_79),
.B2(n_90),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_52),
.B(n_5),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_43),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

XOR2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_17),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_63),
.C(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_43),
.B1(n_32),
.B2(n_25),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_93),
.B(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_69),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_80),
.B1(n_78),
.B2(n_54),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_110),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_12),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_13),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_136),
.B1(n_119),
.B2(n_105),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_82),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_93),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_79),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_138),
.B(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_93),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_96),
.B1(n_83),
.B2(n_78),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_86),
.B(n_96),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_130),
.B1(n_135),
.B2(n_126),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_121),
.B1(n_138),
.B2(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_111),
.C(n_99),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_111),
.C(n_99),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_112),
.C(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_159),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_140),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_114),
.B(n_100),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_110),
.B(n_81),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_167),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_127),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_170),
.C(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_143),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_144),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_149),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_153),
.B(n_160),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_148),
.B(n_151),
.Y(n_181)
);

AOI321xp33_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_158),
.A3(n_142),
.B1(n_10),
.B2(n_116),
.C(n_85),
.Y(n_182)
);

AOI31xp67_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_183),
.A3(n_161),
.B(n_174),
.Y(n_190)
);

BUFx12f_ASAP7_75t_SL g183 ( 
.A(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_158),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_168),
.B1(n_167),
.B2(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_169),
.C(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

AOI321xp33_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_169),
.A3(n_173),
.B1(n_164),
.B2(n_54),
.C(n_51),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_60),
.C(n_59),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_195),
.B(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_4),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_60),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_186),
.C(n_55),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_203),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_186),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_204),
.C(n_7),
.Y(n_207)
);

AOI22x1_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_204)
);

AOI31xp33_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_195),
.A3(n_196),
.B(n_9),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_205),
.B(n_200),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);


endmodule