module real_jpeg_26990_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_0),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_190),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_190),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_57),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_169),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_169),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_169),
.Y(n_266)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_60),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_8),
.B(n_47),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_8),
.A2(n_47),
.B(n_226),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_188),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_8),
.A2(n_31),
.B(n_34),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_138),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_8),
.A2(n_87),
.B1(n_90),
.B2(n_274),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_9),
.A2(n_34),
.B1(n_36),
.B2(n_66),
.Y(n_203)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_54),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_12),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_142),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_142),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_12),
.A2(n_34),
.B1(n_36),
.B2(n_142),
.Y(n_261)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_116),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_20),
.B(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_84),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_21),
.A2(n_22),
.B1(n_74),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_22)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_24),
.A2(n_25),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_41),
.C(n_58),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_37),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_26),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_26),
.A2(n_33),
.B1(n_95),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_26),
.A2(n_37),
.B(n_96),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_26),
.A2(n_33),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_79),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_26),
.A2(n_33),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_26),
.A2(n_33),
.B1(n_233),
.B2(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_28),
.A2(n_48),
.A3(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_224)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_45),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_29),
.A2(n_32),
.B(n_188),
.C(n_253),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_33),
.A2(n_81),
.B(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_33),
.B(n_188),
.Y(n_272)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_36),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_38),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_52),
.B(n_55),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_42),
.A2(n_55),
.B(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_42),
.A2(n_110),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_51),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_43),
.B(n_56),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_43),
.A2(n_51),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_43),
.A2(n_51),
.B1(n_184),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_43),
.A2(n_51),
.B1(n_212),
.B2(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_45),
.Y(n_225)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_47),
.B(n_61),
.Y(n_201)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_48),
.A2(n_69),
.B1(n_187),
.B2(n_201),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_73),
.B1(n_102),
.B2(n_114),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B(n_67),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_63),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_59),
.A2(n_104),
.B1(n_141),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_59),
.A2(n_104),
.B1(n_168),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_61),
.B(n_65),
.C(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_60),
.B(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_60),
.A2(n_68),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_65),
.B(n_188),
.CON(n_187),
.SN(n_187)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_77),
.A2(n_112),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_84),
.A2(n_85),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_93),
.B(n_97),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_97),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_86),
.A2(n_94),
.B1(n_123),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_87),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_87),
.A2(n_134),
.B1(n_160),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_87),
.A2(n_132),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_87),
.A2(n_90),
.B1(n_266),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_88),
.A2(n_92),
.B(n_162),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_88),
.A2(n_133),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_89),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_131),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_90),
.A2(n_129),
.B(n_203),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_94),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_113),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_141),
.B(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_148),
.B(n_319),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_144),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_119),
.B(n_144),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_124),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_125),
.A2(n_126),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_139),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_128),
.B(n_135),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_173),
.B(n_318),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_170),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_150),
.B(n_170),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_155),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_157),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.C(n_166),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_158),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_163),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_312),
.B(n_317),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_216),
.B(n_298),
.C(n_311),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_204),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_176),
.B(n_204),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_178),
.B(n_179),
.C(n_191),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_186),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_193),
.B(n_197),
.C(n_199),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_202),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_210),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_205),
.A2(n_206),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_297),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_290),
.B(n_296),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_244),
.B(n_289),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_220),
.B(n_235),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.C(n_231),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_221),
.A2(n_222),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_236),
.B(n_242),
.C(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_283),
.B(n_288),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_262),
.B(n_282),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_249),
.B1(n_252),
.B2(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_281),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_268),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_275),
.B(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_309),
.B2(n_310),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_306),
.C(n_310),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule