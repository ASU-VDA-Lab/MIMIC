module real_jpeg_30194_n_18 (n_17, n_8, n_0, n_2, n_331, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_331;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_0),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_29),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_0),
.B(n_31),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_0),
.A2(n_55),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_0),
.B(n_55),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_68),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_0),
.A2(n_132),
.B1(n_134),
.B2(n_200),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_0),
.A2(n_32),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_92),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_92),
.Y(n_220)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_5),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_97),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_50),
.B1(n_52),
.B2(n_97),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_153)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_9),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_9),
.A2(n_50),
.B1(n_52),
.B2(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_27),
.B1(n_50),
.B2(n_52),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_10),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_11),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_90),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_90),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_50),
.B1(n_52),
.B2(n_90),
.Y(n_193)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_107),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_50),
.B1(n_52),
.B2(n_107),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_17),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_17),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_34),
.B(n_104),
.C(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_28),
.A2(n_31),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_31),
.B1(n_141),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_28),
.A2(n_31),
.B1(n_160),
.B2(n_255),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_62),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_32),
.A2(n_56),
.A3(n_62),
.B1(n_217),
.B2(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_33),
.B(n_104),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_38),
.A2(n_39),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_40),
.B(n_314),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_282),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_46),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_46),
.A2(n_58),
.B1(n_308),
.B2(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_53),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_47),
.A2(n_53),
.B1(n_130),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_47),
.A2(n_53),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_47),
.A2(n_53),
.B1(n_174),
.B2(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_104),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_47),
.A2(n_53),
.B1(n_96),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_47),
.A2(n_53),
.B1(n_57),
.B2(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_48),
.A2(n_52),
.A3(n_55),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_49),
.B(n_50),
.Y(n_178)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_50),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_55),
.B(n_66),
.Y(n_225)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_68),
.B1(n_89),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_68),
.B1(n_144),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_60),
.A2(n_68),
.B1(n_162),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_65),
.B1(n_88),
.B2(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_65),
.B1(n_91),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_61),
.A2(n_65),
.B1(n_121),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_61),
.A2(n_65),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_69),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_73),
.A2(n_75),
.B1(n_106),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_73),
.A2(n_75),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_322),
.B(n_328),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_299),
.A3(n_318),
.B1(n_320),
.B2(n_321),
.C(n_331),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_251),
.A3(n_288),
.B1(n_293),
.B2(n_298),
.C(n_332),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_146),
.C(n_164),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_125),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_83),
.B(n_125),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_108),
.C(n_117),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_84),
.B(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_102),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_94),
.C(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_98),
.A2(n_101),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_98),
.A2(n_101),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_134),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_249),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_108),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_111),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_112),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g201 ( 
.A(n_113),
.Y(n_201)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_119),
.B(n_236),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_122),
.B(n_124),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_136),
.C(n_137),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_134),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_132),
.A2(n_193),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_132),
.A2(n_134),
.B1(n_188),
.B2(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_132),
.A2(n_134),
.B(n_153),
.Y(n_266)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.C(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_147),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_148),
.B(n_149),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_151),
.B(n_156),
.C(n_163),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_152),
.B(n_154),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_155),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_245),
.B(n_250),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_231),
.B(n_244),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_210),
.B(n_230),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_189),
.B(n_209),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_197),
.B(n_208),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_203),
.B(n_207),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_223),
.B1(n_228),
.B2(n_229),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_222),
.C(n_229),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_240),
.C(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_268),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.C(n_267),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_259),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_253),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.CI(n_258),
.CON(n_253),
.SN(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_256),
.C(n_258),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_255),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_257),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_266),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_266),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_266),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_280),
.B(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_286),
.B2(n_287),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_277),
.C(n_287),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_275),
.B(n_276),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_274),
.Y(n_306)
);

FAx1_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_301),
.CI(n_310),
.CON(n_300),
.SN(n_300)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_311),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_311),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_309),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_303),
.B1(n_313),
.B2(n_316),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.C(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_316),
.C(n_317),
.Y(n_323)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);


endmodule