module fake_netlist_5_1691_n_1153 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1153);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1153;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_1060;
wire n_851;
wire n_1141;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1048;
wire n_932;
wire n_417;
wire n_1008;
wire n_946;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_259;
wire n_448;
wire n_999;
wire n_758;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_1049;
wire n_992;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_919;
wire n_782;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_900;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_1020;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_897;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_1070;
wire n_777;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_1064;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_996;
wire n_921;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_1089;
wire n_1138;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_890;
wire n_1032;
wire n_1056;
wire n_960;
wire n_764;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_38),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_21),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_25),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_8),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_40),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_42),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_118),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_130),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_29),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_44),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_93),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_131),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_86),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_106),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_194),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_46),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_39),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_50),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_88),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_18),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_120),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_196),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_183),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_62),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_2),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_169),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_105),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_174),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_158),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_186),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_76),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_108),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_111),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_221),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_156),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_87),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_137),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_113),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_209),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_222),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_240),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_283),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_242),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_257),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_248),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_232),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_275),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_233),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_225),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_256),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_225),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_229),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_235),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_245),
.B(n_239),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_258),
.B1(n_259),
.B2(n_272),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_258),
.B1(n_259),
.B2(n_272),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_278),
.B1(n_288),
.B2(n_255),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_293),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_335),
.A2(n_249),
.B(n_247),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_250),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_252),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_253),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_292),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_278),
.B1(n_288),
.B2(n_289),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_330),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_295),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_332),
.A2(n_266),
.B(n_265),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_291),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_33),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_286),
.B1(n_285),
.B2(n_284),
.Y(n_378)
);

CKINVDCx11_ASAP7_75t_R g379 ( 
.A(n_294),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_328),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_297),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_321),
.B(n_268),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_303),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_269),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_R g393 ( 
.A(n_315),
.B(n_0),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_326),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_315),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_336),
.A2(n_273),
.B(n_271),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_379),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_276),
.B(n_274),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_390),
.B(n_294),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_379),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_390),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_352),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_380),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_356),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_345),
.Y(n_412)
);

AOI21x1_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_281),
.B(n_279),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_282),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_391),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_358),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_378),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_351),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_360),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

OR2x6_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_396),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

BUFx3_ASAP7_75t_SL g428 ( 
.A(n_377),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_347),
.B(n_0),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_365),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_365),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_353),
.B(n_1),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_393),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_393),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_392),
.B(n_304),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_392),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_363),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_348),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_363),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_363),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_375),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_389),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_375),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_375),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_1),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_395),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_389),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

AO22x2_ASAP7_75t_L g454 ( 
.A1(n_370),
.A2(n_395),
.B1(n_397),
.B2(n_394),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_374),
.Y(n_455)
);

AND3x2_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_2),
.C(n_3),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_371),
.B(n_304),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_374),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_343),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_377),
.B(n_317),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_343),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_382),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_R g468 ( 
.A(n_377),
.B(n_317),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_34),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_355),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_449),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_426),
.B(n_343),
.Y(n_477)
);

NOR2x1p5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_371),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_415),
.B(n_361),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_419),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_400),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_422),
.B(n_457),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_423),
.B(n_373),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_371),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_373),
.Y(n_496)
);

INVx8_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_388),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_418),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_400),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_440),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_367),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_436),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_437),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_451),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_467),
.B(n_367),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_377),
.B1(n_387),
.B2(n_384),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_384),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_372),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_368),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_421),
.A2(n_372),
.B1(n_387),
.B2(n_384),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_410),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_455),
.B(n_368),
.Y(n_516)
);

INVx4_ASAP7_75t_SL g517 ( 
.A(n_425),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_435),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_463),
.B(n_384),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_425),
.B(n_387),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_466),
.B(n_388),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_408),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_454),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_428),
.B(n_377),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_445),
.B(n_387),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_448),
.B(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_443),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_411),
.B(n_381),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_441),
.B(n_381),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_433),
.B(n_381),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_405),
.B(n_3),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_433),
.B(n_366),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_398),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_442),
.B(n_450),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_461),
.B(n_366),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_454),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_456),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_446),
.B(n_366),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_366),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_469),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_508),
.B(n_459),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_498),
.B(n_461),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_462),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_468),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_485),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

AO22x2_ASAP7_75t_L g563 ( 
.A1(n_528),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_531),
.B(n_399),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_494),
.B(n_401),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_479),
.B(n_346),
.Y(n_567)
);

AND3x4_ASAP7_75t_L g568 ( 
.A(n_527),
.B(n_4),
.C(n_5),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_496),
.B(n_7),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_503),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_35),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_484),
.B(n_36),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_518),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_480),
.B(n_346),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_480),
.B(n_346),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_487),
.B(n_476),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_512),
.B(n_9),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_548),
.B(n_346),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_41),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_478),
.B(n_43),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_474),
.B(n_45),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_9),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_489),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_500),
.B(n_10),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_516),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_490),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_488),
.Y(n_595)
);

BUFx8_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_534),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_546),
.B(n_47),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_521),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_529),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_506),
.B(n_11),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_491),
.B(n_48),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_533),
.Y(n_603)
);

AO22x2_ASAP7_75t_L g604 ( 
.A1(n_544),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_519),
.B(n_12),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_513),
.B(n_14),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_541),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

AO22x2_ASAP7_75t_L g611 ( 
.A1(n_545),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_510),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_532),
.A2(n_129),
.B1(n_219),
.B2(n_218),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_504),
.B(n_18),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_517),
.B(n_49),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_530),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_489),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_560),
.A2(n_550),
.B1(n_551),
.B2(n_493),
.Y(n_621)
);

BUFx2_ASAP7_75t_SL g622 ( 
.A(n_579),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_586),
.A2(n_491),
.B(n_552),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_601),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_557),
.B(n_492),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_564),
.A2(n_491),
.B(n_552),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_564),
.A2(n_552),
.B(n_501),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_593),
.B(n_514),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_593),
.A2(n_501),
.B(n_489),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_555),
.A2(n_515),
.B(n_501),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_589),
.A2(n_553),
.B(n_539),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_554),
.B(n_509),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_592),
.B(n_502),
.C(n_481),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_558),
.A2(n_515),
.B(n_543),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_594),
.B(n_540),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_590),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_574),
.A2(n_515),
.B(n_612),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_579),
.B(n_517),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_574),
.A2(n_523),
.B(n_497),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_591),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_619),
.A2(n_523),
.B(n_497),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_617),
.A2(n_537),
.B(n_495),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_569),
.B(n_526),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_617),
.A2(n_542),
.B(n_530),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_583),
.B(n_492),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_572),
.B(n_526),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_578),
.B(n_536),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_609),
.A2(n_525),
.B1(n_472),
.B2(n_530),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_583),
.B(n_472),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_595),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_597),
.B(n_525),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_566),
.B(n_532),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_618),
.A2(n_128),
.B1(n_217),
.B2(n_214),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_571),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_571),
.Y(n_658)
);

NOR2x1_ASAP7_75t_L g659 ( 
.A(n_570),
.B(n_51),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_598),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_565),
.A2(n_126),
.B(n_213),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_565),
.A2(n_125),
.B(n_212),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_559),
.A2(n_124),
.B(n_208),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_573),
.Y(n_664)
);

AOI21x1_ASAP7_75t_L g665 ( 
.A1(n_606),
.A2(n_132),
.B(n_207),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_605),
.B(n_20),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_598),
.B(n_52),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_559),
.A2(n_133),
.B(n_206),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_573),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_561),
.A2(n_123),
.B(n_205),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_615),
.A2(n_122),
.B1(n_204),
.B2(n_203),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_561),
.A2(n_119),
.B(n_202),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_575),
.B(n_22),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_620),
.A2(n_588),
.B(n_607),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_575),
.Y(n_676)
);

NOR2x1p5_ASAP7_75t_SL g677 ( 
.A(n_608),
.B(n_55),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_588),
.A2(n_121),
.B(n_200),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_610),
.A2(n_116),
.B(n_199),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_57),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_587),
.B(n_22),
.C(n_23),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_576),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_587),
.A2(n_134),
.B1(n_197),
.B2(n_195),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_616),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_576),
.B(n_23),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_596),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_624),
.B(n_577),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_632),
.A2(n_613),
.B(n_614),
.C(n_577),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_625),
.B(n_596),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_633),
.B(n_581),
.C(n_580),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_660),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_657),
.B(n_580),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_631),
.A2(n_556),
.B(n_602),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_681),
.A2(n_603),
.B(n_600),
.C(n_556),
.Y(n_694)
);

OAI22x1_ASAP7_75t_L g695 ( 
.A1(n_682),
.A2(n_568),
.B1(n_611),
.B2(n_604),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_628),
.B(n_599),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_666),
.B(n_604),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_635),
.B(n_585),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_664),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_623),
.A2(n_582),
.B(n_567),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_674),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_675),
.A2(n_643),
.B(n_634),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_636),
.B(n_563),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_563),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_645),
.A2(n_611),
.B(n_115),
.Y(n_705)
);

INVx6_ASAP7_75t_L g706 ( 
.A(n_684),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_621),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_667),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_637),
.A2(n_138),
.B(n_192),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_674),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_658),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_648),
.B(n_30),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_669),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_655),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_684),
.B(n_31),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_676),
.A2(n_32),
.B1(n_60),
.B2(n_61),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_639),
.Y(n_717)
);

OAI21xp33_ASAP7_75t_SL g718 ( 
.A1(n_673),
.A2(n_63),
.B(n_64),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_651),
.B(n_65),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_685),
.B(n_66),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_644),
.B(n_67),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_641),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_684),
.B(n_68),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_650),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_647),
.B(n_69),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_674),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_653),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_649),
.B(n_70),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_646),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_654),
.B(n_71),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_653),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_640),
.B(n_642),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_652),
.B(n_72),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_638),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_641),
.B(n_73),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_680),
.B(n_630),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_627),
.A2(n_74),
.B(n_75),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_638),
.Y(n_739)
);

BUFx4f_ASAP7_75t_L g740 ( 
.A(n_680),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_622),
.B(n_78),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_629),
.A2(n_79),
.B(n_80),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_641),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_659),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_626),
.A2(n_81),
.B(n_82),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_683),
.B(n_83),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_680),
.B(n_220),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_677),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_678),
.B(n_84),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_743),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_706),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

BUFx4_ASAP7_75t_SL g753 ( 
.A(n_732),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_692),
.Y(n_754)
);

BUFx5_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_687),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_743),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_722),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_740),
.B(n_680),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

BUFx2_ASAP7_75t_SL g762 ( 
.A(n_701),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_735),
.B(n_661),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_710),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_710),
.Y(n_765)
);

CKINVDCx8_ASAP7_75t_R g766 ( 
.A(n_710),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_740),
.Y(n_767)
);

BUFx2_ASAP7_75t_SL g768 ( 
.A(n_727),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_727),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_691),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_699),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

BUFx4f_ASAP7_75t_L g774 ( 
.A(n_747),
.Y(n_774)
);

INVx11_ASAP7_75t_L g775 ( 
.A(n_706),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_723),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_735),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_739),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_713),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_714),
.A2(n_671),
.B1(n_672),
.B2(n_668),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_730),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_739),
.Y(n_782)
);

BUFx12f_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_696),
.B(n_663),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_747),
.Y(n_785)
);

BUFx4f_ASAP7_75t_SL g786 ( 
.A(n_689),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_728),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_717),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_698),
.B(n_665),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_724),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_729),
.B(n_670),
.Y(n_791)
);

BUFx12f_ASAP7_75t_L g792 ( 
.A(n_741),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_744),
.Y(n_793)
);

BUFx12f_ASAP7_75t_L g794 ( 
.A(n_697),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_736),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_703),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_746),
.B(n_662),
.Y(n_797)
);

BUFx12f_ASAP7_75t_L g798 ( 
.A(n_712),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_704),
.B(n_679),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_734),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_733),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_737),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_720),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_726),
.B(n_89),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_721),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_695),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_688),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_714),
.B(n_90),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_715),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_719),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_718),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_690),
.B(n_91),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_731),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_705),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_749),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_693),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_809),
.B(n_806),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_772),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_783),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_794),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_791),
.A2(n_702),
.B(n_742),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_809),
.B(n_707),
.C(n_708),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_796),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_791),
.A2(n_709),
.B(n_745),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_818),
.A2(n_700),
.B(n_738),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_779),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_775),
.Y(n_829)
);

XOR2xp5_ASAP7_75t_L g830 ( 
.A(n_806),
.B(n_92),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_801),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_769),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_756),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_797),
.A2(n_803),
.B(n_789),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_800),
.B(n_718),
.Y(n_836)
);

OAI211xp5_ASAP7_75t_SL g837 ( 
.A1(n_771),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_753),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_808),
.A2(n_817),
.B1(n_760),
.B2(n_774),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_803),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_756),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_771),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_755),
.Y(n_843)
);

AO31x2_ASAP7_75t_L g844 ( 
.A1(n_802),
.A2(n_99),
.A3(n_100),
.B(n_101),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_797),
.A2(n_103),
.B(n_104),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_817),
.A2(n_804),
.B(n_815),
.C(n_780),
.Y(n_846)
);

OA21x2_ASAP7_75t_L g847 ( 
.A1(n_818),
.A2(n_107),
.B(n_109),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_814),
.B(n_110),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_808),
.A2(n_114),
.B1(n_135),
.B2(n_136),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_754),
.B(n_140),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_SL g851 ( 
.A(n_795),
.B(n_141),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_808),
.A2(n_190),
.B1(n_143),
.B2(n_144),
.Y(n_852)
);

OA21x2_ASAP7_75t_L g853 ( 
.A1(n_815),
.A2(n_142),
.B(n_145),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_808),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_759),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_784),
.A2(n_149),
.B(n_150),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_753),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_754),
.B(n_151),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_780),
.A2(n_784),
.B(n_799),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_789),
.A2(n_153),
.B(n_154),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_755),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_816),
.B(n_155),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_814),
.B(n_157),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_793),
.A2(n_159),
.B(n_160),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_793),
.A2(n_161),
.B(n_162),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_811),
.B(n_163),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_781),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_750),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_816),
.B(n_164),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_787),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_781),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_798),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_787),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_755),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_792),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_778),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_767),
.A2(n_168),
.B(n_170),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_755),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_755),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_767),
.A2(n_171),
.B(n_172),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_750),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_778),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_867),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_836),
.A2(n_856),
.B(n_824),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_820),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_840),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_871),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_828),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_840),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_819),
.B(n_786),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_843),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_819),
.A2(n_774),
.B1(n_786),
.B2(n_807),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_861),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_831),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_823),
.A2(n_805),
.B(n_785),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_859),
.A2(n_813),
.B(n_763),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_874),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_842),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_831),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_878),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_879),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_825),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_856),
.A2(n_763),
.B(n_776),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_832),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_859),
.B(n_755),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_835),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_822),
.Y(n_907)
);

CKINVDCx6p67_ASAP7_75t_R g908 ( 
.A(n_821),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_834),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_825),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_833),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_853),
.B(n_812),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_841),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_842),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_862),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_868),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_844),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_846),
.B(n_790),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_870),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_827),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_881),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_826),
.A2(n_805),
.B(n_785),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_853),
.A2(n_812),
.B1(n_760),
.B2(n_811),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_844),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_857),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_855),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_873),
.B(n_812),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_844),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_876),
.B(n_812),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_882),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_915),
.A2(n_869),
.B1(n_862),
.B2(n_847),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_885),
.Y(n_933)
);

AO31x2_ASAP7_75t_L g934 ( 
.A1(n_917),
.A2(n_848),
.A3(n_863),
.B(n_866),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_885),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_888),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_898),
.B(n_875),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_892),
.B(n_837),
.C(n_839),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_902),
.B(n_846),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_888),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_894),
.B(n_838),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_926),
.B(n_766),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_902),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_904),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_R g945 ( 
.A(n_896),
.B(n_869),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_904),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_916),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_914),
.B(n_866),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_910),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_918),
.A2(n_837),
.B1(n_854),
.B2(n_872),
.C(n_850),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_908),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_915),
.A2(n_852),
.B1(n_849),
.B2(n_872),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_910),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_886),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_890),
.B(n_830),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_913),
.B(n_847),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_886),
.Y(n_957)
);

INVx8_ASAP7_75t_L g958 ( 
.A(n_915),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_899),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_907),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_889),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_889),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_915),
.A2(n_839),
.B(n_854),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_915),
.A2(n_852),
.B(n_862),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_891),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_899),
.B(n_848),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_905),
.B(n_863),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_906),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_958),
.Y(n_969)
);

OAI221xp5_ASAP7_75t_L g970 ( 
.A1(n_932),
.A2(n_884),
.B1(n_923),
.B2(n_907),
.C(n_849),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_960),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_SL g972 ( 
.A1(n_952),
.A2(n_915),
.B1(n_896),
.B2(n_912),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_952),
.A2(n_912),
.B(n_896),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_935),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_954),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_957),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_958),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_961),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_959),
.B(n_917),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_962),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_966),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_936),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_948),
.B(n_883),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_967),
.B(n_887),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_939),
.B(n_911),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_940),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_933),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_944),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_964),
.A2(n_884),
.B(n_963),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_943),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_973),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_986),
.B(n_982),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_990),
.A2(n_950),
.B(n_939),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_980),
.Y(n_995)
);

AO21x2_ASAP7_75t_L g996 ( 
.A1(n_974),
.A2(n_956),
.B(n_924),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_971),
.B(n_908),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_972),
.A2(n_938),
.B(n_903),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_973),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_983),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_969),
.A2(n_956),
.B(n_920),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_980),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_985),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_977),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_977),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_984),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_949),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_979),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_968),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_983),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_978),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1000),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1009),
.B(n_968),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_994),
.B(n_1006),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_997),
.B(n_971),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_993),
.B(n_978),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_995),
.B(n_991),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1007),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1002),
.B(n_975),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1004),
.Y(n_1020)
);

OAI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_998),
.A2(n_970),
.B1(n_945),
.B2(n_907),
.C(n_955),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1005),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1009),
.B(n_969),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1013),
.B(n_996),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1017),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1023),
.B(n_969),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_1011),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_1012),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1019),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1014),
.B(n_998),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1016),
.B(n_1013),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1014),
.B(n_996),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_1030),
.B(n_942),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1028),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1031),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1027),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1025),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1026),
.B(n_1015),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1039),
.B(n_1029),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_1032),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_1018),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1037),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1036),
.B(n_1020),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1036),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1038),
.B(n_1022),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1035),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1034),
.B(n_1024),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_1036),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1043),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1049),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_1015),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1045),
.B(n_1024),
.Y(n_1054)
);

INVxp67_ASAP7_75t_SL g1055 ( 
.A(n_1041),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1048),
.B(n_951),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1044),
.Y(n_1057)
);

AOI222xp33_ASAP7_75t_L g1058 ( 
.A1(n_1055),
.A2(n_1046),
.B1(n_1047),
.B2(n_1042),
.C1(n_1021),
.C2(n_937),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1053),
.B(n_925),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1051),
.Y(n_1060)
);

OAI32xp33_ASAP7_75t_L g1061 ( 
.A1(n_1054),
.A2(n_1012),
.A3(n_921),
.B1(n_996),
.B2(n_947),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_1056),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1055),
.A2(n_941),
.B1(n_968),
.B2(n_916),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1051),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1060),
.B(n_1064),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1062),
.B(n_1059),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1063),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1058),
.B(n_1057),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_1052),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_1066),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1065),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_1050),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1067),
.B(n_829),
.Y(n_1073)
);

OAI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1068),
.A2(n_851),
.B1(n_869),
.B2(n_916),
.C(n_992),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1065),
.B(n_1000),
.Y(n_1075)
);

AOI222xp33_ASAP7_75t_L g1076 ( 
.A1(n_1072),
.A2(n_810),
.B1(n_858),
.B2(n_1001),
.C1(n_999),
.C2(n_992),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1073),
.B(n_941),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_999),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1071),
.Y(n_1079)
);

OAI211xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1074),
.A2(n_751),
.B(n_1008),
.C(n_1010),
.Y(n_1080)
);

NAND4xp75_ASAP7_75t_L g1081 ( 
.A(n_1075),
.B(n_1008),
.C(n_1010),
.D(n_981),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_L g1082 ( 
.A(n_1079),
.B(n_757),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1081),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1078),
.A2(n_1001),
.B(n_752),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1077),
.B(n_987),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1080),
.Y(n_1086)
);

AOI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1086),
.A2(n_1076),
.B1(n_757),
.B2(n_976),
.C(n_981),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1082),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1083),
.B(n_987),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_1084),
.B(n_757),
.C(n_752),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1085),
.A2(n_880),
.B(n_877),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1086),
.B(n_761),
.C(n_764),
.Y(n_1092)
);

OAI31xp33_ASAP7_75t_L g1093 ( 
.A1(n_1086),
.A2(n_912),
.A3(n_770),
.B(n_765),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1086),
.A2(n_976),
.B1(n_765),
.B2(n_770),
.C(n_758),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1089),
.B(n_761),
.C(n_764),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1088),
.B(n_979),
.Y(n_1096)
);

XOR2x2_ASAP7_75t_L g1097 ( 
.A(n_1092),
.B(n_173),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1090),
.Y(n_1098)
);

NOR4xp25_ASAP7_75t_L g1099 ( 
.A(n_1094),
.B(n_953),
.C(n_988),
.D(n_989),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1087),
.A2(n_752),
.B1(n_810),
.B2(n_958),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1091),
.B(n_989),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_752),
.B1(n_988),
.B2(n_911),
.Y(n_1102)
);

AOI322xp5_ASAP7_75t_L g1103 ( 
.A1(n_1092),
.A2(n_924),
.A3(n_928),
.B1(n_929),
.B2(n_905),
.C1(n_894),
.C2(n_931),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1089),
.B(n_934),
.Y(n_1104)
);

AND2x2_ASAP7_75t_SL g1105 ( 
.A(n_1098),
.B(n_758),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1096),
.Y(n_1106)
);

AND4x1_ASAP7_75t_L g1107 ( 
.A(n_1095),
.B(n_175),
.C(n_178),
.D(n_179),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_1102),
.B(n_845),
.C(n_865),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1104),
.B(n_768),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1097),
.A2(n_773),
.B1(n_758),
.B2(n_762),
.Y(n_1110)
);

XNOR2x1_ASAP7_75t_L g1111 ( 
.A(n_1100),
.B(n_180),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1099),
.B(n_934),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1101),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1103),
.B(n_934),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_L g1115 ( 
.A1(n_1098),
.A2(n_773),
.B(n_860),
.C(n_864),
.Y(n_1115)
);

AOI322xp5_ASAP7_75t_L g1116 ( 
.A1(n_1098),
.A2(n_929),
.A3(n_928),
.B1(n_913),
.B2(n_930),
.C1(n_773),
.C2(n_919),
.Y(n_1116)
);

XOR2x1_ASAP7_75t_L g1117 ( 
.A(n_1113),
.B(n_181),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1105),
.B(n_777),
.Y(n_1118)
);

NOR2x1p5_ASAP7_75t_L g1119 ( 
.A(n_1106),
.B(n_782),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1109),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1110),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1107),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1111),
.Y(n_1123)
);

XNOR2xp5_ASAP7_75t_L g1124 ( 
.A(n_1112),
.B(n_1114),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_1117),
.Y(n_1125)
);

XNOR2xp5_ASAP7_75t_L g1126 ( 
.A(n_1122),
.B(n_1108),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1124),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1118),
.Y(n_1128)
);

XNOR2xp5_ASAP7_75t_L g1129 ( 
.A(n_1123),
.B(n_1115),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1120),
.Y(n_1130)
);

AOI22x1_ASAP7_75t_L g1131 ( 
.A1(n_1121),
.A2(n_1119),
.B1(n_1116),
.B2(n_778),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1130),
.Y(n_1132)
);

XNOR2x1_ASAP7_75t_SL g1133 ( 
.A(n_1126),
.B(n_182),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1127),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1135),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1136),
.A2(n_1125),
.B1(n_1134),
.B2(n_1128),
.Y(n_1137)
);

AO21x1_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1133),
.B(n_1129),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1137),
.A2(n_1131),
.B1(n_790),
.B2(n_903),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1137),
.A2(n_790),
.B1(n_782),
.B2(n_906),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1139),
.A2(n_816),
.B1(n_906),
.B2(n_187),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1138),
.Y(n_1142)
);

OAI222xp33_ASAP7_75t_L g1143 ( 
.A1(n_1140),
.A2(n_184),
.B1(n_185),
.B2(n_188),
.C1(n_891),
.C2(n_900),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1138),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_R g1145 ( 
.A1(n_1142),
.A2(n_946),
.B1(n_900),
.B2(n_893),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1144),
.A2(n_930),
.B1(n_901),
.B2(n_893),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1141),
.B(n_901),
.C(n_897),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1143),
.A2(n_897),
.B1(n_896),
.B2(n_909),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_909),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_1147),
.A2(n_922),
.B(n_927),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1145),
.B(n_922),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_895),
.Y(n_1152)
);

AOI211xp5_ASAP7_75t_L g1153 ( 
.A1(n_1152),
.A2(n_1151),
.B(n_1150),
.C(n_895),
.Y(n_1153)
);


endmodule