module fake_jpeg_30782_n_328 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_42),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_57),
.Y(n_63)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_70),
.B1(n_74),
.B2(n_89),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_79),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_27),
.B1(n_19),
.B2(n_36),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_38),
.B1(n_30),
.B2(n_33),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_83),
.B1(n_85),
.B2(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_75),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_20),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_19),
.B1(n_22),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_35),
.B1(n_23),
.B2(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_90),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_1),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_96),
.C(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_59),
.B1(n_58),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_41),
.B1(n_40),
.B2(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_40),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_27),
.B1(n_39),
.B2(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_44),
.A2(n_26),
.B1(n_21),
.B2(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_44),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_96),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_125),
.C(n_128),
.Y(n_166)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_35),
.B1(n_23),
.B2(n_19),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_114),
.A2(n_121),
.B1(n_123),
.B2(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_136),
.B1(n_140),
.B2(n_67),
.Y(n_154)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_1),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_102),
.C(n_65),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_131),
.Y(n_145)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_73),
.B(n_64),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_111),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_91),
.B(n_73),
.C(n_97),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_102),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_138),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_147),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_72),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_65),
.B(n_104),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_144),
.B(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_161),
.B1(n_129),
.B2(n_116),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_91),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_91),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_64),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_8),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_108),
.B(n_109),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_128),
.B(n_118),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_84),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_151),
.Y(n_185)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_182),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_180),
.B(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_127),
.B1(n_170),
.B2(n_169),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_184),
.B(n_194),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_107),
.B1(n_140),
.B2(n_121),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_195),
.B1(n_196),
.B2(n_204),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_107),
.B(n_121),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_145),
.B(n_152),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_125),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_199),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_121),
.B1(n_125),
.B2(n_67),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_69),
.B1(n_84),
.B2(n_80),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_159),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_110),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_110),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_152),
.Y(n_213)
);

AO21x1_ASAP7_75t_SL g202 ( 
.A1(n_143),
.A2(n_133),
.B(n_119),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_69),
.B1(n_80),
.B2(n_62),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_157),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_130),
.B1(n_62),
.B2(n_134),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_187),
.B1(n_181),
.B2(n_206),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_163),
.C(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_214),
.C(n_229),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_234),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_158),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_207),
.B(n_188),
.C(n_194),
.D(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_145),
.B(n_176),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_153),
.B(n_113),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_153),
.B(n_148),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_223),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_192),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_233),
.B1(n_176),
.B2(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_148),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_186),
.B1(n_195),
.B2(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_245),
.C(n_257),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_207),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_191),
.B1(n_202),
.B2(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_182),
.Y(n_245)
);

NAND5xp2_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_201),
.C(n_199),
.D(n_177),
.E(n_208),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_249),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_235),
.B(n_218),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_164),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_227),
.C(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_164),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_205),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_209),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_264),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_261),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_221),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_273),
.C(n_239),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_228),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_250),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_223),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_239),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_244),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_216),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_236),
.B(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_287),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_284),
.C(n_273),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_252),
.B1(n_220),
.B2(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_236),
.B(n_242),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_274),
.B1(n_237),
.B2(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_285),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_254),
.B1(n_248),
.B2(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_255),
.C(n_253),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_297),
.C(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_296),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_267),
.B(n_238),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_205),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_261),
.C(n_262),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_298),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_212),
.Y(n_298)
);

XOR2x2_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_308),
.Y(n_313)
);

AOI31xp33_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_288),
.A3(n_277),
.B(n_280),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_307),
.B(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_289),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_278),
.B(n_212),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_295),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_308),
.CI(n_307),
.CON(n_320),
.SN(n_320)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_315),
.A3(n_295),
.B1(n_12),
.B2(n_15),
.C1(n_11),
.C2(n_8),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_324),
.B(n_317),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_11),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_323),
.Y(n_328)
);


endmodule