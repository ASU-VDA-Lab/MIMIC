module real_jpeg_6957_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_78),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_78),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_1),
.A2(n_78),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_2),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_73),
.B1(n_141),
.B2(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_73),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_3),
.A2(n_73),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_5),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_5),
.Y(n_185)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_5),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_5),
.Y(n_393)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_8),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_10),
.Y(n_435)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_52),
.B1(n_106),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_52),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_12),
.B(n_66),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_12),
.A2(n_336),
.B(n_339),
.C(n_343),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_12),
.B(n_91),
.C(n_274),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_12),
.B(n_22),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_12),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_12),
.B(n_96),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_230),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_13),
.A2(n_230),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_13),
.A2(n_100),
.B1(n_230),
.B2(n_369),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_430),
.B(n_432),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_152),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_18),
.B(n_124),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_55),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_20),
.A2(n_21),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_20),
.B(n_305),
.C(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B(n_49),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_22),
.B(n_114),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_22),
.A2(n_112),
.B(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_22),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_27),
.Y(n_338)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_31),
.Y(n_352)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_34),
.Y(n_171)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_34),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_34),
.Y(n_351)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_37),
.A2(n_140),
.B(n_148),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_37),
.B(n_49),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_37),
.B(n_249),
.Y(n_277)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_38),
.B(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_42),
.Y(n_144)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_48),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_49),
.Y(n_119)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_50),
.Y(n_343)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_51),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_52),
.A2(n_76),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_52),
.B(n_135),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_52),
.A2(n_340),
.B(n_341),
.Y(n_339)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_70),
.B(n_74),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_56),
.A2(n_122),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_57),
.B(n_228),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g264 ( 
.A(n_62),
.B(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_65),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_66),
.B(n_133),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_66),
.B(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_74),
.B(n_227),
.Y(n_296)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_111),
.C(n_120),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_82),
.A2(n_111),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_82),
.B(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_82),
.A2(n_130),
.B1(n_246),
.B2(n_254),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_82),
.B(n_243),
.C(n_246),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_103),
.B(n_104),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_83),
.A2(n_190),
.B(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_84),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_84),
.B(n_105),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_84),
.B(n_348),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_96),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_91),
.B2(n_94),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_87),
.Y(n_342)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_96),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_96),
.B(n_348),
.Y(n_363)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_96)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_98),
.Y(n_221)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_98),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_100),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_101),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_103),
.B(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_103),
.A2(n_168),
.B(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_112),
.Y(n_247)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_115),
.Y(n_253)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_118),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_123),
.B(n_244),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.C(n_138),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_131),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_132),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_134),
.Y(n_263)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_138),
.B(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_144),
.Y(n_259)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_149),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_149),
.B(n_277),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_236),
.B(n_426),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_232),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_199),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_156),
.B(n_199),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_175),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_159),
.B(n_163),
.C(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_165),
.B(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_174),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_166),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_168),
.B(n_363),
.Y(n_406)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_171),
.Y(n_360)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_196),
.B(n_197),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_177),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_196),
.B1(n_197),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_178),
.A2(n_189),
.B1(n_196),
.B2(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_178),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_178),
.A2(n_196),
.B1(n_335),
.B2(n_409),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_186),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_179),
.B(n_186),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_179),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_179),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_180),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_181),
.Y(n_372)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_189),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_195),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_195),
.B(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.C(n_206),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_206),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_223),
.C(n_225),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_207),
.A2(n_208),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_209),
.B(n_222),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_210),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_211),
.A2(n_217),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_216),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_223),
.B(n_225),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_224),
.B(n_248),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_232),
.A2(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_233),
.B(n_235),
.Y(n_429)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_418),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_310),
.C(n_325),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_299),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_285),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_241),
.B(n_285),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_255),
.C(n_275),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_242),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_255),
.A2(n_256),
.B1(n_275),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_268),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_257),
.B(n_268),
.Y(n_294)
);

AOI32xp33_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.A3(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_282),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.C(n_280),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_280),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_281),
.B(n_384),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_282),
.B(n_367),
.Y(n_396)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_288),
.C(n_293),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_292),
.B(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_299),
.A2(n_421),
.B(n_422),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_300),
.B(n_309),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_322),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_311),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_312),
.B(n_319),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_316),
.CI(n_318),
.CON(n_323),
.SN(n_323)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_323),
.B(n_324),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g437 ( 
.A(n_323),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_353),
.B(n_417),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_327),
.B(n_330),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.C(n_344),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_331),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_334),
.A2(n_344),
.B1(n_345),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_336),
.Y(n_340)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx11_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_411),
.B(n_416),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_401),
.B(n_410),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_378),
.B(n_400),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_364),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_364),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_381),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_373),
.Y(n_364)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_385),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_376),
.C(n_403),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_387),
.B(n_399),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_382),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_395),
.B(n_398),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_396),
.B(n_397),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_404),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_407),
.C(n_408),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_415),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_420),
.B(n_423),
.C(n_424),
.D(n_425),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx13_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);


endmodule