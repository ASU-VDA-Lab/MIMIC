module fake_jpeg_864_n_678 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_678);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_678;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_487;
wire n_193;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_60),
.B(n_62),
.Y(n_146)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_63),
.B(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_68),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_79),
.B(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_83),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_91),
.Y(n_169)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g204 ( 
.A(n_98),
.Y(n_204)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_113),
.Y(n_189)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_104),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_118),
.Y(n_135)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_27),
.B(n_8),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_31),
.B(n_8),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_50),
.Y(n_134)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_49),
.B(n_11),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_134),
.B(n_25),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_139),
.A2(n_153),
.B1(n_36),
.B2(n_52),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_56),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_141),
.B(n_175),
.Y(n_249)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_36),
.B1(n_34),
.B2(n_52),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_108),
.B(n_19),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_162),
.B(n_194),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_59),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_56),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_59),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_183),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_25),
.C(n_58),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_178),
.B(n_46),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_55),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_74),
.B(n_21),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_76),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_64),
.A2(n_23),
.B1(n_53),
.B2(n_46),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_199),
.A2(n_37),
.B1(n_30),
.B2(n_23),
.Y(n_283)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_112),
.B(n_55),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_208),
.B(n_39),
.Y(n_271)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_83),
.B(n_34),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_214),
.B(n_37),
.Y(n_282)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_77),
.Y(n_217)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_81),
.B(n_22),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_219),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_82),
.B(n_58),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g322 ( 
.A(n_224),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_68),
.B1(n_110),
.B2(n_103),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_226),
.A2(n_260),
.B1(n_283),
.B2(n_286),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_164),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_228),
.A2(n_229),
.B(n_237),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_124),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_232),
.A2(n_302),
.B1(n_158),
.B2(n_179),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_146),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_234),
.B(n_239),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_154),
.B(n_70),
.C(n_97),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_238),
.B(n_244),
.C(n_166),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_30),
.B(n_19),
.C(n_53),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_241),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_167),
.B(n_25),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_242),
.B(n_248),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_243),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_161),
.B(n_80),
.C(n_96),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_245),
.Y(n_319)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_131),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_146),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_148),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_252),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_167),
.B(n_25),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_253),
.B(n_263),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

CKINVDCx9p33_ASAP7_75t_R g257 ( 
.A(n_204),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_257),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_169),
.A2(n_84),
.B1(n_95),
.B2(n_73),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_261),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_169),
.B(n_25),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_155),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_267),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_52),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_171),
.B(n_98),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_270),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_138),
.B(n_39),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_271),
.B(n_279),
.Y(n_350)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_272),
.Y(n_361)
);

CKINVDCx12_ASAP7_75t_R g273 ( 
.A(n_219),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_273),
.Y(n_363)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_172),
.Y(n_274)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_155),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_280),
.Y(n_315)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_214),
.Y(n_277)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_180),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_165),
.Y(n_281)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_287),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_139),
.A2(n_33),
.B(n_57),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_298),
.Y(n_312)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_144),
.Y(n_285)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_221),
.A2(n_85),
.B1(n_72),
.B2(n_71),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_135),
.A2(n_33),
.B(n_57),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_144),
.Y(n_288)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_180),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_291),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_201),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_137),
.Y(n_294)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_147),
.Y(n_295)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_190),
.A2(n_57),
.B1(n_26),
.B2(n_0),
.Y(n_296)
);

AO22x1_ASAP7_75t_SL g331 ( 
.A1(n_296),
.A2(n_212),
.B1(n_202),
.B2(n_196),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_145),
.B(n_13),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_170),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_166),
.Y(n_300)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_153),
.A2(n_222),
.B1(n_157),
.B2(n_156),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_143),
.Y(n_303)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_304),
.B(n_331),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_140),
.C(n_136),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_307),
.B(n_309),
.C(n_292),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_163),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_260),
.A2(n_187),
.B1(n_184),
.B2(n_200),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_311),
.A2(n_327),
.B1(n_329),
.B2(n_336),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_228),
.A2(n_212),
.B1(n_202),
.B2(n_200),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_258),
.A2(n_279),
.B1(n_228),
.B2(n_229),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_235),
.B(n_142),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_338),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_258),
.A2(n_196),
.B1(n_192),
.B2(n_174),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_181),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_229),
.A2(n_160),
.B1(n_192),
.B2(n_174),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_341),
.A2(n_355),
.B1(n_247),
.B2(n_296),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_231),
.Y(n_347)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_231),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_352),
.Y(n_403)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_233),
.Y(n_353)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_233),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_354),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_267),
.A2(n_236),
.B1(n_284),
.B2(n_286),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_257),
.Y(n_356)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_240),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_364),
.B(n_300),
.Y(n_410)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_365),
.A2(n_386),
.B1(n_398),
.B2(n_401),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_377),
.Y(n_415)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_312),
.A2(n_232),
.B1(n_226),
.B2(n_160),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_371),
.A2(n_406),
.B1(n_311),
.B2(n_339),
.Y(n_427)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_359),
.B(n_239),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_374),
.B(n_393),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_238),
.B(n_244),
.C(n_232),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_375),
.B(n_382),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_225),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_376),
.B(n_378),
.C(n_395),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_315),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_360),
.C(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_304),
.B(n_250),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_380),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_255),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_338),
.B(n_264),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_381),
.B(n_399),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_240),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_151),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_384),
.B(n_392),
.Y(n_452)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_318),
.A2(n_281),
.B1(n_289),
.B2(n_262),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_387),
.A2(n_390),
.B1(n_326),
.B2(n_347),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_345),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_396),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_337),
.A2(n_256),
.B1(n_262),
.B2(n_274),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_407),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_310),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_308),
.B(n_256),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_266),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_243),
.C(n_252),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_345),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_328),
.A2(n_247),
.B1(n_230),
.B2(n_241),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_313),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_404),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_335),
.A2(n_241),
.B1(n_251),
.B2(n_293),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_293),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_305),
.B(n_259),
.Y(n_404)
);

FAx1_ASAP7_75t_SL g405 ( 
.A(n_327),
.B(n_205),
.CI(n_275),
.CON(n_405),
.SN(n_405)
);

OAI32xp33_ASAP7_75t_L g421 ( 
.A1(n_405),
.A2(n_317),
.A3(n_326),
.B1(n_332),
.B2(n_331),
.Y(n_421)
);

OAI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_335),
.A2(n_295),
.B1(n_288),
.B2(n_254),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_305),
.B(n_301),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_320),
.B(n_259),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_408),
.Y(n_449)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_320),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_364),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_335),
.B(n_342),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_416),
.A2(n_424),
.B(n_444),
.Y(n_467)
);

O2A1O1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_411),
.A2(n_331),
.B(n_358),
.C(n_317),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_417),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_421),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_423),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_324),
.B(n_316),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_432),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_368),
.B(n_371),
.Y(n_432)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_340),
.B1(n_339),
.B2(n_361),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_438),
.B1(n_439),
.B2(n_447),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_388),
.A2(n_306),
.B1(n_339),
.B2(n_332),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_368),
.A2(n_340),
.B1(n_361),
.B2(n_321),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_399),
.A2(n_321),
.B1(n_351),
.B2(n_357),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_367),
.A2(n_246),
.B1(n_272),
.B2(n_261),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_442),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_367),
.A2(n_379),
.B1(n_372),
.B2(n_382),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_389),
.A2(n_316),
.B(n_306),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_396),
.A2(n_332),
.B1(n_344),
.B2(n_357),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_446),
.A2(n_362),
.B(n_322),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_372),
.A2(n_351),
.B1(n_342),
.B2(n_314),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g450 ( 
.A1(n_374),
.A2(n_393),
.A3(n_378),
.B1(n_405),
.B2(n_392),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_376),
.Y(n_462)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_453),
.Y(n_498)
);

AO22x1_ASAP7_75t_SL g454 ( 
.A1(n_432),
.A2(n_384),
.B1(n_405),
.B2(n_403),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_454),
.B(n_460),
.Y(n_515)
);

INVx13_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_458),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_424),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_462),
.B(n_465),
.Y(n_503)
);

CKINVDCx10_ASAP7_75t_R g463 ( 
.A(n_444),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_463),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_415),
.B(n_366),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_437),
.B(n_377),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_468),
.B(n_481),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_412),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_469),
.B(n_485),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_391),
.Y(n_472)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_474),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_415),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_475),
.A2(n_489),
.B1(n_416),
.B2(n_428),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_381),
.Y(n_478)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_385),
.B(n_409),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_479),
.A2(n_487),
.B(n_451),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_395),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_480),
.B(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_426),
.B(n_381),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_421),
.B(n_434),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_482),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_432),
.A2(n_400),
.B1(n_403),
.B2(n_410),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_483),
.A2(n_417),
.B1(n_445),
.B2(n_433),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_403),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_448),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_397),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_383),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_486),
.B(n_488),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_423),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_423),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_431),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_490),
.B(n_507),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_492),
.B(n_490),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_437),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_493),
.B(n_495),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_431),
.C(n_443),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_494),
.B(n_496),
.C(n_497),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_414),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_432),
.C(n_414),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_438),
.C(n_425),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_430),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_499),
.B(n_502),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_501),
.A2(n_518),
.B(n_467),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_452),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_457),
.A2(n_464),
.B1(n_482),
.B2(n_459),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_504),
.A2(n_524),
.B1(n_489),
.B2(n_488),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_459),
.A2(n_457),
.B1(n_478),
.B2(n_456),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_505),
.A2(n_508),
.B1(n_514),
.B2(n_520),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_425),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_457),
.A2(n_425),
.B1(n_427),
.B2(n_439),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_474),
.B(n_428),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_526),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_486),
.Y(n_513)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_513),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_456),
.A2(n_441),
.B1(n_447),
.B2(n_417),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_484),
.B(n_409),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_516),
.Y(n_537)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_520),
.A2(n_477),
.B1(n_467),
.B2(n_463),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_522),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_482),
.A2(n_450),
.B1(n_418),
.B2(n_413),
.Y(n_524)
);

AO22x1_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_422),
.B1(n_419),
.B2(n_369),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_527),
.A2(n_530),
.B1(n_542),
.B2(n_543),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_528),
.B(n_534),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_455),
.B1(n_461),
.B2(n_471),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_461),
.Y(n_532)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_500),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_454),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_546),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_522),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_547),
.Y(n_567)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_538),
.B(n_548),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_541),
.A2(n_554),
.B(n_558),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_525),
.A2(n_477),
.B1(n_460),
.B2(n_454),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_454),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_466),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_525),
.A2(n_458),
.B1(n_455),
.B2(n_473),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_498),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_549),
.A2(n_550),
.B1(n_552),
.B2(n_555),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_498),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_513),
.B(n_512),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_551),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_505),
.A2(n_473),
.B1(n_470),
.B2(n_466),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_492),
.B(n_470),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_553),
.B(n_507),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_506),
.A2(n_487),
.B(n_458),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_503),
.A2(n_453),
.B1(n_422),
.B2(n_419),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_512),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_557),
.B(n_521),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_518),
.A2(n_344),
.B(n_386),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_506),
.A2(n_453),
.B1(n_373),
.B2(n_314),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_559),
.A2(n_498),
.B1(n_491),
.B2(n_509),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_573),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_497),
.C(n_491),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_561),
.B(n_571),
.C(n_574),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_SL g599 ( 
.A1(n_562),
.A2(n_579),
.B1(n_538),
.B2(n_559),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_529),
.B(n_516),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_575),
.Y(n_588)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_568),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_556),
.B(n_515),
.C(n_523),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_530),
.A2(n_515),
.B1(n_521),
.B2(n_511),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_572),
.A2(n_580),
.B1(n_365),
.B2(n_227),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_524),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_533),
.B(n_504),
.C(n_514),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_533),
.B(n_526),
.C(n_322),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_528),
.C(n_546),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_576),
.B(n_577),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_535),
.B(n_543),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_547),
.Y(n_578)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_526),
.C(n_509),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_584),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_527),
.A2(n_285),
.B1(n_354),
.B2(n_353),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_531),
.A2(n_352),
.B(n_362),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_583),
.A2(n_558),
.B(n_532),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_386),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_567),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_589),
.B(n_591),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_590),
.A2(n_596),
.B(n_566),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_584),
.B(n_548),
.Y(n_591)
);

AOI321xp33_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_554),
.A3(n_536),
.B1(n_539),
.B2(n_544),
.C(n_540),
.Y(n_592)
);

OAI22x1_ASAP7_75t_L g620 ( 
.A1(n_592),
.A2(n_560),
.B1(n_580),
.B2(n_275),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_586),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_593),
.B(n_188),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_569),
.A2(n_531),
.B1(n_544),
.B2(n_540),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_594),
.A2(n_601),
.B1(n_605),
.B2(n_606),
.Y(n_615)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_585),
.A2(n_545),
.B(n_539),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_561),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_599),
.A2(n_608),
.B1(n_562),
.B2(n_573),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_569),
.A2(n_552),
.B1(n_557),
.B2(n_550),
.Y(n_601)
);

NOR4xp25_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_549),
.C(n_334),
.D(n_227),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_13),
.C(n_2),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_563),
.A2(n_159),
.B1(n_334),
.B2(n_224),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_581),
.A2(n_159),
.B1(n_365),
.B2(n_251),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_563),
.A2(n_572),
.B(n_577),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_607),
.A2(n_206),
.B(n_186),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_152),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_609),
.B(n_575),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_611),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_574),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_612),
.B(n_613),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_566),
.C(n_576),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_587),
.C(n_604),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_614),
.B(n_620),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_604),
.B(n_564),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_616),
.B(n_617),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_618),
.A2(n_592),
.B(n_591),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_564),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_619),
.B(n_622),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_587),
.B(n_191),
.C(n_193),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_624),
.C(n_628),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_206),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_623),
.B(n_12),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_591),
.B(n_149),
.C(n_150),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_625),
.A2(n_626),
.B(n_590),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_601),
.B(n_57),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_615),
.A2(n_589),
.B1(n_600),
.B2(n_603),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_631),
.B(n_632),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_627),
.A2(n_600),
.B1(n_603),
.B2(n_597),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_633),
.B(n_636),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_634),
.A2(n_12),
.B(n_2),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_594),
.C(n_608),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_613),
.B(n_605),
.C(n_609),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_637),
.B(n_638),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_618),
.B(n_57),
.C(n_1),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_641),
.B(n_15),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_1),
.C(n_26),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_643),
.B(n_644),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_1),
.C(n_26),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_648),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_640),
.B(n_637),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_651),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_639),
.B(n_622),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_636),
.B(n_628),
.C(n_620),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_624),
.C(n_621),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_652),
.B(n_655),
.Y(n_664)
);

AOI31xp67_ASAP7_75t_L g658 ( 
.A1(n_653),
.A2(n_638),
.A3(n_644),
.B(n_635),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_629),
.B(n_13),
.Y(n_654)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_654),
.Y(n_663)
);

AOI32xp33_ASAP7_75t_L g655 ( 
.A1(n_634),
.A2(n_26),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_L g657 ( 
.A1(n_646),
.A2(n_630),
.B(n_642),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_657),
.B(n_658),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_649),
.B(n_635),
.C(n_643),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_647),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_650),
.A2(n_7),
.B(n_3),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_660),
.A2(n_656),
.B(n_3),
.Y(n_666)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_666),
.Y(n_672)
);

AOI322xp5_ASAP7_75t_L g671 ( 
.A1(n_667),
.A2(n_668),
.A3(n_669),
.B1(n_664),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_661),
.B(n_652),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_662),
.B(n_651),
.Y(n_669)
);

A2O1A1O1Ixp25_ASAP7_75t_L g670 ( 
.A1(n_665),
.A2(n_664),
.B(n_663),
.C(n_6),
.D(n_7),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_670),
.A2(n_14),
.B(n_16),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_671),
.A2(n_5),
.B(n_14),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_673),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_675),
.B(n_672),
.C(n_674),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_17),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_677),
.B(n_1),
.Y(n_678)
);


endmodule