module fake_jpeg_4645_n_243 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_1),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_18),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_53),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_59),
.B(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_27),
.B1(n_28),
.B2(n_17),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_80),
.B1(n_28),
.B2(n_22),
.Y(n_106)
);

NOR2x1_ASAP7_75t_R g71 ( 
.A(n_37),
.B(n_27),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_83),
.B1(n_85),
.B2(n_59),
.Y(n_96)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_86),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_39),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_4),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_78),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_3),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_115),
.C(n_4),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_28),
.B1(n_33),
.B2(n_45),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_30),
.B1(n_29),
.B2(n_41),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_117),
.B1(n_86),
.B2(n_79),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_53),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_74),
.B1(n_57),
.B2(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_61),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_118),
.A2(n_139),
.B1(n_142),
.B2(n_104),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_56),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_87),
.B(n_68),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_146),
.B(n_91),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_136),
.B1(n_91),
.B2(n_97),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_50),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_109),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_130),
.CI(n_140),
.CON(n_166),
.SN(n_166)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_75),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_93),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_68),
.B1(n_88),
.B2(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_4),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_67),
.B1(n_51),
.B2(n_25),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_5),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_25),
.C(n_16),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_5),
.B(n_6),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_163),
.B1(n_118),
.B2(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_165),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_158),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_159),
.B(n_160),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_99),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_120),
.B(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_104),
.B1(n_94),
.B2(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_100),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_166),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_128),
.C(n_121),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_178),
.C(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_145),
.C(n_138),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_149),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_122),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_150),
.B(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_156),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_134),
.A3(n_137),
.B1(n_141),
.B2(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_189),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_146),
.B(n_135),
.Y(n_186)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_131),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_158),
.B1(n_150),
.B2(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_198),
.B1(n_199),
.B2(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_200),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_170),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_152),
.B(n_164),
.C(n_157),
.D(n_154),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_208),
.Y(n_221)
);

OAI321xp33_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_183),
.A3(n_185),
.B1(n_177),
.B2(n_178),
.C(n_188),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_197),
.B1(n_204),
.B2(n_182),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_179),
.C(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_214),
.C(n_190),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_152),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_152),
.B1(n_184),
.B2(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_200),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_175),
.B1(n_149),
.B2(n_105),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_219),
.B1(n_215),
.B2(n_206),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_201),
.B(n_190),
.C(n_10),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_98),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_223),
.C(n_107),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_175),
.C(n_153),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_229),
.Y(n_231)
);

OAI31xp33_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_213),
.A3(n_205),
.B(n_211),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_230),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_9),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_228),
.B(n_6),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_94),
.C(n_13),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_234),
.B(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_13),
.C(n_10),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_11),
.B1(n_176),
.B2(n_182),
.Y(n_242)
);

NAND2x1p5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_240),
.Y(n_243)
);


endmodule