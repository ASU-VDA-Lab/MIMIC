module fake_jpeg_157_n_584 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_584);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_54),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_59),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_63),
.B(n_74),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_1),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_103),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_1),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_3),
.Y(n_113)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_96),
.Y(n_131)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_2),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

BUFx2_ASAP7_75t_R g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_106),
.Y(n_150)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_53),
.B(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_2),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_30),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_113),
.B(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_118),
.B(n_127),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_93),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_51),
.B1(n_47),
.B2(n_50),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_121),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_52),
.B1(n_35),
.B2(n_51),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_126),
.A2(n_140),
.B1(n_157),
.B2(n_22),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_39),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_34),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_56),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_144),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_54),
.A2(n_35),
.B1(n_47),
.B2(n_51),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_97),
.B(n_25),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_57),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_25),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_78),
.B(n_34),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_98),
.A2(n_47),
.B1(n_22),
.B2(n_29),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_50),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_163),
.B(n_36),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_60),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_48),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_175),
.Y(n_281)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_52),
.B1(n_33),
.B2(n_48),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_180),
.A2(n_205),
.B1(n_234),
.B2(n_110),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_94),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_189),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_187),
.Y(n_278)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_41),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_115),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_190),
.B(n_208),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_108),
.B1(n_62),
.B2(n_106),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_193),
.B1(n_199),
.B2(n_203),
.Y(n_251)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_192),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_64),
.B1(n_101),
.B2(n_100),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_121),
.A2(n_68),
.B1(n_107),
.B2(n_44),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_SL g253 ( 
.A1(n_195),
.A2(n_211),
.B(n_236),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_197),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_140),
.A2(n_80),
.B1(n_95),
.B2(n_90),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_79),
.B1(n_86),
.B2(n_85),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_23),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_207),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_81),
.B1(n_69),
.B2(n_102),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_213),
.Y(n_243)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_44),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_210),
.Y(n_255)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_40),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_223),
.C(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_215),
.B(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_44),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_216),
.B(n_226),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_218),
.Y(n_257)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_225),
.B1(n_129),
.B2(n_161),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_222),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_125),
.B(n_73),
.Y(n_221)
);

NAND2x1_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_166),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_41),
.C(n_40),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_32),
.B1(n_29),
.B2(n_38),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_29),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_136),
.B(n_3),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_136),
.B(n_38),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_3),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_38),
.C(n_31),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_232),
.B(n_117),
.CI(n_31),
.CON(n_290),
.SN(n_290)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_233),
.A2(n_117),
.B1(n_5),
.B2(n_7),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_133),
.A2(n_38),
.B1(n_31),
.B2(n_7),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_159),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_122),
.A2(n_38),
.B1(n_31),
.B2(n_7),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_142),
.B1(n_130),
.B2(n_123),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_242),
.A2(n_261),
.B1(n_272),
.B2(n_282),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_147),
.B(n_122),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_244),
.A2(n_254),
.B(n_276),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_189),
.B(n_168),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_245),
.B(n_252),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_216),
.B(n_226),
.C(n_208),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_246),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_176),
.A2(n_160),
.B(n_151),
.C(n_129),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_286),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_190),
.B(n_130),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_215),
.A2(n_147),
.B(n_160),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_290),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_186),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_258),
.B(n_263),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_179),
.A2(n_160),
.B(n_151),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_260),
.A2(n_31),
.B(n_7),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_201),
.B1(n_197),
.B2(n_175),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_194),
.B(n_142),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_264),
.B(n_267),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_185),
.B(n_129),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_212),
.A2(n_135),
.B1(n_161),
.B2(n_159),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_212),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_274),
.B(n_280),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g276 ( 
.A(n_213),
.B(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_182),
.B(n_155),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_211),
.A2(n_133),
.B1(n_155),
.B2(n_135),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_191),
.A2(n_112),
.B1(n_172),
.B2(n_38),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_288),
.B1(n_229),
.B2(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_223),
.B(n_172),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_285),
.B(n_256),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_184),
.B(n_172),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_203),
.A2(n_112),
.B1(n_110),
.B2(n_151),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_311),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_211),
.B1(n_206),
.B2(n_229),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_SL g351 ( 
.A1(n_296),
.A2(n_243),
.B(n_248),
.C(n_290),
.Y(n_351)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_177),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_299),
.B(n_319),
.C(n_332),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_246),
.A2(n_222),
.B1(n_220),
.B2(n_206),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_300),
.A2(n_335),
.B1(n_243),
.B2(n_254),
.Y(n_352)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_304),
.A2(n_317),
.B1(n_343),
.B2(n_283),
.Y(n_371)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_178),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_306),
.B(n_312),
.Y(n_349)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_258),
.B(n_228),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_313),
.B(n_318),
.Y(n_359)
);

INVx2_ASAP7_75t_R g314 ( 
.A(n_276),
.Y(n_314)
);

INVx11_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_232),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_321),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_235),
.B1(n_218),
.B2(n_187),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_207),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_202),
.C(n_221),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_209),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_333),
.Y(n_344)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_287),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_250),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_330),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_237),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_246),
.B(n_192),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_240),
.B(n_221),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_338),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_241),
.B(n_196),
.C(n_214),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_183),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_274),
.A2(n_188),
.B(n_230),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_334),
.A2(n_244),
.B(n_277),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_251),
.A2(n_210),
.B1(n_174),
.B2(n_233),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_275),
.B(n_241),
.CI(n_290),
.CON(n_336),
.SN(n_336)
);

OAI32xp33_ASAP7_75t_L g370 ( 
.A1(n_336),
.A2(n_277),
.A3(n_238),
.B1(n_265),
.B2(n_266),
.Y(n_370)
);

BUFx8_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

CKINVDCx10_ASAP7_75t_R g380 ( 
.A(n_337),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_240),
.B(n_3),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_267),
.B(n_5),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_265),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_342),
.B(n_277),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_251),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_346),
.B(n_384),
.Y(n_414)
);

AO22x1_ASAP7_75t_SL g347 ( 
.A1(n_300),
.A2(n_243),
.B1(n_272),
.B2(n_242),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_351),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_253),
.B(n_248),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_350),
.A2(n_364),
.B(n_376),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_352),
.A2(n_354),
.B1(n_356),
.B2(n_361),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_253),
.B1(n_243),
.B2(n_262),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_275),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_373),
.C(n_381),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_330),
.B1(n_313),
.B2(n_311),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_264),
.B1(n_290),
.B2(n_245),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_366),
.B(n_387),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_325),
.B(n_277),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_369),
.B(n_370),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_371),
.A2(n_301),
.B1(n_327),
.B2(n_323),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_299),
.B(n_238),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_341),
.A2(n_280),
.B1(n_288),
.B2(n_266),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_375),
.A2(n_295),
.B1(n_314),
.B2(n_338),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_303),
.A2(n_310),
.B(n_337),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_260),
.B1(n_273),
.B2(n_239),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_377),
.A2(n_296),
.B1(n_340),
.B2(n_297),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_294),
.B(n_286),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_383),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_255),
.C(n_270),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_303),
.B(n_255),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_388),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_294),
.B(n_239),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_269),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_298),
.A2(n_292),
.B(n_289),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_298),
.B(n_334),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_308),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_292),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_354),
.A2(n_343),
.B1(n_336),
.B2(n_293),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_404),
.B1(n_407),
.B2(n_369),
.Y(n_435)
);

XOR2x1_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_314),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_391),
.B(n_378),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_348),
.A2(n_337),
.B1(n_328),
.B2(n_320),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_380),
.Y(n_439)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_394),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_326),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_399),
.C(n_413),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_331),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_401),
.A2(n_408),
.B1(n_409),
.B2(n_420),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_349),
.B(n_305),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_405),
.B(n_426),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_361),
.A2(n_296),
.B1(n_332),
.B2(n_302),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_348),
.A2(n_296),
.B1(n_309),
.B2(n_328),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_324),
.Y(n_410)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_348),
.B1(n_367),
.B2(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_321),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_307),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_422),
.C(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

OR2x2_ASAP7_75t_SL g418 ( 
.A(n_376),
.B(n_269),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_418),
.Y(n_433)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_353),
.Y(n_419)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_375),
.A2(n_249),
.B1(n_289),
.B2(n_268),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_379),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_421),
.B(n_400),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_268),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_350),
.A2(n_249),
.B(n_281),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_425),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_344),
.B(n_281),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_385),
.Y(n_436)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_400),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_432),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_410),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_444),
.B1(n_392),
.B2(n_358),
.Y(n_474)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_398),
.B(n_370),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_437),
.B(n_398),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_SL g469 ( 
.A1(n_439),
.A2(n_448),
.B(n_402),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_396),
.A2(n_386),
.B1(n_359),
.B2(n_351),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_449),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_401),
.A2(n_351),
.B1(n_347),
.B2(n_372),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_397),
.B1(n_394),
.B2(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_414),
.B(n_372),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_452),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_374),
.Y(n_454)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_454),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_425),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_460),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_389),
.B(n_360),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_457),
.B(n_461),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_347),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_419),
.B(n_345),
.Y(n_459)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_380),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_395),
.B(n_357),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_469),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_438),
.A2(n_407),
.B1(n_397),
.B2(n_390),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_464),
.A2(n_471),
.B1(n_472),
.B2(n_480),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_416),
.C(n_422),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_470),
.C(n_475),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_416),
.C(n_399),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_351),
.B1(n_418),
.B2(n_413),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_474),
.A2(n_433),
.B1(n_440),
.B2(n_451),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_403),
.C(n_402),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_487),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_364),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_483),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_431),
.A2(n_455),
.B(n_444),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_479),
.A2(n_439),
.B(n_450),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_438),
.A2(n_358),
.B1(n_427),
.B2(n_345),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_437),
.B(n_357),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_249),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_485),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_435),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_17),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_8),
.Y(n_489)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_489),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_431),
.B(n_8),
.C(n_9),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_442),
.C(n_434),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_450),
.Y(n_491)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_491),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_515),
.B(n_478),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_466),
.A2(n_460),
.B(n_439),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_503),
.Y(n_527)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_501),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_533)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_505),
.C(n_506),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_470),
.C(n_475),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_454),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_507),
.A2(n_509),
.B1(n_511),
.B2(n_514),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_441),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_510),
.C(n_513),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_463),
.B(n_456),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_434),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_464),
.A2(n_432),
.B1(n_429),
.B2(n_443),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_479),
.B(n_442),
.C(n_441),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_481),
.A2(n_443),
.B1(n_430),
.B2(n_458),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_L g515 ( 
.A1(n_478),
.A2(n_430),
.B(n_436),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_471),
.B(n_472),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_518),
.A2(n_521),
.B(n_528),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_494),
.B(n_465),
.C(n_462),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_522),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_465),
.C(n_482),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_467),
.C(n_487),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_526),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_459),
.C(n_447),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_491),
.A2(n_447),
.B(n_490),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_491),
.A2(n_501),
.B(n_515),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_529),
.B(n_531),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_512),
.A2(n_9),
.B(n_10),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_498),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_16),
.B1(n_17),
.B2(n_528),
.Y(n_549)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_533),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_513),
.A2(n_11),
.B(n_15),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_534),
.A2(n_508),
.B(n_497),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_524),
.B(n_496),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_537),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_510),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_504),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_538),
.B(n_542),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_502),
.Y(n_543)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_543),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_497),
.C(n_492),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_546),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_517),
.B(n_492),
.C(n_502),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_517),
.B(n_15),
.C(n_16),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_548),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_523),
.B(n_15),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_550),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_16),
.C(n_526),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_16),
.C(n_529),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_531),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_545),
.A2(n_521),
.B(n_520),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_552),
.A2(n_562),
.B1(n_535),
.B2(n_532),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_537),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_560),
.C(n_563),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_558),
.B(n_560),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_520),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_551),
.A2(n_525),
.B(n_530),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_525),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_539),
.A2(n_530),
.B(n_534),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_564),
.A2(n_562),
.B(n_561),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_544),
.C(n_550),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_566),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_552),
.A2(n_540),
.B1(n_533),
.B2(n_547),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_570),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_555),
.B(n_540),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_569),
.B(n_571),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_554),
.A2(n_559),
.B(n_553),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_557),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_565),
.A2(n_556),
.B(n_558),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_575),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_567),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_579),
.A2(n_580),
.B(n_573),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_574),
.B(n_568),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_581),
.A2(n_582),
.B(n_576),
.Y(n_583)
);

BUFx24_ASAP7_75t_SL g582 ( 
.A(n_578),
.Y(n_582)
);

BUFx24_ASAP7_75t_SL g584 ( 
.A(n_583),
.Y(n_584)
);


endmodule