module real_jpeg_28678_n_7 (n_5, n_4, n_0, n_24, n_1, n_26, n_2, n_25, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_24;
input n_1;
input n_26;
input n_2;
input n_25;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_11;
wire n_14;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_25),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_26),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_24),
.Y(n_13)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g7 ( 
.A1(n_5),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

OAI221xp5_ASAP7_75t_L g10 ( 
.A1(n_6),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_16),
.B(n_18),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_14),
.B(n_15),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);


endmodule