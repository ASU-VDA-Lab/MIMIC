module fake_netlist_6_717_n_18607 (n_2542, n_1671, n_2817, n_801, n_4452, n_2576, n_4649, n_1674, n_741, n_1351, n_1212, n_208, n_4251, n_2157, n_5019, n_2332, n_3849, n_578, n_5138, n_4388, n_4395, n_1061, n_3089, n_783, n_4978, n_188, n_1854, n_3088, n_3257, n_1342, n_4829, n_1387, n_3222, n_677, n_4699, n_1151, n_4686, n_2317, n_442, n_1975, n_1930, n_3706, n_2179, n_5055, n_1547, n_3376, n_4868, n_893, n_3801, n_4249, n_1192, n_3564, n_1844, n_1555, n_5057, n_3030, n_830, n_65, n_447, n_2838, n_3427, n_852, n_5101, n_2628, n_3071, n_2926, n_1078, n_544, n_4273, n_35, n_2321, n_2019, n_5102, n_3345, n_2074, n_2919, n_4501, n_2129, n_4724, n_945, n_4997, n_2399, n_4843, n_1232, n_4696, n_4347, n_2480, n_3877, n_3929, n_3048, n_1455, n_2786, n_567, n_1781, n_1971, n_2004, n_1106, n_4814, n_953, n_3979, n_3077, n_2873, n_3452, n_3107, n_155, n_4956, n_454, n_1421, n_3664, n_1936, n_5129, n_1660, n_5070, n_3047, n_4414, n_112, n_713, n_1400, n_2625, n_4646, n_2843, n_3760, n_48, n_1560, n_4262, n_734, n_1088, n_1894, n_3347, n_5136, n_907, n_6, n_4110, n_1658, n_4950, n_4729, n_4268, n_1967, n_3999, n_3928, n_2613, n_3535, n_4751, n_44, n_2708, n_1648, n_5151, n_1911, n_2011, n_281, n_564, n_279, n_686, n_4102, n_1641, n_3871, n_2735, n_4662, n_4671, n_3959, n_2268, n_1367, n_1336, n_4314, n_2080, n_323, n_5099, n_1381, n_331, n_1699, n_2093, n_4296, n_102, n_2770, n_608, n_2101, n_4507, n_32, n_512, n_3484, n_4677, n_792, n_5063, n_1328, n_2917, n_2616, n_3923, n_3900, n_3488, n_939, n_2811, n_3732, n_2832, n_4226, n_1762, n_1910, n_1075, n_3980, n_2998, n_4366, n_3446, n_237, n_1895, n_4294, n_4698, n_4445, n_4810, n_3859, n_2692, n_175, n_3914, n_4456, n_3397, n_3575, n_2469, n_3927, n_3888, n_764, n_2764, n_2895, n_733, n_2922, n_3882, n_4856, n_3492, n_4369, n_30, n_2068, n_4331, n_4972, n_1290, n_4993, n_2072, n_1354, n_586, n_423, n_4375, n_1701, n_2678, n_3935, n_5130, n_4291, n_88, n_1726, n_4613, n_2434, n_2878, n_3012, n_3875, n_1167, n_2428, n_4717, n_4877, n_3247, n_871, n_210, n_2641, n_4731, n_3052, n_178, n_355, n_5046, n_2749, n_3298, n_2254, n_5058, n_1926, n_3273, n_4467, n_1747, n_195, n_780, n_2624, n_2350, n_5042, n_4681, n_4072, n_4752, n_4220, n_835, n_928, n_2092, n_1654, n_1750, n_1462, n_2514, n_604, n_1588, n_3942, n_3997, n_26, n_2468, n_4381, n_5144, n_515, n_2096, n_3968, n_4466, n_4418, n_3434, n_4510, n_4473, n_514, n_687, n_890, n_2812, n_190, n_4518, n_1709, n_2393, n_2657, n_2921, n_2136, n_2409, n_2252, n_3237, n_949, n_3500, n_3834, n_4589, n_2075, n_2972, n_3542, n_91, n_2763, n_2762, n_3192, n_760, n_1546, n_4394, n_2279, n_161, n_1296, n_3352, n_3073, n_2150, n_1294, n_3696, n_1420, n_4082, n_595, n_1779, n_524, n_4921, n_1858, n_4329, n_5135, n_3021, n_2558, n_1164, n_4697, n_4288, n_4289, n_3763, n_2712, n_3733, n_1487, n_3614, n_874, n_382, n_2145, n_898, n_4964, n_4228, n_3423, n_925, n_1932, n_1101, n_15, n_4636, n_4322, n_3644, n_1249, n_4946, n_2706, n_4767, n_4287, n_2693, n_4137, n_1127, n_1512, n_1451, n_320, n_639, n_963, n_2767, n_4576, n_4615, n_1139, n_3179, n_1018, n_3400, n_1521, n_1366, n_4000, n_2897, n_4389, n_3970, n_4345, n_996, n_532, n_173, n_1376, n_413, n_4664, n_2170, n_4156, n_948, n_977, n_536, n_3158, n_1788, n_4873, n_2643, n_3782, n_1835, n_3470, n_5076, n_581, n_4713, n_4098, n_5026, n_4476, n_432, n_3700, n_4995, n_3166, n_3104, n_3435, n_842, n_2239, n_4310, n_1432, n_989, n_2689, n_1473, n_2191, n_1246, n_4528, n_899, n_1035, n_4914, n_4939, n_499, n_1426, n_3418, n_705, n_11, n_1004, n_1529, n_2473, n_4634, n_2069, n_2362, n_4096, n_2539, n_2698, n_4123, n_3119, n_3735, n_2297, n_4379, n_486, n_4718, n_1448, n_3631, n_648, n_2445, n_2057, n_2103, n_3770, n_2772, n_4440, n_4402, n_927, n_5052, n_4541, n_5009, n_4872, n_929, n_4551, n_2857, n_1183, n_4627, n_4079, n_2494, n_3342, n_998, n_5035, n_717, n_1383, n_3390, n_3656, n_1424, n_1000, n_3025, n_2137, n_1626, n_1507, n_2482, n_3810, n_552, n_4798, n_2532, n_1388, n_3006, n_216, n_912, n_5010, n_2296, n_3633, n_5089, n_2849, n_1201, n_1398, n_884, n_4592, n_1395, n_2199, n_2661, n_731, n_1955, n_931, n_474, n_312, n_1791, n_66, n_958, n_5137, n_100, n_3331, n_5104, n_1897, n_2064, n_2773, n_589, n_3606, n_1310, n_819, n_1334, n_3591, n_2788, n_964, n_4756, n_2797, n_4746, n_124, n_3892, n_4970, n_4069, n_211, n_2748, n_1834, n_2331, n_2292, n_3441, n_3534, n_3964, n_2416, n_311, n_1877, n_3944, n_1939, n_2030, n_1769, n_556, n_2209, n_3605, n_1602, n_4633, n_3306, n_276, n_3026, n_221, n_4584, n_3090, n_3724, n_4276, n_5116, n_2990, n_3847, n_1773, n_5001, n_2552, n_1053, n_4428, n_1533, n_3323, n_4, n_266, n_2274, n_518, n_4618, n_4679, n_1745, n_914, n_3479, n_4496, n_317, n_4805, n_1679, n_90, n_3454, n_2160, n_2146, n_2131, n_488, n_3547, n_2575, n_5100, n_4410, n_1933, n_1179, n_324, n_3816, n_4807, n_4411, n_3214, n_1243, n_301, n_2928, n_5166, n_1917, n_1580, n_2822, n_36, n_4180, n_1281, n_3109, n_3354, n_2572, n_1520, n_3126, n_3663, n_2863, n_1419, n_3299, n_351, n_259, n_1731, n_2135, n_4707, n_1645, n_1832, n_4676, n_858, n_2049, n_956, n_663, n_4880, n_3566, n_2781, n_4126, n_410, n_2829, n_1696, n_3845, n_1594, n_664, n_1869, n_3804, n_4207, n_2016, n_4470, n_580, n_4813, n_1030, n_3901, n_1937, n_465, n_1790, n_4014, n_4704, n_341, n_1744, n_828, n_2142, n_4252, n_607, n_4028, n_2448, n_4048, n_4596, n_4444, n_3756, n_3406, n_820, n_951, n_952, n_3919, n_2263, n_974, n_4952, n_2656, n_5023, n_2375, n_1934, n_628, n_1434, n_1573, n_3981, n_3973, n_2756, n_807, n_4761, n_1275, n_2884, n_485, n_67, n_1510, n_3120, n_3797, n_238, n_2024, n_1595, n_4770, n_202, n_1749, n_3474, n_2549, n_4690, n_1669, n_1024, n_3864, n_4932, n_248, n_2302, n_1667, n_1037, n_5143, n_3592, n_468, n_4230, n_2637, n_1639, n_183, n_3967, n_3195, n_466, n_2526, n_4274, n_3277, n_2548, n_991, n_4189, n_3817, n_340, n_1108, n_3659, n_2559, n_2177, n_39, n_2595, n_5003, n_4827, n_1601, n_1960, n_2694, n_3648, n_1686, n_3042, n_5094, n_4610, n_4472, n_3228, n_3657, n_96, n_3081, n_1430, n_1316, n_1287, n_1586, n_2264, n_3464, n_380, n_3723, n_1190, n_397, n_4380, n_4990, n_4996, n_4398, n_2498, n_4515, n_1891, n_5031, n_1213, n_2235, n_4193, n_3570, n_5082, n_1673, n_3828, n_172, n_2392, n_3424, n_4131, n_239, n_97, n_2298, n_2326, n_1539, n_490, n_3594, n_1043, n_4090, n_4165, n_2305, n_2120, n_80, n_4626, n_4144, n_2964, n_352, n_2169, n_3485, n_4077, n_2371, n_1361, n_662, n_3262, n_4008, n_3356, n_1642, n_3210, n_937, n_4689, n_1682, n_4547, n_3329, n_330, n_3826, n_4905, n_1406, n_4601, n_962, n_3647, n_3681, n_1883, n_4300, n_1288, n_1186, n_4623, n_5007, n_3320, n_2518, n_3988, n_1720, n_3476, n_4842, n_204, n_482, n_3439, n_4135, n_2688, n_394, n_1845, n_1489, n_942, n_2798, n_2852, n_1524, n_1964, n_1920, n_2753, n_1496, n_3292, n_2007, n_2039, n_1225, n_1544, n_1485, n_1846, n_3437, n_4111, n_533, n_3712, n_4608, n_879, n_2310, n_2506, n_4859, n_94, n_2626, n_1567, n_4037, n_3562, n_2973, n_41, n_3665, n_273, n_3007, n_3528, n_4571, n_3698, n_3355, n_2454, n_2114, n_3174, n_1066, n_1948, n_157, n_4215, n_2154, n_1484, n_4185, n_3752, n_2283, n_5145, n_4219, n_1229, n_1373, n_3958, n_3985, n_2427, n_4196, n_1447, n_4774, n_2056, n_4242, n_5109, n_3389, n_4232, n_4190, n_4902, n_3000, n_5149, n_2680, n_1047, n_3375, n_3899, n_1385, n_3713, n_1931, n_502, n_2668, n_1257, n_3197, n_4987, n_2128, n_4736, n_2398, n_1725, n_3743, n_834, n_5033, n_2695, n_4035, n_3818, n_3124, n_1741, n_1002, n_1949, n_3759, n_545, n_2671, n_4516, n_2715, n_1804, n_251, n_2508, n_3511, n_2054, n_1337, n_1477, n_2614, n_4492, n_2833, n_2758, n_3694, n_2937, n_4789, n_4376, n_1001, n_2241, n_4708, n_4657, n_1690, n_1191, n_1076, n_4512, n_1378, n_855, n_1377, n_695, n_4081, n_1542, n_4542, n_4462, n_1716, n_278, n_4931, n_4536, n_3303, n_978, n_4324, n_384, n_1976, n_4382, n_2905, n_1291, n_749, n_1824, n_3954, n_2122, n_2140, n_3503, n_3160, n_1065, n_1255, n_568, n_5124, n_143, n_3951, n_823, n_1074, n_698, n_3569, n_739, n_3874, n_2528, n_5123, n_4639, n_1338, n_1097, n_3027, n_781, n_4083, n_1810, n_182, n_573, n_1583, n_4480, n_1730, n_2295, n_2746, n_389, n_814, n_1643, n_2020, n_4171, n_3652, n_222, n_4023, n_1105, n_721, n_1461, n_742, n_691, n_3617, n_2076, n_3567, n_377, n_1598, n_4344, n_2935, n_4705, n_4046, n_3807, n_918, n_1114, n_56, n_763, n_4027, n_3154, n_1227, n_2485, n_3898, n_3520, n_191, n_4391, n_946, n_1303, n_4095, n_2881, n_1116, n_1570, n_1702, n_1219, n_3551, n_4947, n_3064, n_1780, n_3897, n_1689, n_8, n_3372, n_1944, n_1347, n_795, n_1221, n_1245, n_3215, n_448, n_3853, n_4740, n_4631, n_1561, n_1112, n_2081, n_2168, n_5068, n_234, n_1460, n_911, n_82, n_27, n_5159, n_2862, n_472, n_2615, n_4068, n_4625, n_2474, n_3703, n_2437, n_2444, n_25, n_3962, n_2743, n_4766, n_4863, n_2267, n_3035, n_668, n_4166, n_1821, n_1058, n_3378, n_3745, n_3362, n_4744, n_103, n_4188, n_2934, n_3667, n_3523, n_2222, n_712, n_3176, n_31, n_2505, n_334, n_4817, n_4115, n_2999, n_2014, n_1239, n_3697, n_1584, n_470, n_3680, n_2408, n_3468, n_5045, n_1972, n_4383, n_4491, n_455, n_363, n_4486, n_1816, n_393, n_503, n_3024, n_4612, n_2531, n_5163, n_307, n_4529, n_500, n_3361, n_714, n_3478, n_3936, n_1349, n_291, n_2723, n_2800, n_3496, n_4390, n_3096, n_2651, n_2095, n_3239, n_3161, n_2799, n_3902, n_4062, n_3295, n_4396, n_1998, n_1574, n_3101, n_240, n_756, n_1981, n_4233, n_1606, n_3374, n_2640, n_253, n_1552, n_2918, n_583, n_3288, n_4307, n_3992, n_3876, n_249, n_3125, n_4293, n_941, n_3552, n_1031, n_115, n_849, n_4684, n_3116, n_4091, n_1753, n_5027, n_3095, n_2471, n_4412, n_2807, n_1921, n_3618, n_4580, n_1055, n_2217, n_2197, n_4758, n_4781, n_4148, n_2461, n_271, n_206, n_4057, n_633, n_1170, n_308, n_3444, n_1040, n_3059, n_2634, n_1761, n_1890, n_3017, n_1805, n_2477, n_2308, n_2333, n_3001, n_1089, n_3795, n_3852, n_1365, n_4138, n_5018, n_3815, n_3896, n_3274, n_4457, n_4093, n_1616, n_1862, n_339, n_434, n_64, n_288, n_4928, n_4794, n_722, n_2223, n_4197, n_4482, n_629, n_1621, n_2547, n_2415, n_5073, n_827, n_4834, n_4762, n_192, n_3113, n_992, n_3813, n_3660, n_3766, n_1613, n_1458, n_1027, n_3266, n_3574, n_1189, n_223, n_4154, n_4907, n_5077, n_5034, n_726, n_50, n_4504, n_365, n_3844, n_1237, n_2534, n_4975, n_3741, n_2451, n_2243, n_4815, n_4898, n_3443, n_509, n_4819, n_1209, n_1708, n_805, n_396, n_350, n_78, n_2051, n_4370, n_2359, n_5112, n_480, n_142, n_1402, n_1691, n_3332, n_4134, n_1238, n_2570, n_4092, n_4645, n_3668, n_2491, n_1264, n_4755, n_4359, n_4960, n_4087, n_1700, n_4933, n_5091, n_3487, n_4591, n_287, n_4302, n_5111, n_3340, n_230, n_461, n_873, n_3946, n_2989, n_3395, n_4474, n_2509, n_2513, n_3757, n_4178, n_5165, n_1704, n_2247, n_250, n_1711, n_4884, n_1579, n_3275, n_836, n_522, n_3678, n_3440, n_2094, n_1511, n_2356, n_1422, n_1772, n_4692, n_616, n_3165, n_1119, n_1433, n_1902, n_1842, n_1620, n_2739, n_1735, n_3890, n_1541, n_1300, n_641, n_3750, n_1313, n_3607, n_3316, n_516, n_2418, n_2864, n_4311, n_1180, n_2703, n_3371, n_4722, n_4606, n_3261, n_666, n_4187, n_940, n_2058, n_405, n_213, n_2660, n_1094, n_4962, n_4563, n_494, n_5056, n_4820, n_2394, n_3532, n_3948, n_2124, n_4619, n_381, n_4327, n_1961, n_3765, n_4125, n_5036, n_4221, n_3297, n_976, n_3067, n_2155, n_2686, n_2364, n_4392, n_2996, n_3803, n_2085, n_917, n_5014, n_3639, n_4334, n_659, n_3351, n_808, n_4047, n_3413, n_1193, n_3412, n_3791, n_3164, n_4575, n_551, n_699, n_4320, n_3884, n_451, n_5139, n_757, n_594, n_2190, n_3438, n_166, n_4141, n_2850, n_572, n_1481, n_1441, n_3373, n_92, n_2104, n_513, n_3883, n_261, n_3728, n_2925, n_4499, n_121, n_433, n_3949, n_2792, n_219, n_3315, n_263, n_3798, n_788, n_1543, n_1599, n_329, n_4257, n_4458, n_2674, n_5103, n_4641, n_4720, n_4893, n_61, n_3857, n_1876, n_4107, n_243, n_1873, n_3630, n_3518, n_1866, n_117, n_2130, n_1330, n_1413, n_3714, n_2228, n_5039, n_2455, n_2876, n_4772, n_3099, n_4468, n_4161, n_1663, n_4172, n_3403, n_2714, n_2245, n_4961, n_4454, n_1107, n_2457, n_3294, n_4119, n_3686, n_4502, n_318, n_2971, n_1713, n_715, n_4277, n_4526, n_1265, n_3490, n_4849, n_530, n_277, n_4319, n_3369, n_618, n_199, n_3581, n_3069, n_2028, n_3715, n_1069, n_612, n_3725, n_3933, n_1175, n_2311, n_429, n_1012, n_3691, n_4485, n_4066, n_903, n_4146, n_1802, n_1504, n_4340, n_286, n_254, n_3961, n_4855, n_1801, n_2347, n_3917, n_47, n_816, n_1188, n_2206, n_4004, n_2967, n_2916, n_4292, n_2467, n_267, n_3145, n_1124, n_1624, n_3983, n_4940, n_3538, n_3280, n_1515, n_961, n_4356, n_3510, n_2824, n_593, n_637, n_2377, n_701, n_950, n_3009, n_3719, n_2525, n_4361, n_3827, n_891, n_5154, n_2067, n_3889, n_2687, n_1630, n_2887, n_4245, n_4136, n_3526, n_2194, n_2619, n_4367, n_1987, n_507, n_968, n_2271, n_1008, n_2583, n_4560, n_2606, n_4899, n_1033, n_462, n_1052, n_2794, n_5164, n_2391, n_304, n_2431, n_125, n_2078, n_2932, n_1767, n_3431, n_3450, n_449, n_4663, n_2893, n_1208, n_2954, n_2728, n_1072, n_815, n_3421, n_3183, n_2493, n_4802, n_2705, n_1067, n_3405, n_255, n_284, n_1952, n_5074, n_4044, n_3436, n_1026, n_1880, n_3442, n_3366, n_2631, n_38, n_289, n_3937, n_1293, n_3159, n_4701, n_108, n_794, n_727, n_894, n_685, n_353, n_3240, n_3576, n_1863, n_3385, n_4851, n_3293, n_872, n_3922, n_86, n_847, n_644, n_682, n_851, n_4991, n_72, n_2554, n_1513, n_1913, n_4934, n_837, n_5087, n_2517, n_2713, n_5000, n_2765, n_2590, n_3150, n_2060, n_4479, n_2608, n_4011, n_5131, n_1959, n_3133, n_765, n_1492, n_1340, n_4688, n_4753, n_4058, n_631, n_2262, n_3611, n_3082, n_4848, n_5059, n_156, n_843, n_2604, n_2407, n_1277, n_2816, n_3799, n_2574, n_4475, n_2675, n_3537, n_4443, n_3887, n_1022, n_614, n_2667, n_4587, n_1615, n_4114, n_1474, n_1571, n_2948, n_1577, n_2119, n_947, n_1117, n_1992, n_3223, n_3140, n_3185, n_4749, n_2605, n_5155, n_118, n_926, n_3654, n_1849, n_2848, n_919, n_1698, n_4100, n_4264, n_3788, n_89, n_4891, n_777, n_1299, n_3837, n_2718, n_1436, n_1384, n_3325, n_2238, n_4085, n_4464, n_4624, n_4818, n_4659, n_3600, n_18, n_5015, n_4339, n_1178, n_98, n_2338, n_3324, n_796, n_1195, n_184, n_1811, n_1857, n_3987, n_1519, n_2144, n_1284, n_1604, n_4487, n_4889, n_4866, n_1142, n_623, n_1048, n_3638, n_4816, n_2110, n_1502, n_1659, n_3393, n_3451, n_1418, n_1250, n_292, n_4937, n_3615, n_3072, n_3087, n_2053, n_2259, n_2121, n_4222, n_4874, n_4401, n_889, n_2710, n_3142, n_4015, n_1966, n_477, n_1110, n_4709, n_2213, n_4976, n_2389, n_2132, n_2892, n_4120, n_1564, n_4658, n_231, n_2860, n_2330, n_40, n_1457, n_505, n_3718, n_1787, n_537, n_1993, n_2281, n_2617, n_2776, n_1466, n_10, n_1919, n_3705, n_3211, n_3909, n_546, n_386, n_1220, n_1893, n_2301, n_4665, n_3582, n_4223, n_2387, n_3270, n_2846, n_970, n_2488, n_1980, n_2237, n_1060, n_1951, n_444, n_4362, n_1252, n_3311, n_3913, n_1223, n_511, n_5121, n_1286, n_2115, n_4430, n_3302, n_4348, n_5013, n_1597, n_4489, n_4839, n_2596, n_3163, n_775, n_4404, n_1153, n_439, n_1531, n_2828, n_453, n_2384, n_4261, n_4204, n_759, n_2724, n_426, n_2585, n_4825, n_2352, n_1625, n_3986, n_5006, n_4513, n_4006, n_2226, n_2801, n_1901, n_3869, n_2556, n_4747, n_1647, n_3753, n_2306, n_1614, n_1892, n_3742, n_3683, n_4801, n_401, n_3260, n_2550, n_3175, n_3736, n_4448, n_1096, n_2227, n_3284, n_4869, n_427, n_2159, n_4386, n_688, n_1077, n_2315, n_4132, n_2995, n_1437, n_4844, n_4438, n_4836, n_4955, n_4149, n_4355, n_501, n_2276, n_3234, n_856, n_2803, n_379, n_1668, n_2777, n_3202, n_2830, n_3220, n_1129, n_602, n_2181, n_171, n_2911, n_169, n_4655, n_1429, n_2826, n_3429, n_2379, n_326, n_587, n_3554, n_1593, n_1202, n_1635, n_4067, n_4357, n_28, n_3462, n_2851, n_4374, n_5132, n_106, n_358, n_160, n_2420, n_3722, n_186, n_4400, n_4846, n_2984, n_575, n_4024, n_1508, n_732, n_2983, n_2240, n_392, n_2538, n_724, n_3250, n_1042, n_4582, n_1728, n_557, n_1871, n_4860, n_845, n_140, n_3414, n_1549, n_4870, n_768, n_3651, n_2102, n_2563, n_4989, n_3449, n_1683, n_1916, n_2598, n_597, n_280, n_1187, n_4304, n_4558, n_1403, n_4488, n_3767, n_2544, n_3550, n_4211, n_1206, n_4016, n_621, n_750, n_4656, n_3839, n_2823, n_4915, n_4328, n_1057, n_2785, n_235, n_1997, n_2636, n_3131, n_710, n_1818, n_3730, n_1298, n_4397, n_3399, n_2088, n_1611, n_5050, n_2740, n_746, n_4808, n_3416, n_3498, n_2401, n_101, n_1589, n_4712, n_2309, n_2900, n_2957, n_1740, n_2737, n_3994, n_1497, n_133, n_3672, n_3533, n_1622, n_4725, n_4406, n_1694, n_1535, n_3382, n_3132, n_2571, n_3138, n_20, n_5053, n_2171, n_2988, n_4908, n_3136, n_1350, n_4109, n_4192, n_4824, n_2037, n_2808, n_4567, n_5150, n_782, n_809, n_3819, n_4778, n_1797, n_986, n_2050, n_4595, n_2164, n_4174, n_402, n_1870, n_1171, n_460, n_1827, n_4904, n_2187, n_1152, n_450, n_3544, n_4150, n_2904, n_711, n_3105, n_2872, n_3692, n_4616, n_4982, n_370, n_1695, n_2046, n_2272, n_2760, n_1979, n_4643, n_2738, n_972, n_1332, n_4323, n_624, n_2346, n_4831, n_936, n_3045, n_3821, n_885, n_83, n_2342, n_2167, n_2970, n_3676, n_4896, n_2882, n_3666, n_3675, n_4017, n_4260, n_4916, n_2541, n_2940, n_4739, n_599, n_105, n_1974, n_4122, n_934, n_4209, n_2768, n_3858, n_1341, n_4298, n_2314, n_3502, n_3003, n_4128, n_543, n_5147, n_4271, n_4644, n_1355, n_2258, n_325, n_804, n_2390, n_959, n_2562, n_4716, n_4312, n_1343, n_1522, n_76, n_2734, n_1782, n_707, n_1900, n_5048, n_3246, n_1548, n_3381, n_1155, n_2195, n_3208, n_4944, n_4343, n_4715, n_4935, n_4694, n_4672, n_5054, n_2962, n_2939, n_1672, n_1925, n_4407, n_737, n_4045, n_3517, n_2945, n_4598, n_3061, n_3893, n_3932, n_21, n_3469, n_2960, n_138, n_3258, n_4524, n_3143, n_333, n_4084, n_3149, n_3365, n_3379, n_24, n_459, n_4850, n_4424, n_3008, n_1751, n_2840, n_285, n_3939, n_4776, n_1375, n_3972, n_4153, n_85, n_3506, n_1650, n_1962, n_3855, n_1928, n_3091, n_4317, n_4723, n_4269, n_4088, n_3398, n_2761, n_2793, n_3776, n_3711, n_4235, n_1019, n_4143, n_4170, n_729, n_876, n_774, n_3642, n_2845, n_4650, n_438, n_4719, n_1860, n_5016, n_1904, n_2874, n_1200, n_2588, n_479, n_1353, n_1777, n_4967, n_3308, n_1113, n_1600, n_2253, n_2366, n_4912, n_4799, n_2261, n_4423, n_5086, n_2210, n_4735, n_3602, n_187, n_3300, n_2978, n_2516, n_1050, n_1411, n_2827, n_1177, n_3515, n_1150, n_566, n_1023, n_2951, n_1118, n_194, n_2949, n_1807, n_5028, n_1814, n_1631, n_1879, n_256, n_440, n_3806, n_2931, n_209, n_367, n_2569, n_3866, n_671, n_4543, n_740, n_703, n_4157, n_4229, n_3865, n_4073, n_1324, n_3629, n_1435, n_3920, n_969, n_4892, n_3255, n_1401, n_1516, n_3846, n_180, n_3512, n_2029, n_4439, n_1394, n_1326, n_4783, n_1379, n_214, n_935, n_4910, n_1130, n_3083, n_676, n_832, n_3049, n_5142, n_3830, n_3679, n_3541, n_74, n_3117, n_4930, n_372, n_111, n_314, n_378, n_338, n_1283, n_2385, n_4112, n_506, n_360, n_2149, n_2396, n_4557, n_4917, n_895, n_2450, n_3739, n_4432, n_2284, n_4352, n_4416, n_4593, n_344, n_2769, n_4465, n_3622, n_5114, n_4980, n_1392, n_4495, n_5117, n_1924, n_525, n_2463, n_3363, n_1677, n_611, n_3721, n_3062, n_2679, n_5024, n_4559, n_838, n_3969, n_129, n_3336, n_4160, n_4231, n_2952, n_1017, n_4256, n_2779, n_4938, n_109, n_445, n_930, n_2620, n_5162, n_1945, n_1656, n_2112, n_1464, n_2430, n_653, n_1414, n_2721, n_944, n_4335, n_2034, n_576, n_270, n_2683, n_563, n_2744, n_1011, n_4521, n_1566, n_626, n_990, n_3204, n_1104, n_4920, n_498, n_870, n_1253, n_366, n_1693, n_3256, n_348, n_3802, n_376, n_2118, n_2111, n_390, n_2915, n_1148, n_2188, n_1989, n_2802, n_3643, n_2425, n_4265, n_2950, n_719, n_3060, n_3098, n_4105, n_1851, n_1090, n_4861, n_4064, n_4926, n_1518, n_1362, n_3123, n_3380, n_1829, n_1450, n_4828, n_1638, n_3038, n_570, n_1789, n_620, n_519, n_2523, n_2413, n_3769, n_1482, n_3863, n_3669, n_3130, n_4316, n_4640, n_5122, n_1710, n_2161, n_1301, n_2805, n_33, n_4769, n_2282, n_4628, n_2047, n_1609, n_3344, n_2334, n_5133, n_409, n_1763, n_3989, n_2490, n_4460, n_4108, n_635, n_3786, n_3841, n_4254, n_1996, n_2867, n_1442, n_2726, n_4303, n_1158, n_2248, n_5011, n_2662, n_4909, n_3147, n_753, n_3925, n_3180, n_2795, n_3472, n_5106, n_269, n_359, n_1479, n_4768, n_1675, n_3717, n_571, n_2215, n_404, n_158, n_1884, n_665, n_2055, n_5156, n_2553, n_149, n_632, n_2038, n_4447, n_4826, n_3445, n_373, n_87, n_1833, n_3903, n_1494, n_2325, n_1850, n_3854, n_3235, n_1417, n_3673, n_4281, n_681, n_4648, n_3094, n_412, n_965, n_1428, n_1576, n_1856, n_2077, n_1059, n_4951, n_422, n_4957, n_3079, n_165, n_4360, n_540, n_4039, n_457, n_3070, n_3800, n_4566, n_3263, n_4853, n_1748, n_3504, n_531, n_4272, n_2930, n_1025, n_3111, n_336, n_12, n_1885, n_3054, n_1538, n_1240, n_1, n_4730, n_1234, n_3254, n_3684, n_4670, n_4882, n_4620, n_3152, n_4738, n_3579, n_3335, n_4177, n_3783, n_700, n_1307, n_3178, n_4127, n_1003, n_168, n_2353, n_4099, n_4517, n_77, n_4168, n_1738, n_4490, n_1575, n_1923, n_2260, n_3952, n_3911, n_1688, n_4285, n_3465, n_1743, n_2997, n_1991, n_2386, n_5161, n_1724, n_3708, n_4078, n_3046, n_2956, n_1553, n_3619, n_1415, n_1370, n_1786, n_4198, n_2382, n_3754, n_2291, n_415, n_1371, n_383, n_2886, n_2974, n_4213, n_200, n_2184, n_2982, n_1803, n_4065, n_229, n_2645, n_3904, n_1393, n_1517, n_1867, n_2630, n_1444, n_1603, n_2470, n_4446, n_1263, n_4417, n_4733, n_4764, n_1261, n_3879, n_2286, n_4743, n_2018, n_3080, n_1903, n_1143, n_658, n_1874, n_2865, n_2825, n_2013, n_2044, n_3023, n_3232, n_693, n_1056, n_758, n_2256, n_943, n_4060, n_5110, n_4879, n_42, n_772, n_2806, n_770, n_3028, n_3662, n_2981, n_3076, n_886, n_343, n_3624, n_1345, n_1820, n_4556, n_539, n_45, n_4117, n_4687, n_2836, n_638, n_1404, n_2378, n_887, n_2655, n_4600, n_126, n_1467, n_4250, n_3906, n_224, n_4954, n_1231, n_2599, n_3963, n_3368, n_9, n_2370, n_2612, n_2591, n_4881, n_1815, n_2214, n_4253, n_407, n_913, n_2593, n_4255, n_867, n_4071, n_3568, n_1230, n_3850, n_1333, n_2496, n_3313, n_4605, n_3189, n_163, n_1644, n_2725, n_2277, n_4691, n_1558, n_1732, n_2300, n_3943, n_4305, n_824, n_4297, n_2907, n_577, n_1843, n_619, n_4227, n_521, n_2778, n_395, n_1909, n_5020, n_606, n_1123, n_1309, n_2961, n_916, n_3934, n_4033, n_4415, n_483, n_1970, n_630, n_2059, n_2669, n_4094, n_4765, n_2546, n_3193, n_2522, n_476, n_4364, n_1957, n_4354, n_4732, n_3912, n_3118, n_3720, n_1907, n_2529, n_264, n_860, n_1530, n_4745, n_938, n_1302, n_4581, n_549, n_4377, n_2143, n_905, n_4792, n_1680, n_3842, n_322, n_993, n_689, n_2031, n_4878, n_1605, n_3514, n_4979, n_1988, n_558, n_2654, n_3036, n_966, n_4511, n_2908, n_3357, n_692, n_1233, n_3895, n_487, n_241, n_4520, n_3455, n_4118, n_4503, n_2176, n_2459, n_1111, n_3599, n_1251, n_2711, n_4199, n_1912, n_4441, n_1982, n_3872, n_3772, n_1312, n_5038, n_268, n_1760, n_4585, n_2664, n_5, n_1664, n_1722, n_3022, n_247, n_1165, n_4773, n_2008, n_2192, n_3281, n_2345, n_328, n_1386, n_4427, n_5113, n_3549, n_2804, n_2453, n_2676, n_3940, n_4822, n_1214, n_690, n_850, n_4800, n_1157, n_3453, n_3410, n_1752, n_1813, n_3768, n_4958, n_2810, n_4043, n_2319, n_825, n_3785, n_2963, n_2602, n_55, n_3873, n_2980, n_696, n_4886, n_1082, n_1317, n_3227, n_2733, n_3289, n_4055, n_2178, n_2644, n_2036, n_3326, n_4200, n_3460, n_2411, n_1796, n_2082, n_3519, n_678, n_5078, n_3707, n_283, n_3578, n_909, n_4737, n_590, n_4925, n_4116, n_362, n_22, n_1990, n_3805, n_2943, n_1634, n_3252, n_627, n_3253, n_1465, n_342, n_2622, n_2658, n_2665, n_2133, n_1712, n_4603, n_1523, n_1627, n_5080, n_3128, n_1527, n_495, n_2691, n_840, n_2913, n_4471, n_2230, n_1969, n_2690, n_1565, n_1493, n_2573, n_2646, n_2535, n_1364, n_3078, n_2436, n_615, n_3838, n_4651, n_3941, n_3793, n_4854, n_5071, n_3789, n_605, n_1514, n_3037, n_1646, n_3729, n_4994, n_2537, n_4483, n_5168, n_4661, n_1308, n_4988, n_3171, n_3608, n_4540, n_2097, n_79, n_3459, n_2853, n_1808, n_3053, n_3358, n_3499, n_4284, n_1005, n_1947, n_3426, n_4971, n_1469, n_5125, n_2650, n_987, n_720, n_153, n_3229, n_3348, n_1707, n_656, n_797, n_2933, n_2717, n_1723, n_1878, n_189, n_738, n_2012, n_3497, n_5066, n_2842, n_3580, n_2335, n_529, n_2307, n_3704, n_684, n_1809, n_4280, n_1181, n_37, n_3173, n_3677, n_3996, n_1049, n_4097, n_1666, n_803, n_4218, n_1717, n_1817, n_2449, n_3880, n_3685, n_2868, n_2231, n_3609, n_1228, n_417, n_4459, n_4545, n_272, n_2896, n_3019, n_2639, n_3471, n_2898, n_69, n_2368, n_53, n_458, n_4175, n_16, n_3200, n_4771, n_3259, n_2524, n_3167, n_2460, n_3867, n_3593, n_4455, n_1073, n_252, n_4514, n_3191, n_4140, n_2481, n_3561, n_4806, n_2682, n_3032, n_5160, n_2877, n_5098, n_1021, n_811, n_683, n_1207, n_5140, n_4992, n_880, n_3505, n_3540, n_3577, n_2432, n_150, n_1478, n_4796, n_3598, n_4442, n_2581, n_1363, n_3641, n_3777, n_4203, n_767, n_1837, n_2218, n_4533, n_831, n_3590, n_2435, n_954, n_4419, n_1410, n_1382, n_1736, n_4053, n_1483, n_3848, n_1372, n_3327, n_1719, n_319, n_2701, n_2511, n_4167, n_1427, n_2745, n_1080, n_123, n_562, n_2323, n_2784, n_162, n_4431, n_2421, n_1136, n_4387, n_2618, n_3265, n_2464, n_128, n_1125, n_3755, n_4042, n_5128, n_2224, n_2329, n_1092, n_441, n_4299, n_4890, n_146, n_1784, n_3571, n_193, n_1775, n_2410, n_1093, n_1783, n_2929, n_4176, n_296, n_651, n_3407, n_217, n_1185, n_3856, n_4236, n_3425, n_215, n_3894, n_3127, n_1831, n_2621, n_3623, n_5079, n_54, n_1453, n_2502, n_3646, n_497, n_4830, n_4706, n_1315, n_4570, n_2754, n_1224, n_2783, n_3188, n_1459, n_2462, n_3243, n_1135, n_2889, n_4034, n_4056, n_4622, n_3960, n_1470, n_4887, n_2732, n_4693, n_4206, n_2249, n_1091, n_2000, n_3862, n_4267, n_2270, n_1425, n_5049, n_983, n_906, n_1390, n_2289, n_1733, n_2955, n_2158, n_4609, n_1855, n_3051, n_3367, n_385, n_1687, n_1439, n_2328, n_2859, n_2202, n_1331, n_613, n_736, n_3314, n_3525, n_2100, n_5157, n_2993, n_4754, n_3016, n_4647, n_1134, n_3688, n_4003, n_554, n_1995, n_3751, n_4894, n_4113, n_1889, n_4760, n_435, n_1905, n_3466, n_762, n_4983, n_1778, n_1079, n_2139, n_419, n_5083, n_4509, n_2875, n_1103, n_3907, n_3338, n_144, n_4217, n_4906, n_2219, n_1203, n_3636, n_2327, n_999, n_1254, n_2841, n_4897, n_3539, n_3291, n_4399, n_2304, n_2487, n_3276, n_2597, n_3194, n_5084, n_3572, n_349, n_3886, n_4710, n_4420, n_443, n_892, n_3637, n_4574, n_1468, n_2855, n_1859, n_2156, n_1718, n_4234, n_4101, n_3548, n_5017, n_1768, n_3974, n_198, n_1847, n_3634, n_1397, n_3236, n_901, n_2755, n_3141, n_923, n_5096, n_1841, n_4660, n_1623, n_1015, n_3112, n_4797, n_3108, n_4270, n_4151, n_4945, n_3417, n_4124, n_73, n_785, n_5153, n_609, n_4611, n_2337, n_1356, n_3213, n_4333, n_127, n_3820, n_2607, n_2890, n_1168, n_5115, n_1943, n_3249, n_1320, n_2722, n_1452, n_2854, n_2499, n_4152, n_302, n_137, n_1596, n_5092, n_1734, n_3172, n_4832, n_2902, n_3217, n_1983, n_1938, n_2472, n_3394, n_1715, n_3536, n_1443, n_1272, n_2894, n_3957, n_3710, n_4195, n_4554, n_3040, n_3279, n_2402, n_2225, n_1081, n_1692, n_1084, n_1864, n_2006, n_3402, n_3475, n_3501, n_374, n_1705, n_3905, n_4680, n_3013, n_921, n_579, n_2789, n_5152, n_2257, n_4927, n_4258, n_1828, n_2699, n_2200, n_650, n_1940, n_4548, n_4862, n_1405, n_2376, n_456, n_3878, n_2670, n_313, n_2700, n_1041, n_565, n_3134, n_1569, n_3115, n_1062, n_896, n_4553, n_3278, n_2084, n_4875, n_654, n_411, n_2458, n_1222, n_3050, n_2673, n_2456, n_2527, n_2635, n_1637, n_3307, n_1407, n_1795, n_2871, n_420, n_4321, n_4183, n_164, n_1271, n_4901, n_1545, n_4821, n_4145, n_3121, n_1640, n_4040, n_2406, n_806, n_584, n_2141, n_244, n_548, n_282, n_833, n_523, n_345, n_3930, n_4943, n_799, n_3044, n_4757, n_2196, n_2629, n_2809, n_787, n_2172, n_4682, n_4530, n_1528, n_1146, n_2021, n_4942, n_159, n_1086, n_2125, n_2561, n_652, n_4604, n_1906, n_3305, n_2992, n_1241, n_3157, n_4841, n_1758, n_3221, n_3267, n_2422, n_1914, n_1318, n_4338, n_3457, n_306, n_3762, n_3005, n_3151, n_3411, n_4840, n_1029, n_4519, n_3779, n_2388, n_3984, n_1706, n_1498, n_2417, n_1210, n_5093, n_1556, n_4052, n_3558, n_1984, n_2236, n_4326, n_1269, n_2083, n_2834, n_3207, n_2441, n_3401, n_3242, n_3613, n_655, n_4726, n_1045, n_786, n_1559, n_1872, n_19, n_29, n_75, n_5040, n_1325, n_3761, n_4315, n_2888, n_2923, n_1727, n_4301, n_151, n_3744, n_4788, n_2041, n_1360, n_3814, n_3781, n_1908, n_2484, n_2126, n_3843, n_1098, n_2045, n_817, n_3687, n_2216, n_3543, n_3621, n_2903, n_3216, n_332, n_3808, n_398, n_4365, n_1882, n_3726, n_1007, n_1929, n_2369, n_1592, n_2719, n_591, n_3758, n_2587, n_3199, n_680, n_3339, n_4923, n_2400, n_1953, n_4741, n_3343, n_2752, n_4885, n_751, n_1399, n_4550, n_4652, n_2358, n_3658, n_4900, n_2163, n_2186, n_2815, n_3034, n_4408, n_4577, n_4748, n_643, n_400, n_337, n_2814, n_789, n_3231, n_4212, n_2979, n_181, n_2953, n_327, n_4295, n_2946, n_2500, n_3430, n_2269, n_1729, n_4225, n_300, n_747, n_2565, n_1389, n_535, n_3583, n_3860, n_3851, n_5064, n_3015, n_2175, n_601, n_2182, n_4009, n_1848, n_5002, n_1506, n_119, n_3473, n_1652, n_957, n_1994, n_2566, n_387, n_744, n_971, n_2702, n_3241, n_2906, n_4342, n_4568, n_1205, n_1258, n_2438, n_2914, n_3100, n_2180, n_2858, n_3573, n_1016, n_4106, n_1501, n_3604, n_4373, n_197, n_4711, n_3068, n_2685, n_1083, n_3553, n_2275, n_2465, n_2568, n_2022, n_3811, n_910, n_3494, n_1721, n_1737, n_3486, n_4086, n_752, n_908, n_1028, n_2106, n_2265, n_2032, n_4812, n_4409, n_4629, n_4638, n_708, n_1973, n_3181, n_1500, n_3699, n_854, n_4913, n_2312, n_904, n_709, n_1266, n_2242, n_3328, n_185, n_3868, n_1276, n_4266, n_2466, n_2530, n_1085, n_2042, n_771, n_475, n_924, n_298, n_1582, n_492, n_2318, n_3286, n_4012, n_1149, n_3170, n_265, n_3645, n_5075, n_3682, n_3304, n_2592, n_4968, n_3771, n_2666, n_1585, n_1799, n_2564, n_5085, n_4259, n_2433, n_829, n_2035, n_3422, n_4572, n_859, n_3086, n_2033, n_406, n_4104, n_4845, n_1770, n_878, n_5120, n_130, n_3285, n_4208, n_981, n_4089, n_1144, n_2071, n_3219, n_3702, n_2233, n_4779, n_481, n_3233, n_4599, n_997, n_4437, n_3310, n_1306, n_3264, n_2010, n_1198, n_4061, n_2174, n_436, n_3881, n_4508, n_4727, n_4594, n_2426, n_2478, n_1133, n_95, n_4429, n_4642, n_4051, n_1051, n_4865, n_1039, n_2043, n_1480, n_3206, n_1305, n_2363, n_2578, n_4562, n_553, n_3383, n_4903, n_3709, n_3738, n_4186, n_2540, n_973, n_3610, n_4998, n_3330, n_2065, n_2879, n_967, n_4522, n_2001, n_4341, n_679, n_1629, n_4263, n_225, n_1260, n_1819, n_309, n_3555, n_915, n_812, n_1131, n_3155, n_1006, n_3110, n_1632, n_257, n_1888, n_1311, n_4780, n_670, n_2697, n_3908, n_4973, n_3467, n_1887, n_1587, n_3916, n_3527, n_4803, n_2512, n_3950, n_1242, n_2086, n_2927, n_4750, n_3039, n_1226, n_3740, n_2166, n_2899, n_3186, n_640, n_1322, n_1958, n_315, n_1197, n_3065, n_2632, n_4984, n_2579, n_2105, n_135, n_1423, n_3387, n_364, n_3420, n_5041, n_1915, n_4275, n_4283, n_4959, n_900, n_4426, n_2912, n_60, n_2659, n_4425, n_3409, n_4449, n_2116, n_2320, n_1013, n_1259, n_2183, n_3002, n_51, n_649, n_1612, n_4809, n_1199, n_3392, n_625, n_226, n_68, n_212, n_3773, n_2003, n_1038, n_1581, n_3301, n_1357, n_4241, n_1853, n_798, n_2324, n_245, n_1348, n_2977, n_1739, n_1380, n_2847, n_2557, n_1009, n_62, n_2405, n_4050, n_1160, n_883, n_2647, n_1032, n_2336, n_1247, n_2521, n_1099, n_471, n_424, n_4578, n_2211, n_4777, n_369, n_2672, n_4702, n_2299, n_4179, n_4895, n_141, n_1285, n_1985, n_1172, n_4026, n_71, n_4531, n_3282, n_1590, n_3626, n_1532, n_2313, n_5072, n_3106, n_1140, n_1670, n_2344, n_2365, n_4666, n_3031, n_4029, n_375, n_2447, n_4617, n_2340, n_4010, n_1649, n_4555, n_4969, n_5105, n_1572, n_4308, n_5021, n_3463, n_428, n_2510, n_1954, n_822, n_2791, n_4325, n_3251, n_4602, n_5044, n_5134, n_2212, n_3063, n_1163, n_2729, n_2582, n_1798, n_1550, n_491, n_3998, n_1591, n_3632, n_3122, n_1344, n_2730, n_2495, n_371, n_2090, n_2603, n_538, n_3829, n_4164, n_2173, n_1471, n_4919, n_3737, n_3655, n_493, n_3825, n_2880, n_3225, n_2108, n_5158, n_1211, n_5022, n_1280, n_3296, n_58, n_1445, n_2551, n_1526, n_5047, n_196, n_2985, n_1978, n_574, n_3792, n_4202, n_1446, n_14, n_3938, n_4791, n_3507, n_4403, n_3269, n_3531, n_473, n_1054, n_559, n_1956, n_4139, n_4549, n_1986, n_2397, n_3931, n_4349, n_5141, n_2113, n_1918, n_3603, n_813, n_3822, n_4163, n_818, n_645, n_3812, n_3910, n_2633, n_2207, n_4948, n_2696, n_3482, n_4080, n_2198, n_3319, n_541, n_2073, n_2273, n_3748, n_3272, n_4941, n_2, n_3396, n_4393, n_1162, n_4372, n_821, n_1068, n_982, n_408, n_932, n_2831, n_4318, n_4158, n_3317, n_3978, n_2123, n_1697, n_979, n_4074, n_3716, n_4795, n_4918, n_3824, n_5067, n_4013, n_4544, n_3248, n_354, n_134, n_2941, n_1278, n_547, n_5108, n_4032, n_1064, n_1396, n_634, n_2355, n_4147, n_136, n_4477, n_3168, n_2751, n_4337, n_4130, n_2009, n_1793, n_3601, n_3092, n_1289, n_3055, n_3966, n_2866, n_4742, n_1014, n_3734, n_1703, n_2580, n_882, n_3649, n_2821, n_1875, n_1865, n_3746, n_3384, n_1950, n_1563, n_3419, n_1297, n_1662, n_4478, n_1359, n_2818, n_3794, n_674, n_3921, n_922, n_1335, n_1927, n_4838, n_702, n_4965, n_347, n_3346, n_1896, n_2965, n_3058, n_3861, n_675, n_1540, n_1977, n_3891, n_2193, n_4523, n_1655, n_242, n_1886, n_4371, n_2994, n_3428, n_3153, n_4552, n_3689, n_877, n_4673, n_2519, n_728, n_3415, n_1063, n_4607, n_4041, n_2947, n_3918, n_1965, n_4837, n_2476, n_598, n_437, n_4169, n_697, n_3271, n_295, n_5088, n_4248, n_388, n_484, n_2976, n_2152, n_2652, n_1825, n_1757, n_170, n_1792, n_1412, n_2497, n_3809, n_3139, n_4070, n_3545, n_3885, n_1369, n_881, n_3993, n_4685, n_63, n_4031, n_148, n_4675, n_2663, n_4018, n_2987, n_694, n_2938, n_3780, n_297, n_3337, n_4002, n_3209, n_1044, n_2165, n_1391, n_131, n_2750, n_2775, n_1295, n_3477, n_2349, n_2684, n_3146, n_1495, n_1438, n_3953, n_4588, n_1100, n_585, n_4653, n_4435, n_1756, n_1128, n_673, n_4019, n_1071, n_1968, n_4728, n_4999, n_4385, n_4922, n_865, n_3616, n_4191, n_2870, n_59, n_2151, n_1839, n_2341, n_1765, n_3727, n_2707, n_826, n_4350, n_3747, n_1714, n_104, n_718, n_4330, n_542, n_305, n_2089, n_3522, n_2747, n_3924, n_791, n_4621, n_4216, n_510, n_4240, n_3491, n_1488, n_704, n_2148, n_4162, n_2339, n_2861, n_1999, n_2731, n_622, n_147, n_3353, n_3018, n_3975, n_1838, n_2638, n_4785, n_4683, n_1766, n_1776, n_2002, n_2138, n_4021, n_2414, n_3014, n_1771, n_2316, n_4103, n_5060, n_3148, n_4022, n_4986, n_145, n_2208, n_4775, n_4864, n_4674, n_4481, n_1304, n_294, n_3775, n_4669, n_2134, n_1176, n_425, n_1431, n_3312, n_3835, n_4286, n_2958, n_3731, n_1822, n_2936, n_3224, n_2489, n_1087, n_657, n_2771, n_3020, n_4525, n_1505, n_290, n_3557, n_2610, n_3129, n_3620, n_478, n_107, n_3832, n_2520, n_4484, n_3693, n_446, n_4497, n_1568, n_2372, n_1490, n_526, n_2251, n_3674, n_2959, n_2501, n_3203, n_4871, n_293, n_1070, n_2403, n_2837, n_4700, n_4883, n_1665, n_4306, n_154, n_4224, n_2127, n_3341, n_4453, n_3559, n_4005, n_3546, n_1358, n_3661, n_4564, n_5146, n_3056, n_745, n_2424, n_3201, n_3447, n_3971, n_716, n_1475, n_1774, n_2354, n_3103, n_4573, n_2589, n_4535, n_755, n_527, n_2442, n_3627, n_3480, n_1368, n_1137, n_3612, n_4695, n_2545, n_3509, n_4368, n_2966, n_2294, n_1942, n_1314, n_600, n_3196, n_864, n_2504, n_2623, n_399, n_1440, n_2063, n_1534, n_5005, n_1339, n_2475, n_403, n_723, n_3144, n_3244, n_596, n_1141, n_1268, n_3287, n_3322, n_1755, n_5043, n_2025, n_2357, n_4654, n_3640, n_642, n_995, n_1159, n_3481, n_2250, n_3033, n_303, n_2374, n_416, n_1681, n_520, n_418, n_4597, n_113, n_3364, n_3226, n_2780, n_4020, n_1618, n_4867, n_5061, n_1653, n_4063, n_4237, n_2601, n_5029, n_5127, n_2920, n_773, n_920, n_99, n_1374, n_2648, n_3212, n_13, n_1169, n_1617, n_3370, n_3386, n_335, n_4721, n_463, n_3093, n_848, n_120, n_274, n_4247, n_3169, n_3205, n_1881, n_1267, n_1806, n_2023, n_2204, n_2720, n_496, n_4614, n_177, n_3360, n_2087, n_1636, n_3956, n_4001, n_1323, n_2627, n_4422, n_960, n_778, n_3004, n_3870, n_3625, n_1764, n_4632, n_1610, n_3084, n_2343, n_793, n_4546, n_4583, n_4963, n_3749, n_2942, n_4966, n_4714, n_5037, n_2515, n_316, n_1551, n_4847, n_4054, n_2555, n_3586, n_3653, n_2201, n_725, n_3349, n_4668, n_4635, n_0, n_368, n_994, n_2278, n_1020, n_1273, n_4214, n_3448, n_617, n_2924, n_1036, n_3595, n_1138, n_1661, n_421, n_3991, n_3516, n_3926, n_1095, n_1270, n_4405, n_610, n_4413, n_1852, n_4036, n_4759, n_2153, n_3670, n_2381, n_2052, n_179, n_4667, n_5081, n_517, n_4182, n_667, n_3230, n_1279, n_1115, n_1499, n_504, n_1409, n_1503, n_2819, n_3041, n_4637, n_2423, n_603, n_1657, n_1126, n_2412, n_2439, n_2404, n_1182, n_3635, n_5118, n_4155, n_4238, n_3011, n_2061, n_2757, n_4977, n_167, n_1216, n_2716, n_2452, n_3650, n_3010, n_3043, n_4590, n_2543, n_5090, n_3137, n_2486, n_3560, n_3177, n_4929, n_122, n_2220, n_2577, n_34, n_1262, n_3238, n_218, n_3529, n_70, n_4835, n_2232, n_4038, n_2790, n_4565, n_4159, n_3784, n_220, n_4586, n_1608, n_2373, n_1472, n_3628, n_800, n_4734, n_1491, n_1840, n_4434, n_2244, n_4290, n_2586, n_1684, n_2446, n_1346, n_1352, n_2017, n_3029, n_3597, n_1046, n_2560, n_2704, n_1145, n_1121, n_1102, n_1963, n_258, n_3790, n_2766, n_260, n_356, n_3318, n_4833, n_5062, n_152, n_4888, n_776, n_321, n_1823, n_2479, n_3350, n_2782, n_3977, n_227, n_3588, n_4279, n_5008, n_1456, n_5004, n_23, n_2229, n_4133, n_4527, n_2288, n_2099, n_3388, n_4790, n_1946, n_4181, n_3184, n_4561, n_4461, n_464, n_3245, n_3075, n_4007, n_4949, n_2642, n_4239, n_2383, n_4184, n_1676, n_1830, n_2351, n_1319, n_5069, n_2986, n_2536, n_3915, n_139, n_1633, n_3489, n_2835, n_1416, n_2820, n_2293, n_3074, n_3102, n_2026, n_1282, n_550, n_3321, n_2567, n_2322, n_275, n_2727, n_3377, n_560, n_4782, n_1321, n_2533, n_569, n_3530, n_2869, n_4378, n_1235, n_2759, n_2361, n_1292, n_2266, n_4876, n_346, n_3, n_790, n_2611, n_2901, n_4358, n_2653, n_49, n_299, n_1248, n_902, n_2189, n_2246, n_4469, n_431, n_3156, n_672, n_1941, n_3483, n_706, n_1794, n_1236, n_4493, n_4924, n_743, n_766, n_430, n_1746, n_3524, n_489, n_2885, n_636, n_110, n_3097, n_660, n_2062, n_4539, n_2975, n_4421, n_2839, n_2856, n_4793, n_4498, n_2070, n_1607, n_1454, n_4953, n_2348, n_2944, n_3831, n_869, n_1154, n_646, n_528, n_391, n_1329, n_5167, n_3589, n_262, n_897, n_846, n_2066, n_841, n_1476, n_3391, n_508, n_1800, n_1463, n_3458, n_4505, n_3190, n_1562, n_1826, n_57, n_5126, n_1759, n_5051, n_52, n_853, n_875, n_5012, n_1678, n_661, n_3787, n_1256, n_3585, n_3565, n_4450, n_7, n_5025, n_933, n_4173, n_3135, n_4630, n_1217, n_3990, n_310, n_1628, n_2109, n_988, n_2796, n_2507, n_84, n_4534, n_1536, n_1204, n_1132, n_233, n_1327, n_955, n_246, n_2787, n_2969, n_2395, n_1554, n_4494, n_769, n_2380, n_4786, n_1120, n_555, n_4579, n_669, n_2290, n_4811, n_2048, n_176, n_114, n_2005, n_4857, n_3432, n_2736, n_2883, n_1408, n_4282, n_1196, n_3493, n_863, n_3774, n_2910, n_748, n_3268, n_1785, n_1147, n_1754, n_3057, n_3701, n_5148, n_2584, n_1812, n_866, n_2287, n_452, n_761, n_2492, n_3778, n_174, n_1173, n_4974, n_4911, n_4436, n_5119, n_4569, n_1174, n_3334, n_647, n_5097, n_844, n_17, n_4985, n_2117, n_2234, n_3823, n_4384, n_2741, n_3114, n_888, n_2203, n_2255, n_3584, n_236, n_4858, n_4678, n_2649, n_3556, n_3836, n_414, n_1922, n_4823, n_4309, n_4363, n_1215, n_93, n_839, n_5107, n_3456, n_5095, n_779, n_1537, n_2205, n_4243, n_4025, n_3404, n_1122, n_4059, n_1509, n_4121, n_3290, n_1109, n_4313, n_3309, n_3671, n_4142, n_2015, n_3982, n_2609, n_1161, n_3796, n_232, n_3840, n_46, n_3461, n_3408, n_4246, n_3513, n_3690, n_1184, n_2483, n_4532, n_228, n_1525, n_3995, n_4076, n_2594, n_4244, n_2147, n_592, n_2503, n_4049, n_1156, n_2600, n_984, n_3508, n_132, n_868, n_4353, n_735, n_4787, n_469, n_1218, n_3596, n_4537, n_4346, n_4351, n_357, n_2429, n_985, n_2440, n_3521, n_802, n_561, n_980, n_2681, n_1651, n_2360, n_3764, n_4784, n_4075, n_116, n_3947, n_1244, n_1685, n_3066, n_2844, n_2303, n_1619, n_2285, n_4451, n_4332, n_810, n_1194, n_4538, n_4506, n_2742, n_3695, n_3976, n_3563, n_2367, n_201, n_3198, n_3495, n_1034, n_2909, n_754, n_975, n_43, n_3359, n_467, n_3187, n_3218, n_582, n_861, n_857, n_2107, n_2040, n_2968, n_4201, n_4336, n_2221, n_588, n_4852, n_1010, n_4210, n_4981, n_1166, n_2891, n_2709, n_534, n_1578, n_1861, n_3955, n_1557, n_2280, n_3945, n_730, n_203, n_1898, n_2443, n_4936, n_4205, n_2162, n_1868, n_207, n_2079, n_4763, n_3587, n_4278, n_3433, n_4463, n_205, n_2185, n_1836, n_3833, n_2774, n_3162, n_1274, n_1486, n_3333, n_4129, n_81, n_5032, n_1899, n_784, n_4804, n_3965, n_4500, n_5065, n_862, n_2098, n_3085, n_4433, n_2813, n_1935, n_2027, n_2091, n_2991, n_5030, n_4194, n_1449, n_4703, n_361, n_2419, n_2677, n_3182, n_3283, n_1742, n_4030, n_18607);

input n_2542;
input n_1671;
input n_2817;
input n_801;
input n_4452;
input n_2576;
input n_4649;
input n_1674;
input n_741;
input n_1351;
input n_1212;
input n_208;
input n_4251;
input n_2157;
input n_5019;
input n_2332;
input n_3849;
input n_578;
input n_5138;
input n_4388;
input n_4395;
input n_1061;
input n_3089;
input n_783;
input n_4978;
input n_188;
input n_1854;
input n_3088;
input n_3257;
input n_1342;
input n_4829;
input n_1387;
input n_3222;
input n_677;
input n_4699;
input n_1151;
input n_4686;
input n_2317;
input n_442;
input n_1975;
input n_1930;
input n_3706;
input n_2179;
input n_5055;
input n_1547;
input n_3376;
input n_4868;
input n_893;
input n_3801;
input n_4249;
input n_1192;
input n_3564;
input n_1844;
input n_1555;
input n_5057;
input n_3030;
input n_830;
input n_65;
input n_447;
input n_2838;
input n_3427;
input n_852;
input n_5101;
input n_2628;
input n_3071;
input n_2926;
input n_1078;
input n_544;
input n_4273;
input n_35;
input n_2321;
input n_2019;
input n_5102;
input n_3345;
input n_2074;
input n_2919;
input n_4501;
input n_2129;
input n_4724;
input n_945;
input n_4997;
input n_2399;
input n_4843;
input n_1232;
input n_4696;
input n_4347;
input n_2480;
input n_3877;
input n_3929;
input n_3048;
input n_1455;
input n_2786;
input n_567;
input n_1781;
input n_1971;
input n_2004;
input n_1106;
input n_4814;
input n_953;
input n_3979;
input n_3077;
input n_2873;
input n_3452;
input n_3107;
input n_155;
input n_4956;
input n_454;
input n_1421;
input n_3664;
input n_1936;
input n_5129;
input n_1660;
input n_5070;
input n_3047;
input n_4414;
input n_112;
input n_713;
input n_1400;
input n_2625;
input n_4646;
input n_2843;
input n_3760;
input n_48;
input n_1560;
input n_4262;
input n_734;
input n_1088;
input n_1894;
input n_3347;
input n_5136;
input n_907;
input n_6;
input n_4110;
input n_1658;
input n_4950;
input n_4729;
input n_4268;
input n_1967;
input n_3999;
input n_3928;
input n_2613;
input n_3535;
input n_4751;
input n_44;
input n_2708;
input n_1648;
input n_5151;
input n_1911;
input n_2011;
input n_281;
input n_564;
input n_279;
input n_686;
input n_4102;
input n_1641;
input n_3871;
input n_2735;
input n_4662;
input n_4671;
input n_3959;
input n_2268;
input n_1367;
input n_1336;
input n_4314;
input n_2080;
input n_323;
input n_5099;
input n_1381;
input n_331;
input n_1699;
input n_2093;
input n_4296;
input n_102;
input n_2770;
input n_608;
input n_2101;
input n_4507;
input n_32;
input n_512;
input n_3484;
input n_4677;
input n_792;
input n_5063;
input n_1328;
input n_2917;
input n_2616;
input n_3923;
input n_3900;
input n_3488;
input n_939;
input n_2811;
input n_3732;
input n_2832;
input n_4226;
input n_1762;
input n_1910;
input n_1075;
input n_3980;
input n_2998;
input n_4366;
input n_3446;
input n_237;
input n_1895;
input n_4294;
input n_4698;
input n_4445;
input n_4810;
input n_3859;
input n_2692;
input n_175;
input n_3914;
input n_4456;
input n_3397;
input n_3575;
input n_2469;
input n_3927;
input n_3888;
input n_764;
input n_2764;
input n_2895;
input n_733;
input n_2922;
input n_3882;
input n_4856;
input n_3492;
input n_4369;
input n_30;
input n_2068;
input n_4331;
input n_4972;
input n_1290;
input n_4993;
input n_2072;
input n_1354;
input n_586;
input n_423;
input n_4375;
input n_1701;
input n_2678;
input n_3935;
input n_5130;
input n_4291;
input n_88;
input n_1726;
input n_4613;
input n_2434;
input n_2878;
input n_3012;
input n_3875;
input n_1167;
input n_2428;
input n_4717;
input n_4877;
input n_3247;
input n_871;
input n_210;
input n_2641;
input n_4731;
input n_3052;
input n_178;
input n_355;
input n_5046;
input n_2749;
input n_3298;
input n_2254;
input n_5058;
input n_1926;
input n_3273;
input n_4467;
input n_1747;
input n_195;
input n_780;
input n_2624;
input n_2350;
input n_5042;
input n_4681;
input n_4072;
input n_4752;
input n_4220;
input n_835;
input n_928;
input n_2092;
input n_1654;
input n_1750;
input n_1462;
input n_2514;
input n_604;
input n_1588;
input n_3942;
input n_3997;
input n_26;
input n_2468;
input n_4381;
input n_5144;
input n_515;
input n_2096;
input n_3968;
input n_4466;
input n_4418;
input n_3434;
input n_4510;
input n_4473;
input n_514;
input n_687;
input n_890;
input n_2812;
input n_190;
input n_4518;
input n_1709;
input n_2393;
input n_2657;
input n_2921;
input n_2136;
input n_2409;
input n_2252;
input n_3237;
input n_949;
input n_3500;
input n_3834;
input n_4589;
input n_2075;
input n_2972;
input n_3542;
input n_91;
input n_2763;
input n_2762;
input n_3192;
input n_760;
input n_1546;
input n_4394;
input n_2279;
input n_161;
input n_1296;
input n_3352;
input n_3073;
input n_2150;
input n_1294;
input n_3696;
input n_1420;
input n_4082;
input n_595;
input n_1779;
input n_524;
input n_4921;
input n_1858;
input n_4329;
input n_5135;
input n_3021;
input n_2558;
input n_1164;
input n_4697;
input n_4288;
input n_4289;
input n_3763;
input n_2712;
input n_3733;
input n_1487;
input n_3614;
input n_874;
input n_382;
input n_2145;
input n_898;
input n_4964;
input n_4228;
input n_3423;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_4636;
input n_4322;
input n_3644;
input n_1249;
input n_4946;
input n_2706;
input n_4767;
input n_4287;
input n_2693;
input n_4137;
input n_1127;
input n_1512;
input n_1451;
input n_320;
input n_639;
input n_963;
input n_2767;
input n_4576;
input n_4615;
input n_1139;
input n_3179;
input n_1018;
input n_3400;
input n_1521;
input n_1366;
input n_4000;
input n_2897;
input n_4389;
input n_3970;
input n_4345;
input n_996;
input n_532;
input n_173;
input n_1376;
input n_413;
input n_4664;
input n_2170;
input n_4156;
input n_948;
input n_977;
input n_536;
input n_3158;
input n_1788;
input n_4873;
input n_2643;
input n_3782;
input n_1835;
input n_3470;
input n_5076;
input n_581;
input n_4713;
input n_4098;
input n_5026;
input n_4476;
input n_432;
input n_3700;
input n_4995;
input n_3166;
input n_3104;
input n_3435;
input n_842;
input n_2239;
input n_4310;
input n_1432;
input n_989;
input n_2689;
input n_1473;
input n_2191;
input n_1246;
input n_4528;
input n_899;
input n_1035;
input n_4914;
input n_4939;
input n_499;
input n_1426;
input n_3418;
input n_705;
input n_11;
input n_1004;
input n_1529;
input n_2473;
input n_4634;
input n_2069;
input n_2362;
input n_4096;
input n_2539;
input n_2698;
input n_4123;
input n_3119;
input n_3735;
input n_2297;
input n_4379;
input n_486;
input n_4718;
input n_1448;
input n_3631;
input n_648;
input n_2445;
input n_2057;
input n_2103;
input n_3770;
input n_2772;
input n_4440;
input n_4402;
input n_927;
input n_5052;
input n_4541;
input n_5009;
input n_4872;
input n_929;
input n_4551;
input n_2857;
input n_1183;
input n_4627;
input n_4079;
input n_2494;
input n_3342;
input n_998;
input n_5035;
input n_717;
input n_1383;
input n_3390;
input n_3656;
input n_1424;
input n_1000;
input n_3025;
input n_2137;
input n_1626;
input n_1507;
input n_2482;
input n_3810;
input n_552;
input n_4798;
input n_2532;
input n_1388;
input n_3006;
input n_216;
input n_912;
input n_5010;
input n_2296;
input n_3633;
input n_5089;
input n_2849;
input n_1201;
input n_1398;
input n_884;
input n_4592;
input n_1395;
input n_2199;
input n_2661;
input n_731;
input n_1955;
input n_931;
input n_474;
input n_312;
input n_1791;
input n_66;
input n_958;
input n_5137;
input n_100;
input n_3331;
input n_5104;
input n_1897;
input n_2064;
input n_2773;
input n_589;
input n_3606;
input n_1310;
input n_819;
input n_1334;
input n_3591;
input n_2788;
input n_964;
input n_4756;
input n_2797;
input n_4746;
input n_124;
input n_3892;
input n_4970;
input n_4069;
input n_211;
input n_2748;
input n_1834;
input n_2331;
input n_2292;
input n_3441;
input n_3534;
input n_3964;
input n_2416;
input n_311;
input n_1877;
input n_3944;
input n_1939;
input n_2030;
input n_1769;
input n_556;
input n_2209;
input n_3605;
input n_1602;
input n_4633;
input n_3306;
input n_276;
input n_3026;
input n_221;
input n_4584;
input n_3090;
input n_3724;
input n_4276;
input n_5116;
input n_2990;
input n_3847;
input n_1773;
input n_5001;
input n_2552;
input n_1053;
input n_4428;
input n_1533;
input n_3323;
input n_4;
input n_266;
input n_2274;
input n_518;
input n_4618;
input n_4679;
input n_1745;
input n_914;
input n_3479;
input n_4496;
input n_317;
input n_4805;
input n_1679;
input n_90;
input n_3454;
input n_2160;
input n_2146;
input n_2131;
input n_488;
input n_3547;
input n_2575;
input n_5100;
input n_4410;
input n_1933;
input n_1179;
input n_324;
input n_3816;
input n_4807;
input n_4411;
input n_3214;
input n_1243;
input n_301;
input n_2928;
input n_5166;
input n_1917;
input n_1580;
input n_2822;
input n_36;
input n_4180;
input n_1281;
input n_3109;
input n_3354;
input n_2572;
input n_1520;
input n_3126;
input n_3663;
input n_2863;
input n_1419;
input n_3299;
input n_351;
input n_259;
input n_1731;
input n_2135;
input n_4707;
input n_1645;
input n_1832;
input n_4676;
input n_858;
input n_2049;
input n_956;
input n_663;
input n_4880;
input n_3566;
input n_2781;
input n_4126;
input n_410;
input n_2829;
input n_1696;
input n_3845;
input n_1594;
input n_664;
input n_1869;
input n_3804;
input n_4207;
input n_2016;
input n_4470;
input n_580;
input n_4813;
input n_1030;
input n_3901;
input n_1937;
input n_465;
input n_1790;
input n_4014;
input n_4704;
input n_341;
input n_1744;
input n_828;
input n_2142;
input n_4252;
input n_607;
input n_4028;
input n_2448;
input n_4048;
input n_4596;
input n_4444;
input n_3756;
input n_3406;
input n_820;
input n_951;
input n_952;
input n_3919;
input n_2263;
input n_974;
input n_4952;
input n_2656;
input n_5023;
input n_2375;
input n_1934;
input n_628;
input n_1434;
input n_1573;
input n_3981;
input n_3973;
input n_2756;
input n_807;
input n_4761;
input n_1275;
input n_2884;
input n_485;
input n_67;
input n_1510;
input n_3120;
input n_3797;
input n_238;
input n_2024;
input n_1595;
input n_4770;
input n_202;
input n_1749;
input n_3474;
input n_2549;
input n_4690;
input n_1669;
input n_1024;
input n_3864;
input n_4932;
input n_248;
input n_2302;
input n_1667;
input n_1037;
input n_5143;
input n_3592;
input n_468;
input n_4230;
input n_2637;
input n_1639;
input n_183;
input n_3967;
input n_3195;
input n_466;
input n_2526;
input n_4274;
input n_3277;
input n_2548;
input n_991;
input n_4189;
input n_3817;
input n_340;
input n_1108;
input n_3659;
input n_2559;
input n_2177;
input n_39;
input n_2595;
input n_5003;
input n_4827;
input n_1601;
input n_1960;
input n_2694;
input n_3648;
input n_1686;
input n_3042;
input n_5094;
input n_4610;
input n_4472;
input n_3228;
input n_3657;
input n_96;
input n_3081;
input n_1430;
input n_1316;
input n_1287;
input n_1586;
input n_2264;
input n_3464;
input n_380;
input n_3723;
input n_1190;
input n_397;
input n_4380;
input n_4990;
input n_4996;
input n_4398;
input n_2498;
input n_4515;
input n_1891;
input n_5031;
input n_1213;
input n_2235;
input n_4193;
input n_3570;
input n_5082;
input n_1673;
input n_3828;
input n_172;
input n_2392;
input n_3424;
input n_4131;
input n_239;
input n_97;
input n_2298;
input n_2326;
input n_1539;
input n_490;
input n_3594;
input n_1043;
input n_4090;
input n_4165;
input n_2305;
input n_2120;
input n_80;
input n_4626;
input n_4144;
input n_2964;
input n_352;
input n_2169;
input n_3485;
input n_4077;
input n_2371;
input n_1361;
input n_662;
input n_3262;
input n_4008;
input n_3356;
input n_1642;
input n_3210;
input n_937;
input n_4689;
input n_1682;
input n_4547;
input n_3329;
input n_330;
input n_3826;
input n_4905;
input n_1406;
input n_4601;
input n_962;
input n_3647;
input n_3681;
input n_1883;
input n_4300;
input n_1288;
input n_1186;
input n_4623;
input n_5007;
input n_3320;
input n_2518;
input n_3988;
input n_1720;
input n_3476;
input n_4842;
input n_204;
input n_482;
input n_3439;
input n_4135;
input n_2688;
input n_394;
input n_1845;
input n_1489;
input n_942;
input n_2798;
input n_2852;
input n_1524;
input n_1964;
input n_1920;
input n_2753;
input n_1496;
input n_3292;
input n_2007;
input n_2039;
input n_1225;
input n_1544;
input n_1485;
input n_1846;
input n_3437;
input n_4111;
input n_533;
input n_3712;
input n_4608;
input n_879;
input n_2310;
input n_2506;
input n_4859;
input n_94;
input n_2626;
input n_1567;
input n_4037;
input n_3562;
input n_2973;
input n_41;
input n_3665;
input n_273;
input n_3007;
input n_3528;
input n_4571;
input n_3698;
input n_3355;
input n_2454;
input n_2114;
input n_3174;
input n_1066;
input n_1948;
input n_157;
input n_4215;
input n_2154;
input n_1484;
input n_4185;
input n_3752;
input n_2283;
input n_5145;
input n_4219;
input n_1229;
input n_1373;
input n_3958;
input n_3985;
input n_2427;
input n_4196;
input n_1447;
input n_4774;
input n_2056;
input n_4242;
input n_5109;
input n_3389;
input n_4232;
input n_4190;
input n_4902;
input n_3000;
input n_5149;
input n_2680;
input n_1047;
input n_3375;
input n_3899;
input n_1385;
input n_3713;
input n_1931;
input n_502;
input n_2668;
input n_1257;
input n_3197;
input n_4987;
input n_2128;
input n_4736;
input n_2398;
input n_1725;
input n_3743;
input n_834;
input n_5033;
input n_2695;
input n_4035;
input n_3818;
input n_3124;
input n_1741;
input n_1002;
input n_1949;
input n_3759;
input n_545;
input n_2671;
input n_4516;
input n_2715;
input n_1804;
input n_251;
input n_2508;
input n_3511;
input n_2054;
input n_1337;
input n_1477;
input n_2614;
input n_4492;
input n_2833;
input n_2758;
input n_3694;
input n_2937;
input n_4789;
input n_4376;
input n_1001;
input n_2241;
input n_4708;
input n_4657;
input n_1690;
input n_1191;
input n_1076;
input n_4512;
input n_1378;
input n_855;
input n_1377;
input n_695;
input n_4081;
input n_1542;
input n_4542;
input n_4462;
input n_1716;
input n_278;
input n_4931;
input n_4536;
input n_3303;
input n_978;
input n_4324;
input n_384;
input n_1976;
input n_4382;
input n_2905;
input n_1291;
input n_749;
input n_1824;
input n_3954;
input n_2122;
input n_2140;
input n_3503;
input n_3160;
input n_1065;
input n_1255;
input n_568;
input n_5124;
input n_143;
input n_3951;
input n_823;
input n_1074;
input n_698;
input n_3569;
input n_739;
input n_3874;
input n_2528;
input n_5123;
input n_4639;
input n_1338;
input n_1097;
input n_3027;
input n_781;
input n_4083;
input n_1810;
input n_182;
input n_573;
input n_1583;
input n_4480;
input n_1730;
input n_2295;
input n_2746;
input n_389;
input n_814;
input n_1643;
input n_2020;
input n_4171;
input n_3652;
input n_222;
input n_4023;
input n_1105;
input n_721;
input n_1461;
input n_742;
input n_691;
input n_3617;
input n_2076;
input n_3567;
input n_377;
input n_1598;
input n_4344;
input n_2935;
input n_4705;
input n_4046;
input n_3807;
input n_918;
input n_1114;
input n_56;
input n_763;
input n_4027;
input n_3154;
input n_1227;
input n_2485;
input n_3898;
input n_3520;
input n_191;
input n_4391;
input n_946;
input n_1303;
input n_4095;
input n_2881;
input n_1116;
input n_1570;
input n_1702;
input n_1219;
input n_3551;
input n_4947;
input n_3064;
input n_1780;
input n_3897;
input n_1689;
input n_8;
input n_3372;
input n_1944;
input n_1347;
input n_795;
input n_1221;
input n_1245;
input n_3215;
input n_448;
input n_3853;
input n_4740;
input n_4631;
input n_1561;
input n_1112;
input n_2081;
input n_2168;
input n_5068;
input n_234;
input n_1460;
input n_911;
input n_82;
input n_27;
input n_5159;
input n_2862;
input n_472;
input n_2615;
input n_4068;
input n_4625;
input n_2474;
input n_3703;
input n_2437;
input n_2444;
input n_25;
input n_3962;
input n_2743;
input n_4766;
input n_4863;
input n_2267;
input n_3035;
input n_668;
input n_4166;
input n_1821;
input n_1058;
input n_3378;
input n_3745;
input n_3362;
input n_4744;
input n_103;
input n_4188;
input n_2934;
input n_3667;
input n_3523;
input n_2222;
input n_712;
input n_3176;
input n_31;
input n_2505;
input n_334;
input n_4817;
input n_4115;
input n_2999;
input n_2014;
input n_1239;
input n_3697;
input n_1584;
input n_470;
input n_3680;
input n_2408;
input n_3468;
input n_5045;
input n_1972;
input n_4383;
input n_4491;
input n_455;
input n_363;
input n_4486;
input n_1816;
input n_393;
input n_503;
input n_3024;
input n_4612;
input n_2531;
input n_5163;
input n_307;
input n_4529;
input n_500;
input n_3361;
input n_714;
input n_3478;
input n_3936;
input n_1349;
input n_291;
input n_2723;
input n_2800;
input n_3496;
input n_4390;
input n_3096;
input n_2651;
input n_2095;
input n_3239;
input n_3161;
input n_2799;
input n_3902;
input n_4062;
input n_3295;
input n_4396;
input n_1998;
input n_1574;
input n_3101;
input n_240;
input n_756;
input n_1981;
input n_4233;
input n_1606;
input n_3374;
input n_2640;
input n_253;
input n_1552;
input n_2918;
input n_583;
input n_3288;
input n_4307;
input n_3992;
input n_3876;
input n_249;
input n_3125;
input n_4293;
input n_941;
input n_3552;
input n_1031;
input n_115;
input n_849;
input n_4684;
input n_3116;
input n_4091;
input n_1753;
input n_5027;
input n_3095;
input n_2471;
input n_4412;
input n_2807;
input n_1921;
input n_3618;
input n_4580;
input n_1055;
input n_2217;
input n_2197;
input n_4758;
input n_4781;
input n_4148;
input n_2461;
input n_271;
input n_206;
input n_4057;
input n_633;
input n_1170;
input n_308;
input n_3444;
input n_1040;
input n_3059;
input n_2634;
input n_1761;
input n_1890;
input n_3017;
input n_1805;
input n_2477;
input n_2308;
input n_2333;
input n_3001;
input n_1089;
input n_3795;
input n_3852;
input n_1365;
input n_4138;
input n_5018;
input n_3815;
input n_3896;
input n_3274;
input n_4457;
input n_4093;
input n_1616;
input n_1862;
input n_339;
input n_434;
input n_64;
input n_288;
input n_4928;
input n_4794;
input n_722;
input n_2223;
input n_4197;
input n_4482;
input n_629;
input n_1621;
input n_2547;
input n_2415;
input n_5073;
input n_827;
input n_4834;
input n_4762;
input n_192;
input n_3113;
input n_992;
input n_3813;
input n_3660;
input n_3766;
input n_1613;
input n_1458;
input n_1027;
input n_3266;
input n_3574;
input n_1189;
input n_223;
input n_4154;
input n_4907;
input n_5077;
input n_5034;
input n_726;
input n_50;
input n_4504;
input n_365;
input n_3844;
input n_1237;
input n_2534;
input n_4975;
input n_3741;
input n_2451;
input n_2243;
input n_4815;
input n_4898;
input n_3443;
input n_509;
input n_4819;
input n_1209;
input n_1708;
input n_805;
input n_396;
input n_350;
input n_78;
input n_2051;
input n_4370;
input n_2359;
input n_5112;
input n_480;
input n_142;
input n_1402;
input n_1691;
input n_3332;
input n_4134;
input n_1238;
input n_2570;
input n_4092;
input n_4645;
input n_3668;
input n_2491;
input n_1264;
input n_4755;
input n_4359;
input n_4960;
input n_4087;
input n_1700;
input n_4933;
input n_5091;
input n_3487;
input n_4591;
input n_287;
input n_4302;
input n_5111;
input n_3340;
input n_230;
input n_461;
input n_873;
input n_3946;
input n_2989;
input n_3395;
input n_4474;
input n_2509;
input n_2513;
input n_3757;
input n_4178;
input n_5165;
input n_1704;
input n_2247;
input n_250;
input n_1711;
input n_4884;
input n_1579;
input n_3275;
input n_836;
input n_522;
input n_3678;
input n_3440;
input n_2094;
input n_1511;
input n_2356;
input n_1422;
input n_1772;
input n_4692;
input n_616;
input n_3165;
input n_1119;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2739;
input n_1735;
input n_3890;
input n_1541;
input n_1300;
input n_641;
input n_3750;
input n_1313;
input n_3607;
input n_3316;
input n_516;
input n_2418;
input n_2864;
input n_4311;
input n_1180;
input n_2703;
input n_3371;
input n_4722;
input n_4606;
input n_3261;
input n_666;
input n_4187;
input n_940;
input n_2058;
input n_405;
input n_213;
input n_2660;
input n_1094;
input n_4962;
input n_4563;
input n_494;
input n_5056;
input n_4820;
input n_2394;
input n_3532;
input n_3948;
input n_2124;
input n_4619;
input n_381;
input n_4327;
input n_1961;
input n_3765;
input n_4125;
input n_5036;
input n_4221;
input n_3297;
input n_976;
input n_3067;
input n_2155;
input n_2686;
input n_2364;
input n_4392;
input n_2996;
input n_3803;
input n_2085;
input n_917;
input n_5014;
input n_3639;
input n_4334;
input n_659;
input n_3351;
input n_808;
input n_4047;
input n_3413;
input n_1193;
input n_3412;
input n_3791;
input n_3164;
input n_4575;
input n_551;
input n_699;
input n_4320;
input n_3884;
input n_451;
input n_5139;
input n_757;
input n_594;
input n_2190;
input n_3438;
input n_166;
input n_4141;
input n_2850;
input n_572;
input n_1481;
input n_1441;
input n_3373;
input n_92;
input n_2104;
input n_513;
input n_3883;
input n_261;
input n_3728;
input n_2925;
input n_4499;
input n_121;
input n_433;
input n_3949;
input n_2792;
input n_219;
input n_3315;
input n_263;
input n_3798;
input n_788;
input n_1543;
input n_1599;
input n_329;
input n_4257;
input n_4458;
input n_2674;
input n_5103;
input n_4641;
input n_4720;
input n_4893;
input n_61;
input n_3857;
input n_1876;
input n_4107;
input n_243;
input n_1873;
input n_3630;
input n_3518;
input n_1866;
input n_117;
input n_2130;
input n_1330;
input n_1413;
input n_3714;
input n_2228;
input n_5039;
input n_2455;
input n_2876;
input n_4772;
input n_3099;
input n_4468;
input n_4161;
input n_1663;
input n_4172;
input n_3403;
input n_2714;
input n_2245;
input n_4961;
input n_4454;
input n_1107;
input n_2457;
input n_3294;
input n_4119;
input n_3686;
input n_4502;
input n_318;
input n_2971;
input n_1713;
input n_715;
input n_4277;
input n_4526;
input n_1265;
input n_3490;
input n_4849;
input n_530;
input n_277;
input n_4319;
input n_3369;
input n_618;
input n_199;
input n_3581;
input n_3069;
input n_2028;
input n_3715;
input n_1069;
input n_612;
input n_3725;
input n_3933;
input n_1175;
input n_2311;
input n_429;
input n_1012;
input n_3691;
input n_4485;
input n_4066;
input n_903;
input n_4146;
input n_1802;
input n_1504;
input n_4340;
input n_286;
input n_254;
input n_3961;
input n_4855;
input n_1801;
input n_2347;
input n_3917;
input n_47;
input n_816;
input n_1188;
input n_2206;
input n_4004;
input n_2967;
input n_2916;
input n_4292;
input n_2467;
input n_267;
input n_3145;
input n_1124;
input n_1624;
input n_3983;
input n_4940;
input n_3538;
input n_3280;
input n_1515;
input n_961;
input n_4356;
input n_3510;
input n_2824;
input n_593;
input n_637;
input n_2377;
input n_701;
input n_950;
input n_3009;
input n_3719;
input n_2525;
input n_4361;
input n_3827;
input n_891;
input n_5154;
input n_2067;
input n_3889;
input n_2687;
input n_1630;
input n_2887;
input n_4245;
input n_4136;
input n_3526;
input n_2194;
input n_2619;
input n_4367;
input n_1987;
input n_507;
input n_968;
input n_2271;
input n_1008;
input n_2583;
input n_4560;
input n_2606;
input n_4899;
input n_1033;
input n_462;
input n_1052;
input n_2794;
input n_5164;
input n_2391;
input n_304;
input n_2431;
input n_125;
input n_2078;
input n_2932;
input n_1767;
input n_3431;
input n_3450;
input n_449;
input n_4663;
input n_2893;
input n_1208;
input n_2954;
input n_2728;
input n_1072;
input n_815;
input n_3421;
input n_3183;
input n_2493;
input n_4802;
input n_2705;
input n_1067;
input n_3405;
input n_255;
input n_284;
input n_1952;
input n_5074;
input n_4044;
input n_3436;
input n_1026;
input n_1880;
input n_3442;
input n_3366;
input n_2631;
input n_38;
input n_289;
input n_3937;
input n_1293;
input n_3159;
input n_4701;
input n_108;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_3240;
input n_3576;
input n_1863;
input n_3385;
input n_4851;
input n_3293;
input n_872;
input n_3922;
input n_86;
input n_847;
input n_644;
input n_682;
input n_851;
input n_4991;
input n_72;
input n_2554;
input n_1513;
input n_1913;
input n_4934;
input n_837;
input n_5087;
input n_2517;
input n_2713;
input n_5000;
input n_2765;
input n_2590;
input n_3150;
input n_2060;
input n_4479;
input n_2608;
input n_4011;
input n_5131;
input n_1959;
input n_3133;
input n_765;
input n_1492;
input n_1340;
input n_4688;
input n_4753;
input n_4058;
input n_631;
input n_2262;
input n_3611;
input n_3082;
input n_4848;
input n_5059;
input n_156;
input n_843;
input n_2604;
input n_2407;
input n_1277;
input n_2816;
input n_3799;
input n_2574;
input n_4475;
input n_2675;
input n_3537;
input n_4443;
input n_3887;
input n_1022;
input n_614;
input n_2667;
input n_4587;
input n_1615;
input n_4114;
input n_1474;
input n_1571;
input n_2948;
input n_1577;
input n_2119;
input n_947;
input n_1117;
input n_1992;
input n_3223;
input n_3140;
input n_3185;
input n_4749;
input n_2605;
input n_5155;
input n_118;
input n_926;
input n_3654;
input n_1849;
input n_2848;
input n_919;
input n_1698;
input n_4100;
input n_4264;
input n_3788;
input n_89;
input n_4891;
input n_777;
input n_1299;
input n_3837;
input n_2718;
input n_1436;
input n_1384;
input n_3325;
input n_2238;
input n_4085;
input n_4464;
input n_4624;
input n_4818;
input n_4659;
input n_3600;
input n_18;
input n_5015;
input n_4339;
input n_1178;
input n_98;
input n_2338;
input n_3324;
input n_796;
input n_1195;
input n_184;
input n_1811;
input n_1857;
input n_3987;
input n_1519;
input n_2144;
input n_1284;
input n_1604;
input n_4487;
input n_4889;
input n_4866;
input n_1142;
input n_623;
input n_1048;
input n_3638;
input n_4816;
input n_2110;
input n_1502;
input n_1659;
input n_3393;
input n_3451;
input n_1418;
input n_1250;
input n_292;
input n_4937;
input n_3615;
input n_3072;
input n_3087;
input n_2053;
input n_2259;
input n_2121;
input n_4222;
input n_4874;
input n_4401;
input n_889;
input n_2710;
input n_3142;
input n_4015;
input n_1966;
input n_477;
input n_1110;
input n_4709;
input n_2213;
input n_4976;
input n_2389;
input n_2132;
input n_2892;
input n_4120;
input n_1564;
input n_4658;
input n_231;
input n_2860;
input n_2330;
input n_40;
input n_1457;
input n_505;
input n_3718;
input n_1787;
input n_537;
input n_1993;
input n_2281;
input n_2617;
input n_2776;
input n_1466;
input n_10;
input n_1919;
input n_3705;
input n_3211;
input n_3909;
input n_546;
input n_386;
input n_1220;
input n_1893;
input n_2301;
input n_4665;
input n_3582;
input n_4223;
input n_2387;
input n_3270;
input n_2846;
input n_970;
input n_2488;
input n_1980;
input n_2237;
input n_1060;
input n_1951;
input n_444;
input n_4362;
input n_1252;
input n_3311;
input n_3913;
input n_1223;
input n_511;
input n_5121;
input n_1286;
input n_2115;
input n_4430;
input n_3302;
input n_4348;
input n_5013;
input n_1597;
input n_4489;
input n_4839;
input n_2596;
input n_3163;
input n_775;
input n_4404;
input n_1153;
input n_439;
input n_1531;
input n_2828;
input n_453;
input n_2384;
input n_4261;
input n_4204;
input n_759;
input n_2724;
input n_426;
input n_2585;
input n_4825;
input n_2352;
input n_1625;
input n_3986;
input n_5006;
input n_4513;
input n_4006;
input n_2226;
input n_2801;
input n_1901;
input n_3869;
input n_2556;
input n_4747;
input n_1647;
input n_3753;
input n_2306;
input n_1614;
input n_1892;
input n_3742;
input n_3683;
input n_4801;
input n_401;
input n_3260;
input n_2550;
input n_3175;
input n_3736;
input n_4448;
input n_1096;
input n_2227;
input n_3284;
input n_4869;
input n_427;
input n_2159;
input n_4386;
input n_688;
input n_1077;
input n_2315;
input n_4132;
input n_2995;
input n_1437;
input n_4844;
input n_4438;
input n_4836;
input n_4955;
input n_4149;
input n_4355;
input n_501;
input n_2276;
input n_3234;
input n_856;
input n_2803;
input n_379;
input n_1668;
input n_2777;
input n_3202;
input n_2830;
input n_3220;
input n_1129;
input n_602;
input n_2181;
input n_171;
input n_2911;
input n_169;
input n_4655;
input n_1429;
input n_2826;
input n_3429;
input n_2379;
input n_326;
input n_587;
input n_3554;
input n_1593;
input n_1202;
input n_1635;
input n_4067;
input n_4357;
input n_28;
input n_3462;
input n_2851;
input n_4374;
input n_5132;
input n_106;
input n_358;
input n_160;
input n_2420;
input n_3722;
input n_186;
input n_4400;
input n_4846;
input n_2984;
input n_575;
input n_4024;
input n_1508;
input n_732;
input n_2983;
input n_2240;
input n_392;
input n_2538;
input n_724;
input n_3250;
input n_1042;
input n_4582;
input n_1728;
input n_557;
input n_1871;
input n_4860;
input n_845;
input n_140;
input n_3414;
input n_1549;
input n_4870;
input n_768;
input n_3651;
input n_2102;
input n_2563;
input n_4989;
input n_3449;
input n_1683;
input n_1916;
input n_2598;
input n_597;
input n_280;
input n_1187;
input n_4304;
input n_4558;
input n_1403;
input n_4488;
input n_3767;
input n_2544;
input n_3550;
input n_4211;
input n_1206;
input n_4016;
input n_621;
input n_750;
input n_4656;
input n_3839;
input n_2823;
input n_4915;
input n_4328;
input n_1057;
input n_2785;
input n_235;
input n_1997;
input n_2636;
input n_3131;
input n_710;
input n_1818;
input n_3730;
input n_1298;
input n_4397;
input n_3399;
input n_2088;
input n_1611;
input n_5050;
input n_2740;
input n_746;
input n_4808;
input n_3416;
input n_3498;
input n_2401;
input n_101;
input n_1589;
input n_4712;
input n_2309;
input n_2900;
input n_2957;
input n_1740;
input n_2737;
input n_3994;
input n_1497;
input n_133;
input n_3672;
input n_3533;
input n_1622;
input n_4725;
input n_4406;
input n_1694;
input n_1535;
input n_3382;
input n_3132;
input n_2571;
input n_3138;
input n_20;
input n_5053;
input n_2171;
input n_2988;
input n_4908;
input n_3136;
input n_1350;
input n_4109;
input n_4192;
input n_4824;
input n_2037;
input n_2808;
input n_4567;
input n_5150;
input n_782;
input n_809;
input n_3819;
input n_4778;
input n_1797;
input n_986;
input n_2050;
input n_4595;
input n_2164;
input n_4174;
input n_402;
input n_1870;
input n_1171;
input n_460;
input n_1827;
input n_4904;
input n_2187;
input n_1152;
input n_450;
input n_3544;
input n_4150;
input n_2904;
input n_711;
input n_3105;
input n_2872;
input n_3692;
input n_4616;
input n_4982;
input n_370;
input n_1695;
input n_2046;
input n_2272;
input n_2760;
input n_1979;
input n_4643;
input n_2738;
input n_972;
input n_1332;
input n_4323;
input n_624;
input n_2346;
input n_4831;
input n_936;
input n_3045;
input n_3821;
input n_885;
input n_83;
input n_2342;
input n_2167;
input n_2970;
input n_3676;
input n_4896;
input n_2882;
input n_3666;
input n_3675;
input n_4017;
input n_4260;
input n_4916;
input n_2541;
input n_2940;
input n_4739;
input n_599;
input n_105;
input n_1974;
input n_4122;
input n_934;
input n_4209;
input n_2768;
input n_3858;
input n_1341;
input n_4298;
input n_2314;
input n_3502;
input n_3003;
input n_4128;
input n_543;
input n_5147;
input n_4271;
input n_4644;
input n_1355;
input n_2258;
input n_325;
input n_804;
input n_2390;
input n_959;
input n_2562;
input n_4716;
input n_4312;
input n_1343;
input n_1522;
input n_76;
input n_2734;
input n_1782;
input n_707;
input n_1900;
input n_5048;
input n_3246;
input n_1548;
input n_3381;
input n_1155;
input n_2195;
input n_3208;
input n_4944;
input n_4343;
input n_4715;
input n_4935;
input n_4694;
input n_4672;
input n_5054;
input n_2962;
input n_2939;
input n_1672;
input n_1925;
input n_4407;
input n_737;
input n_4045;
input n_3517;
input n_2945;
input n_4598;
input n_3061;
input n_3893;
input n_3932;
input n_21;
input n_3469;
input n_2960;
input n_138;
input n_3258;
input n_4524;
input n_3143;
input n_333;
input n_4084;
input n_3149;
input n_3365;
input n_3379;
input n_24;
input n_459;
input n_4850;
input n_4424;
input n_3008;
input n_1751;
input n_2840;
input n_285;
input n_3939;
input n_4776;
input n_1375;
input n_3972;
input n_4153;
input n_85;
input n_3506;
input n_1650;
input n_1962;
input n_3855;
input n_1928;
input n_3091;
input n_4317;
input n_4723;
input n_4269;
input n_4088;
input n_3398;
input n_2761;
input n_2793;
input n_3776;
input n_3711;
input n_4235;
input n_1019;
input n_4143;
input n_4170;
input n_729;
input n_876;
input n_774;
input n_3642;
input n_2845;
input n_4650;
input n_438;
input n_4719;
input n_1860;
input n_5016;
input n_1904;
input n_2874;
input n_1200;
input n_2588;
input n_479;
input n_1353;
input n_1777;
input n_4967;
input n_3308;
input n_1113;
input n_1600;
input n_2253;
input n_2366;
input n_4912;
input n_4799;
input n_2261;
input n_4423;
input n_5086;
input n_2210;
input n_4735;
input n_3602;
input n_187;
input n_3300;
input n_2978;
input n_2516;
input n_1050;
input n_1411;
input n_2827;
input n_1177;
input n_3515;
input n_1150;
input n_566;
input n_1023;
input n_2951;
input n_1118;
input n_194;
input n_2949;
input n_1807;
input n_5028;
input n_1814;
input n_1631;
input n_1879;
input n_256;
input n_440;
input n_3806;
input n_2931;
input n_209;
input n_367;
input n_2569;
input n_3866;
input n_671;
input n_4543;
input n_740;
input n_703;
input n_4157;
input n_4229;
input n_3865;
input n_4073;
input n_1324;
input n_3629;
input n_1435;
input n_3920;
input n_969;
input n_4892;
input n_3255;
input n_1401;
input n_1516;
input n_3846;
input n_180;
input n_3512;
input n_2029;
input n_4439;
input n_1394;
input n_1326;
input n_4783;
input n_1379;
input n_214;
input n_935;
input n_4910;
input n_1130;
input n_3083;
input n_676;
input n_832;
input n_3049;
input n_5142;
input n_3830;
input n_3679;
input n_3541;
input n_74;
input n_3117;
input n_4930;
input n_372;
input n_111;
input n_314;
input n_378;
input n_338;
input n_1283;
input n_2385;
input n_4112;
input n_506;
input n_360;
input n_2149;
input n_2396;
input n_4557;
input n_4917;
input n_895;
input n_2450;
input n_3739;
input n_4432;
input n_2284;
input n_4352;
input n_4416;
input n_4593;
input n_344;
input n_2769;
input n_4465;
input n_3622;
input n_5114;
input n_4980;
input n_1392;
input n_4495;
input n_5117;
input n_1924;
input n_525;
input n_2463;
input n_3363;
input n_1677;
input n_611;
input n_3721;
input n_3062;
input n_2679;
input n_5024;
input n_4559;
input n_838;
input n_3969;
input n_129;
input n_3336;
input n_4160;
input n_4231;
input n_2952;
input n_1017;
input n_4256;
input n_2779;
input n_4938;
input n_109;
input n_445;
input n_930;
input n_2620;
input n_5162;
input n_1945;
input n_1656;
input n_2112;
input n_1464;
input n_2430;
input n_653;
input n_1414;
input n_2721;
input n_944;
input n_4335;
input n_2034;
input n_576;
input n_270;
input n_2683;
input n_563;
input n_2744;
input n_1011;
input n_4521;
input n_1566;
input n_626;
input n_990;
input n_3204;
input n_1104;
input n_4920;
input n_498;
input n_870;
input n_1253;
input n_366;
input n_1693;
input n_3256;
input n_348;
input n_3802;
input n_376;
input n_2118;
input n_2111;
input n_390;
input n_2915;
input n_1148;
input n_2188;
input n_1989;
input n_2802;
input n_3643;
input n_2425;
input n_4265;
input n_2950;
input n_719;
input n_3060;
input n_3098;
input n_4105;
input n_1851;
input n_1090;
input n_4861;
input n_4064;
input n_4926;
input n_1518;
input n_1362;
input n_3123;
input n_3380;
input n_1829;
input n_1450;
input n_4828;
input n_1638;
input n_3038;
input n_570;
input n_1789;
input n_620;
input n_519;
input n_2523;
input n_2413;
input n_3769;
input n_1482;
input n_3863;
input n_3669;
input n_3130;
input n_4316;
input n_4640;
input n_5122;
input n_1710;
input n_2161;
input n_1301;
input n_2805;
input n_33;
input n_4769;
input n_2282;
input n_4628;
input n_2047;
input n_1609;
input n_3344;
input n_2334;
input n_5133;
input n_409;
input n_1763;
input n_3989;
input n_2490;
input n_4460;
input n_4108;
input n_635;
input n_3786;
input n_3841;
input n_4254;
input n_1996;
input n_2867;
input n_1442;
input n_2726;
input n_4303;
input n_1158;
input n_2248;
input n_5011;
input n_2662;
input n_4909;
input n_3147;
input n_753;
input n_3925;
input n_3180;
input n_2795;
input n_3472;
input n_5106;
input n_269;
input n_359;
input n_1479;
input n_4768;
input n_1675;
input n_3717;
input n_571;
input n_2215;
input n_404;
input n_158;
input n_1884;
input n_665;
input n_2055;
input n_5156;
input n_2553;
input n_149;
input n_632;
input n_2038;
input n_4447;
input n_4826;
input n_3445;
input n_373;
input n_87;
input n_1833;
input n_3903;
input n_1494;
input n_2325;
input n_1850;
input n_3854;
input n_3235;
input n_1417;
input n_3673;
input n_4281;
input n_681;
input n_4648;
input n_3094;
input n_412;
input n_965;
input n_1428;
input n_1576;
input n_1856;
input n_2077;
input n_1059;
input n_4951;
input n_422;
input n_4957;
input n_3079;
input n_165;
input n_4360;
input n_540;
input n_4039;
input n_457;
input n_3070;
input n_3800;
input n_4566;
input n_3263;
input n_4853;
input n_1748;
input n_3504;
input n_531;
input n_4272;
input n_2930;
input n_1025;
input n_3111;
input n_336;
input n_12;
input n_1885;
input n_3054;
input n_1538;
input n_1240;
input n_1;
input n_4730;
input n_1234;
input n_3254;
input n_3684;
input n_4670;
input n_4882;
input n_4620;
input n_3152;
input n_4738;
input n_3579;
input n_3335;
input n_4177;
input n_3783;
input n_700;
input n_1307;
input n_3178;
input n_4127;
input n_1003;
input n_168;
input n_2353;
input n_4099;
input n_4517;
input n_77;
input n_4168;
input n_1738;
input n_4490;
input n_1575;
input n_1923;
input n_2260;
input n_3952;
input n_3911;
input n_1688;
input n_4285;
input n_3465;
input n_1743;
input n_2997;
input n_1991;
input n_2386;
input n_5161;
input n_1724;
input n_3708;
input n_4078;
input n_3046;
input n_2956;
input n_1553;
input n_3619;
input n_1415;
input n_1370;
input n_1786;
input n_4198;
input n_2382;
input n_3754;
input n_2291;
input n_415;
input n_1371;
input n_383;
input n_2886;
input n_2974;
input n_4213;
input n_200;
input n_2184;
input n_2982;
input n_1803;
input n_4065;
input n_229;
input n_2645;
input n_3904;
input n_1393;
input n_1517;
input n_1867;
input n_2630;
input n_1444;
input n_1603;
input n_2470;
input n_4446;
input n_1263;
input n_4417;
input n_4733;
input n_4764;
input n_1261;
input n_3879;
input n_2286;
input n_4743;
input n_2018;
input n_3080;
input n_1903;
input n_1143;
input n_658;
input n_1874;
input n_2865;
input n_2825;
input n_2013;
input n_2044;
input n_3023;
input n_3232;
input n_693;
input n_1056;
input n_758;
input n_2256;
input n_943;
input n_4060;
input n_5110;
input n_4879;
input n_42;
input n_772;
input n_2806;
input n_770;
input n_3028;
input n_3662;
input n_2981;
input n_3076;
input n_886;
input n_343;
input n_3624;
input n_1345;
input n_1820;
input n_4556;
input n_539;
input n_45;
input n_4117;
input n_4687;
input n_2836;
input n_638;
input n_1404;
input n_2378;
input n_887;
input n_2655;
input n_4600;
input n_126;
input n_1467;
input n_4250;
input n_3906;
input n_224;
input n_4954;
input n_1231;
input n_2599;
input n_3963;
input n_3368;
input n_9;
input n_2370;
input n_2612;
input n_2591;
input n_4881;
input n_1815;
input n_2214;
input n_4253;
input n_407;
input n_913;
input n_2593;
input n_4255;
input n_867;
input n_4071;
input n_3568;
input n_1230;
input n_3850;
input n_1333;
input n_2496;
input n_3313;
input n_4605;
input n_3189;
input n_163;
input n_1644;
input n_2725;
input n_2277;
input n_4691;
input n_1558;
input n_1732;
input n_2300;
input n_3943;
input n_4305;
input n_824;
input n_4297;
input n_2907;
input n_577;
input n_1843;
input n_619;
input n_4227;
input n_521;
input n_2778;
input n_395;
input n_1909;
input n_5020;
input n_606;
input n_1123;
input n_1309;
input n_2961;
input n_916;
input n_3934;
input n_4033;
input n_4415;
input n_483;
input n_1970;
input n_630;
input n_2059;
input n_2669;
input n_4094;
input n_4765;
input n_2546;
input n_3193;
input n_2522;
input n_476;
input n_4364;
input n_1957;
input n_4354;
input n_4732;
input n_3912;
input n_3118;
input n_3720;
input n_1907;
input n_2529;
input n_264;
input n_860;
input n_1530;
input n_4745;
input n_938;
input n_1302;
input n_4581;
input n_549;
input n_4377;
input n_2143;
input n_905;
input n_4792;
input n_1680;
input n_3842;
input n_322;
input n_993;
input n_689;
input n_2031;
input n_4878;
input n_1605;
input n_3514;
input n_4979;
input n_1988;
input n_558;
input n_2654;
input n_3036;
input n_966;
input n_4511;
input n_2908;
input n_3357;
input n_692;
input n_1233;
input n_3895;
input n_487;
input n_241;
input n_4520;
input n_3455;
input n_4118;
input n_4503;
input n_2176;
input n_2459;
input n_1111;
input n_3599;
input n_1251;
input n_2711;
input n_4199;
input n_1912;
input n_4441;
input n_1982;
input n_3872;
input n_3772;
input n_1312;
input n_5038;
input n_268;
input n_1760;
input n_4585;
input n_2664;
input n_5;
input n_1664;
input n_1722;
input n_3022;
input n_247;
input n_1165;
input n_4773;
input n_2008;
input n_2192;
input n_3281;
input n_2345;
input n_328;
input n_1386;
input n_4427;
input n_5113;
input n_3549;
input n_2804;
input n_2453;
input n_2676;
input n_3940;
input n_4822;
input n_1214;
input n_690;
input n_850;
input n_4800;
input n_1157;
input n_3453;
input n_3410;
input n_1752;
input n_1813;
input n_3768;
input n_4958;
input n_2810;
input n_4043;
input n_2319;
input n_825;
input n_3785;
input n_2963;
input n_2602;
input n_55;
input n_3873;
input n_2980;
input n_696;
input n_4886;
input n_1082;
input n_1317;
input n_3227;
input n_2733;
input n_3289;
input n_4055;
input n_2178;
input n_2644;
input n_2036;
input n_3326;
input n_4200;
input n_3460;
input n_2411;
input n_1796;
input n_2082;
input n_3519;
input n_678;
input n_5078;
input n_3707;
input n_283;
input n_3578;
input n_909;
input n_4737;
input n_590;
input n_4925;
input n_4116;
input n_362;
input n_22;
input n_1990;
input n_3805;
input n_2943;
input n_1634;
input n_3252;
input n_627;
input n_3253;
input n_1465;
input n_342;
input n_2622;
input n_2658;
input n_2665;
input n_2133;
input n_1712;
input n_4603;
input n_1523;
input n_1627;
input n_5080;
input n_3128;
input n_1527;
input n_495;
input n_2691;
input n_840;
input n_2913;
input n_4471;
input n_2230;
input n_1969;
input n_2690;
input n_1565;
input n_1493;
input n_2573;
input n_2646;
input n_2535;
input n_1364;
input n_3078;
input n_2436;
input n_615;
input n_3838;
input n_4651;
input n_3941;
input n_3793;
input n_4854;
input n_5071;
input n_3789;
input n_605;
input n_1514;
input n_3037;
input n_1646;
input n_3729;
input n_4994;
input n_2537;
input n_4483;
input n_5168;
input n_4661;
input n_1308;
input n_4988;
input n_3171;
input n_3608;
input n_4540;
input n_2097;
input n_79;
input n_3459;
input n_2853;
input n_1808;
input n_3053;
input n_3358;
input n_3499;
input n_4284;
input n_1005;
input n_1947;
input n_3426;
input n_4971;
input n_1469;
input n_5125;
input n_2650;
input n_987;
input n_720;
input n_153;
input n_3229;
input n_3348;
input n_1707;
input n_656;
input n_797;
input n_2933;
input n_2717;
input n_1723;
input n_1878;
input n_189;
input n_738;
input n_2012;
input n_3497;
input n_5066;
input n_2842;
input n_3580;
input n_2335;
input n_529;
input n_2307;
input n_3704;
input n_684;
input n_1809;
input n_4280;
input n_1181;
input n_37;
input n_3173;
input n_3677;
input n_3996;
input n_1049;
input n_4097;
input n_1666;
input n_803;
input n_4218;
input n_1717;
input n_1817;
input n_2449;
input n_3880;
input n_3685;
input n_2868;
input n_2231;
input n_3609;
input n_1228;
input n_417;
input n_4459;
input n_4545;
input n_272;
input n_2896;
input n_3019;
input n_2639;
input n_3471;
input n_2898;
input n_69;
input n_2368;
input n_53;
input n_458;
input n_4175;
input n_16;
input n_3200;
input n_4771;
input n_3259;
input n_2524;
input n_3167;
input n_2460;
input n_3867;
input n_3593;
input n_4455;
input n_1073;
input n_252;
input n_4514;
input n_3191;
input n_4140;
input n_2481;
input n_3561;
input n_4806;
input n_2682;
input n_3032;
input n_5160;
input n_2877;
input n_5098;
input n_1021;
input n_811;
input n_683;
input n_1207;
input n_5140;
input n_4992;
input n_880;
input n_3505;
input n_3540;
input n_3577;
input n_2432;
input n_150;
input n_1478;
input n_4796;
input n_3598;
input n_4442;
input n_2581;
input n_1363;
input n_3641;
input n_3777;
input n_4203;
input n_767;
input n_1837;
input n_2218;
input n_4533;
input n_831;
input n_3590;
input n_2435;
input n_954;
input n_4419;
input n_1410;
input n_1382;
input n_1736;
input n_4053;
input n_1483;
input n_3848;
input n_1372;
input n_3327;
input n_1719;
input n_319;
input n_2701;
input n_2511;
input n_4167;
input n_1427;
input n_2745;
input n_1080;
input n_123;
input n_562;
input n_2323;
input n_2784;
input n_162;
input n_4431;
input n_2421;
input n_1136;
input n_4387;
input n_2618;
input n_3265;
input n_2464;
input n_128;
input n_1125;
input n_3755;
input n_4042;
input n_5128;
input n_2224;
input n_2329;
input n_1092;
input n_441;
input n_4299;
input n_4890;
input n_146;
input n_1784;
input n_3571;
input n_193;
input n_1775;
input n_2410;
input n_1093;
input n_1783;
input n_2929;
input n_4176;
input n_296;
input n_651;
input n_3407;
input n_217;
input n_1185;
input n_3856;
input n_4236;
input n_3425;
input n_215;
input n_3894;
input n_3127;
input n_1831;
input n_2621;
input n_3623;
input n_5079;
input n_54;
input n_1453;
input n_2502;
input n_3646;
input n_497;
input n_4830;
input n_4706;
input n_1315;
input n_4570;
input n_2754;
input n_1224;
input n_2783;
input n_3188;
input n_1459;
input n_2462;
input n_3243;
input n_1135;
input n_2889;
input n_4034;
input n_4056;
input n_4622;
input n_3960;
input n_1470;
input n_4887;
input n_2732;
input n_4693;
input n_4206;
input n_2249;
input n_1091;
input n_2000;
input n_3862;
input n_4267;
input n_2270;
input n_1425;
input n_5049;
input n_983;
input n_906;
input n_1390;
input n_2289;
input n_1733;
input n_2955;
input n_2158;
input n_4609;
input n_1855;
input n_3051;
input n_3367;
input n_385;
input n_1687;
input n_1439;
input n_2328;
input n_2859;
input n_2202;
input n_1331;
input n_613;
input n_736;
input n_3314;
input n_3525;
input n_2100;
input n_5157;
input n_2993;
input n_4754;
input n_3016;
input n_4647;
input n_1134;
input n_3688;
input n_4003;
input n_554;
input n_1995;
input n_3751;
input n_4894;
input n_4113;
input n_1889;
input n_4760;
input n_435;
input n_1905;
input n_3466;
input n_762;
input n_4983;
input n_1778;
input n_1079;
input n_2139;
input n_419;
input n_5083;
input n_4509;
input n_2875;
input n_1103;
input n_3907;
input n_3338;
input n_144;
input n_4217;
input n_4906;
input n_2219;
input n_1203;
input n_3636;
input n_2327;
input n_999;
input n_1254;
input n_2841;
input n_4897;
input n_3539;
input n_3291;
input n_4399;
input n_2304;
input n_2487;
input n_3276;
input n_2597;
input n_3194;
input n_5084;
input n_3572;
input n_349;
input n_3886;
input n_4710;
input n_4420;
input n_443;
input n_892;
input n_3637;
input n_4574;
input n_1468;
input n_2855;
input n_1859;
input n_2156;
input n_1718;
input n_4234;
input n_4101;
input n_3548;
input n_5017;
input n_1768;
input n_3974;
input n_198;
input n_1847;
input n_3634;
input n_1397;
input n_3236;
input n_901;
input n_2755;
input n_3141;
input n_923;
input n_5096;
input n_1841;
input n_4660;
input n_1623;
input n_1015;
input n_3112;
input n_4797;
input n_3108;
input n_4270;
input n_4151;
input n_4945;
input n_3417;
input n_4124;
input n_73;
input n_785;
input n_5153;
input n_609;
input n_4611;
input n_2337;
input n_1356;
input n_3213;
input n_4333;
input n_127;
input n_3820;
input n_2607;
input n_2890;
input n_1168;
input n_5115;
input n_1943;
input n_3249;
input n_1320;
input n_2722;
input n_1452;
input n_2854;
input n_2499;
input n_4152;
input n_302;
input n_137;
input n_1596;
input n_5092;
input n_1734;
input n_3172;
input n_4832;
input n_2902;
input n_3217;
input n_1983;
input n_1938;
input n_2472;
input n_3394;
input n_1715;
input n_3536;
input n_1443;
input n_1272;
input n_2894;
input n_3957;
input n_3710;
input n_4195;
input n_4554;
input n_3040;
input n_3279;
input n_2402;
input n_2225;
input n_1081;
input n_1692;
input n_1084;
input n_1864;
input n_2006;
input n_3402;
input n_3475;
input n_3501;
input n_374;
input n_1705;
input n_3905;
input n_4680;
input n_3013;
input n_921;
input n_579;
input n_2789;
input n_5152;
input n_2257;
input n_4927;
input n_4258;
input n_1828;
input n_2699;
input n_2200;
input n_650;
input n_1940;
input n_4548;
input n_4862;
input n_1405;
input n_2376;
input n_456;
input n_3878;
input n_2670;
input n_313;
input n_2700;
input n_1041;
input n_565;
input n_3134;
input n_1569;
input n_3115;
input n_1062;
input n_896;
input n_4553;
input n_3278;
input n_2084;
input n_4875;
input n_654;
input n_411;
input n_2458;
input n_1222;
input n_3050;
input n_2673;
input n_2456;
input n_2527;
input n_2635;
input n_1637;
input n_3307;
input n_1407;
input n_1795;
input n_2871;
input n_420;
input n_4321;
input n_4183;
input n_164;
input n_1271;
input n_4901;
input n_1545;
input n_4821;
input n_4145;
input n_3121;
input n_1640;
input n_4040;
input n_2406;
input n_806;
input n_584;
input n_2141;
input n_244;
input n_548;
input n_282;
input n_833;
input n_523;
input n_345;
input n_3930;
input n_4943;
input n_799;
input n_3044;
input n_4757;
input n_2196;
input n_2629;
input n_2809;
input n_787;
input n_2172;
input n_4682;
input n_4530;
input n_1528;
input n_1146;
input n_2021;
input n_4942;
input n_159;
input n_1086;
input n_2125;
input n_2561;
input n_652;
input n_4604;
input n_1906;
input n_3305;
input n_2992;
input n_1241;
input n_3157;
input n_4841;
input n_1758;
input n_3221;
input n_3267;
input n_2422;
input n_1914;
input n_1318;
input n_4338;
input n_3457;
input n_306;
input n_3762;
input n_3005;
input n_3151;
input n_3411;
input n_4840;
input n_1029;
input n_4519;
input n_3779;
input n_2388;
input n_3984;
input n_1706;
input n_1498;
input n_2417;
input n_1210;
input n_5093;
input n_1556;
input n_4052;
input n_3558;
input n_1984;
input n_2236;
input n_4326;
input n_1269;
input n_2083;
input n_2834;
input n_3207;
input n_2441;
input n_3401;
input n_3242;
input n_3613;
input n_655;
input n_4726;
input n_1045;
input n_786;
input n_1559;
input n_1872;
input n_19;
input n_29;
input n_75;
input n_5040;
input n_1325;
input n_3761;
input n_4315;
input n_2888;
input n_2923;
input n_1727;
input n_4301;
input n_151;
input n_3744;
input n_4788;
input n_2041;
input n_1360;
input n_3814;
input n_3781;
input n_1908;
input n_2484;
input n_2126;
input n_3843;
input n_1098;
input n_2045;
input n_817;
input n_3687;
input n_2216;
input n_3543;
input n_3621;
input n_2903;
input n_3216;
input n_332;
input n_3808;
input n_398;
input n_4365;
input n_1882;
input n_3726;
input n_1007;
input n_1929;
input n_2369;
input n_1592;
input n_2719;
input n_591;
input n_3758;
input n_2587;
input n_3199;
input n_680;
input n_3339;
input n_4923;
input n_2400;
input n_1953;
input n_4741;
input n_3343;
input n_2752;
input n_4885;
input n_751;
input n_1399;
input n_4550;
input n_4652;
input n_2358;
input n_3658;
input n_4900;
input n_2163;
input n_2186;
input n_2815;
input n_3034;
input n_4408;
input n_4577;
input n_4748;
input n_643;
input n_400;
input n_337;
input n_2814;
input n_789;
input n_3231;
input n_4212;
input n_2979;
input n_181;
input n_2953;
input n_327;
input n_4295;
input n_2946;
input n_2500;
input n_3430;
input n_2269;
input n_1729;
input n_4225;
input n_300;
input n_747;
input n_2565;
input n_1389;
input n_535;
input n_3583;
input n_3860;
input n_3851;
input n_5064;
input n_3015;
input n_2175;
input n_601;
input n_2182;
input n_4009;
input n_1848;
input n_5002;
input n_1506;
input n_119;
input n_3473;
input n_1652;
input n_957;
input n_1994;
input n_2566;
input n_387;
input n_744;
input n_971;
input n_2702;
input n_3241;
input n_2906;
input n_4342;
input n_4568;
input n_1205;
input n_1258;
input n_2438;
input n_2914;
input n_3100;
input n_2180;
input n_2858;
input n_3573;
input n_1016;
input n_4106;
input n_1501;
input n_3604;
input n_4373;
input n_197;
input n_4711;
input n_3068;
input n_2685;
input n_1083;
input n_3553;
input n_2275;
input n_2465;
input n_2568;
input n_2022;
input n_3811;
input n_910;
input n_3494;
input n_1721;
input n_1737;
input n_3486;
input n_4086;
input n_752;
input n_908;
input n_1028;
input n_2106;
input n_2265;
input n_2032;
input n_4812;
input n_4409;
input n_4629;
input n_4638;
input n_708;
input n_1973;
input n_3181;
input n_1500;
input n_3699;
input n_854;
input n_4913;
input n_2312;
input n_904;
input n_709;
input n_1266;
input n_2242;
input n_3328;
input n_185;
input n_3868;
input n_1276;
input n_4266;
input n_2466;
input n_2530;
input n_1085;
input n_2042;
input n_771;
input n_475;
input n_924;
input n_298;
input n_1582;
input n_492;
input n_2318;
input n_3286;
input n_4012;
input n_1149;
input n_3170;
input n_265;
input n_3645;
input n_5075;
input n_3682;
input n_3304;
input n_2592;
input n_4968;
input n_3771;
input n_2666;
input n_1585;
input n_1799;
input n_2564;
input n_5085;
input n_4259;
input n_2433;
input n_829;
input n_2035;
input n_3422;
input n_4572;
input n_859;
input n_3086;
input n_2033;
input n_406;
input n_4104;
input n_4845;
input n_1770;
input n_878;
input n_5120;
input n_130;
input n_3285;
input n_4208;
input n_981;
input n_4089;
input n_1144;
input n_2071;
input n_3219;
input n_3702;
input n_2233;
input n_4779;
input n_481;
input n_3233;
input n_4599;
input n_997;
input n_4437;
input n_3310;
input n_1306;
input n_3264;
input n_2010;
input n_1198;
input n_4061;
input n_2174;
input n_436;
input n_3881;
input n_4508;
input n_4727;
input n_4594;
input n_2426;
input n_2478;
input n_1133;
input n_95;
input n_4429;
input n_4642;
input n_4051;
input n_1051;
input n_4865;
input n_1039;
input n_2043;
input n_1480;
input n_3206;
input n_1305;
input n_2363;
input n_2578;
input n_4562;
input n_553;
input n_3383;
input n_4903;
input n_3709;
input n_3738;
input n_4186;
input n_2540;
input n_973;
input n_3610;
input n_4998;
input n_3330;
input n_2065;
input n_2879;
input n_967;
input n_4522;
input n_2001;
input n_4341;
input n_679;
input n_1629;
input n_4263;
input n_225;
input n_1260;
input n_1819;
input n_309;
input n_3555;
input n_915;
input n_812;
input n_1131;
input n_3155;
input n_1006;
input n_3110;
input n_1632;
input n_257;
input n_1888;
input n_1311;
input n_4780;
input n_670;
input n_2697;
input n_3908;
input n_4973;
input n_3467;
input n_1887;
input n_1587;
input n_3916;
input n_3527;
input n_4803;
input n_2512;
input n_3950;
input n_1242;
input n_2086;
input n_2927;
input n_4750;
input n_3039;
input n_1226;
input n_3740;
input n_2166;
input n_2899;
input n_3186;
input n_640;
input n_1322;
input n_1958;
input n_315;
input n_1197;
input n_3065;
input n_2632;
input n_4984;
input n_2579;
input n_2105;
input n_135;
input n_1423;
input n_3387;
input n_364;
input n_3420;
input n_5041;
input n_1915;
input n_4275;
input n_4283;
input n_4959;
input n_900;
input n_4426;
input n_2912;
input n_60;
input n_2659;
input n_4425;
input n_3409;
input n_4449;
input n_2116;
input n_2320;
input n_1013;
input n_1259;
input n_2183;
input n_3002;
input n_51;
input n_649;
input n_1612;
input n_4809;
input n_1199;
input n_3392;
input n_625;
input n_226;
input n_68;
input n_212;
input n_3773;
input n_2003;
input n_1038;
input n_1581;
input n_3301;
input n_1357;
input n_4241;
input n_1853;
input n_798;
input n_2324;
input n_245;
input n_1348;
input n_2977;
input n_1739;
input n_1380;
input n_2847;
input n_2557;
input n_1009;
input n_62;
input n_2405;
input n_4050;
input n_1160;
input n_883;
input n_2647;
input n_1032;
input n_2336;
input n_1247;
input n_2521;
input n_1099;
input n_471;
input n_424;
input n_4578;
input n_2211;
input n_4777;
input n_369;
input n_2672;
input n_4702;
input n_2299;
input n_4179;
input n_4895;
input n_141;
input n_1285;
input n_1985;
input n_1172;
input n_4026;
input n_71;
input n_4531;
input n_3282;
input n_1590;
input n_3626;
input n_1532;
input n_2313;
input n_5072;
input n_3106;
input n_1140;
input n_1670;
input n_2344;
input n_2365;
input n_4666;
input n_3031;
input n_4029;
input n_375;
input n_2447;
input n_4617;
input n_2340;
input n_4010;
input n_1649;
input n_4555;
input n_4969;
input n_5105;
input n_1572;
input n_4308;
input n_5021;
input n_3463;
input n_428;
input n_2510;
input n_1954;
input n_822;
input n_2791;
input n_4325;
input n_3251;
input n_4602;
input n_5044;
input n_5134;
input n_2212;
input n_3063;
input n_1163;
input n_2729;
input n_2582;
input n_1798;
input n_1550;
input n_491;
input n_3998;
input n_1591;
input n_3632;
input n_3122;
input n_1344;
input n_2730;
input n_2495;
input n_371;
input n_2090;
input n_2603;
input n_538;
input n_3829;
input n_4164;
input n_2173;
input n_1471;
input n_4919;
input n_3737;
input n_3655;
input n_493;
input n_3825;
input n_2880;
input n_3225;
input n_2108;
input n_5158;
input n_1211;
input n_5022;
input n_1280;
input n_3296;
input n_58;
input n_1445;
input n_2551;
input n_1526;
input n_5047;
input n_196;
input n_2985;
input n_1978;
input n_574;
input n_3792;
input n_4202;
input n_1446;
input n_14;
input n_3938;
input n_4791;
input n_3507;
input n_4403;
input n_3269;
input n_3531;
input n_473;
input n_1054;
input n_559;
input n_1956;
input n_4139;
input n_4549;
input n_1986;
input n_2397;
input n_3931;
input n_4349;
input n_5141;
input n_2113;
input n_1918;
input n_3603;
input n_813;
input n_3822;
input n_4163;
input n_818;
input n_645;
input n_3812;
input n_3910;
input n_2633;
input n_2207;
input n_4948;
input n_2696;
input n_3482;
input n_4080;
input n_2198;
input n_3319;
input n_541;
input n_2073;
input n_2273;
input n_3748;
input n_3272;
input n_4941;
input n_2;
input n_3396;
input n_4393;
input n_1162;
input n_4372;
input n_821;
input n_1068;
input n_982;
input n_408;
input n_932;
input n_2831;
input n_4318;
input n_4158;
input n_3317;
input n_3978;
input n_2123;
input n_1697;
input n_979;
input n_4074;
input n_3716;
input n_4795;
input n_4918;
input n_3824;
input n_5067;
input n_4013;
input n_4544;
input n_3248;
input n_354;
input n_134;
input n_2941;
input n_1278;
input n_547;
input n_5108;
input n_4032;
input n_1064;
input n_1396;
input n_634;
input n_2355;
input n_4147;
input n_136;
input n_4477;
input n_3168;
input n_2751;
input n_4337;
input n_4130;
input n_2009;
input n_1793;
input n_3601;
input n_3092;
input n_1289;
input n_3055;
input n_3966;
input n_2866;
input n_4742;
input n_1014;
input n_3734;
input n_1703;
input n_2580;
input n_882;
input n_3649;
input n_2821;
input n_1875;
input n_1865;
input n_3746;
input n_3384;
input n_1950;
input n_1563;
input n_3419;
input n_1297;
input n_1662;
input n_4478;
input n_1359;
input n_2818;
input n_3794;
input n_674;
input n_3921;
input n_922;
input n_1335;
input n_1927;
input n_4838;
input n_702;
input n_4965;
input n_347;
input n_3346;
input n_1896;
input n_2965;
input n_3058;
input n_3861;
input n_675;
input n_1540;
input n_1977;
input n_3891;
input n_2193;
input n_4523;
input n_1655;
input n_242;
input n_1886;
input n_4371;
input n_2994;
input n_3428;
input n_3153;
input n_4552;
input n_3689;
input n_877;
input n_4673;
input n_2519;
input n_728;
input n_3415;
input n_1063;
input n_4607;
input n_4041;
input n_2947;
input n_3918;
input n_1965;
input n_4837;
input n_2476;
input n_598;
input n_437;
input n_4169;
input n_697;
input n_3271;
input n_295;
input n_5088;
input n_4248;
input n_388;
input n_484;
input n_2976;
input n_2152;
input n_2652;
input n_1825;
input n_1757;
input n_170;
input n_1792;
input n_1412;
input n_2497;
input n_3809;
input n_3139;
input n_4070;
input n_3545;
input n_3885;
input n_1369;
input n_881;
input n_3993;
input n_4685;
input n_63;
input n_4031;
input n_148;
input n_4675;
input n_2663;
input n_4018;
input n_2987;
input n_694;
input n_2938;
input n_3780;
input n_297;
input n_3337;
input n_4002;
input n_3209;
input n_1044;
input n_2165;
input n_1391;
input n_131;
input n_2750;
input n_2775;
input n_1295;
input n_3477;
input n_2349;
input n_2684;
input n_3146;
input n_1495;
input n_1438;
input n_3953;
input n_4588;
input n_1100;
input n_585;
input n_4653;
input n_4435;
input n_1756;
input n_1128;
input n_673;
input n_4019;
input n_1071;
input n_1968;
input n_4728;
input n_4999;
input n_4385;
input n_4922;
input n_865;
input n_3616;
input n_4191;
input n_2870;
input n_59;
input n_2151;
input n_1839;
input n_2341;
input n_1765;
input n_3727;
input n_2707;
input n_826;
input n_4350;
input n_3747;
input n_1714;
input n_104;
input n_718;
input n_4330;
input n_542;
input n_305;
input n_2089;
input n_3522;
input n_2747;
input n_3924;
input n_791;
input n_4621;
input n_4216;
input n_510;
input n_4240;
input n_3491;
input n_1488;
input n_704;
input n_2148;
input n_4162;
input n_2339;
input n_2861;
input n_1999;
input n_2731;
input n_622;
input n_147;
input n_3353;
input n_3018;
input n_3975;
input n_1838;
input n_2638;
input n_4785;
input n_4683;
input n_1766;
input n_1776;
input n_2002;
input n_2138;
input n_4021;
input n_2414;
input n_3014;
input n_1771;
input n_2316;
input n_4103;
input n_5060;
input n_3148;
input n_4022;
input n_4986;
input n_145;
input n_2208;
input n_4775;
input n_4864;
input n_4674;
input n_4481;
input n_1304;
input n_294;
input n_3775;
input n_4669;
input n_2134;
input n_1176;
input n_425;
input n_1431;
input n_3312;
input n_3835;
input n_4286;
input n_2958;
input n_3731;
input n_1822;
input n_2936;
input n_3224;
input n_2489;
input n_1087;
input n_657;
input n_2771;
input n_3020;
input n_4525;
input n_1505;
input n_290;
input n_3557;
input n_2610;
input n_3129;
input n_3620;
input n_478;
input n_107;
input n_3832;
input n_2520;
input n_4484;
input n_3693;
input n_446;
input n_4497;
input n_1568;
input n_2372;
input n_1490;
input n_526;
input n_2251;
input n_3674;
input n_2959;
input n_2501;
input n_3203;
input n_4871;
input n_293;
input n_1070;
input n_2403;
input n_2837;
input n_4700;
input n_4883;
input n_1665;
input n_4306;
input n_154;
input n_4224;
input n_2127;
input n_3341;
input n_4453;
input n_3559;
input n_4005;
input n_3546;
input n_1358;
input n_3661;
input n_4564;
input n_5146;
input n_3056;
input n_745;
input n_2424;
input n_3201;
input n_3447;
input n_3971;
input n_716;
input n_1475;
input n_1774;
input n_2354;
input n_3103;
input n_4573;
input n_2589;
input n_4535;
input n_755;
input n_527;
input n_2442;
input n_3627;
input n_3480;
input n_1368;
input n_1137;
input n_3612;
input n_4695;
input n_2545;
input n_3509;
input n_4368;
input n_2966;
input n_2294;
input n_1942;
input n_1314;
input n_600;
input n_3196;
input n_864;
input n_2504;
input n_2623;
input n_399;
input n_1440;
input n_2063;
input n_1534;
input n_5005;
input n_1339;
input n_2475;
input n_403;
input n_723;
input n_3144;
input n_3244;
input n_596;
input n_1141;
input n_1268;
input n_3287;
input n_3322;
input n_1755;
input n_5043;
input n_2025;
input n_2357;
input n_4654;
input n_3640;
input n_642;
input n_995;
input n_1159;
input n_3481;
input n_2250;
input n_3033;
input n_303;
input n_2374;
input n_416;
input n_1681;
input n_520;
input n_418;
input n_4597;
input n_113;
input n_3364;
input n_3226;
input n_2780;
input n_4020;
input n_1618;
input n_4867;
input n_5061;
input n_1653;
input n_4063;
input n_4237;
input n_2601;
input n_5029;
input n_5127;
input n_2920;
input n_773;
input n_920;
input n_99;
input n_1374;
input n_2648;
input n_3212;
input n_13;
input n_1169;
input n_1617;
input n_3370;
input n_3386;
input n_335;
input n_4721;
input n_463;
input n_3093;
input n_848;
input n_120;
input n_274;
input n_4247;
input n_3169;
input n_3205;
input n_1881;
input n_1267;
input n_1806;
input n_2023;
input n_2204;
input n_2720;
input n_496;
input n_4614;
input n_177;
input n_3360;
input n_2087;
input n_1636;
input n_3956;
input n_4001;
input n_1323;
input n_2627;
input n_4422;
input n_960;
input n_778;
input n_3004;
input n_3870;
input n_3625;
input n_1764;
input n_4632;
input n_1610;
input n_3084;
input n_2343;
input n_793;
input n_4546;
input n_4583;
input n_4963;
input n_3749;
input n_2942;
input n_4966;
input n_4714;
input n_5037;
input n_2515;
input n_316;
input n_1551;
input n_4847;
input n_4054;
input n_2555;
input n_3586;
input n_3653;
input n_2201;
input n_725;
input n_3349;
input n_4668;
input n_4635;
input n_0;
input n_368;
input n_994;
input n_2278;
input n_1020;
input n_1273;
input n_4214;
input n_3448;
input n_617;
input n_2924;
input n_1036;
input n_3595;
input n_1138;
input n_1661;
input n_421;
input n_3991;
input n_3516;
input n_3926;
input n_1095;
input n_1270;
input n_4405;
input n_610;
input n_4413;
input n_1852;
input n_4036;
input n_4759;
input n_2153;
input n_3670;
input n_2381;
input n_2052;
input n_179;
input n_4667;
input n_5081;
input n_517;
input n_4182;
input n_667;
input n_3230;
input n_1279;
input n_1115;
input n_1499;
input n_504;
input n_1409;
input n_1503;
input n_2819;
input n_3041;
input n_4637;
input n_2423;
input n_603;
input n_1657;
input n_1126;
input n_2412;
input n_2439;
input n_2404;
input n_1182;
input n_3635;
input n_5118;
input n_4155;
input n_4238;
input n_3011;
input n_2061;
input n_2757;
input n_4977;
input n_167;
input n_1216;
input n_2716;
input n_2452;
input n_3650;
input n_3010;
input n_3043;
input n_4590;
input n_2543;
input n_5090;
input n_3137;
input n_2486;
input n_3560;
input n_3177;
input n_4929;
input n_122;
input n_2220;
input n_2577;
input n_34;
input n_1262;
input n_3238;
input n_218;
input n_3529;
input n_70;
input n_4835;
input n_2232;
input n_4038;
input n_2790;
input n_4565;
input n_4159;
input n_3784;
input n_220;
input n_4586;
input n_1608;
input n_2373;
input n_1472;
input n_3628;
input n_800;
input n_4734;
input n_1491;
input n_1840;
input n_4434;
input n_2244;
input n_4290;
input n_2586;
input n_1684;
input n_2446;
input n_1346;
input n_1352;
input n_2017;
input n_3029;
input n_3597;
input n_1046;
input n_2560;
input n_2704;
input n_1145;
input n_1121;
input n_1102;
input n_1963;
input n_258;
input n_3790;
input n_2766;
input n_260;
input n_356;
input n_3318;
input n_4833;
input n_5062;
input n_152;
input n_4888;
input n_776;
input n_321;
input n_1823;
input n_2479;
input n_3350;
input n_2782;
input n_3977;
input n_227;
input n_3588;
input n_4279;
input n_5008;
input n_1456;
input n_5004;
input n_23;
input n_2229;
input n_4133;
input n_4527;
input n_2288;
input n_2099;
input n_3388;
input n_4790;
input n_1946;
input n_4181;
input n_3184;
input n_4561;
input n_4461;
input n_464;
input n_3245;
input n_3075;
input n_4007;
input n_4949;
input n_2642;
input n_4239;
input n_2383;
input n_4184;
input n_1676;
input n_1830;
input n_2351;
input n_1319;
input n_5069;
input n_2986;
input n_2536;
input n_3915;
input n_139;
input n_1633;
input n_3489;
input n_2835;
input n_1416;
input n_2820;
input n_2293;
input n_3074;
input n_3102;
input n_2026;
input n_1282;
input n_550;
input n_3321;
input n_2567;
input n_2322;
input n_275;
input n_2727;
input n_3377;
input n_560;
input n_4782;
input n_1321;
input n_2533;
input n_569;
input n_3530;
input n_2869;
input n_4378;
input n_1235;
input n_2759;
input n_2361;
input n_1292;
input n_2266;
input n_4876;
input n_346;
input n_3;
input n_790;
input n_2611;
input n_2901;
input n_4358;
input n_2653;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_2189;
input n_2246;
input n_4469;
input n_431;
input n_3156;
input n_672;
input n_1941;
input n_3483;
input n_706;
input n_1794;
input n_1236;
input n_4493;
input n_4924;
input n_743;
input n_766;
input n_430;
input n_1746;
input n_3524;
input n_489;
input n_2885;
input n_636;
input n_110;
input n_3097;
input n_660;
input n_2062;
input n_4539;
input n_2975;
input n_4421;
input n_2839;
input n_2856;
input n_4793;
input n_4498;
input n_2070;
input n_1607;
input n_1454;
input n_4953;
input n_2348;
input n_2944;
input n_3831;
input n_869;
input n_1154;
input n_646;
input n_528;
input n_391;
input n_1329;
input n_5167;
input n_3589;
input n_262;
input n_897;
input n_846;
input n_2066;
input n_841;
input n_1476;
input n_3391;
input n_508;
input n_1800;
input n_1463;
input n_3458;
input n_4505;
input n_3190;
input n_1562;
input n_1826;
input n_57;
input n_5126;
input n_1759;
input n_5051;
input n_52;
input n_853;
input n_875;
input n_5012;
input n_1678;
input n_661;
input n_3787;
input n_1256;
input n_3585;
input n_3565;
input n_4450;
input n_7;
input n_5025;
input n_933;
input n_4173;
input n_3135;
input n_4630;
input n_1217;
input n_3990;
input n_310;
input n_1628;
input n_2109;
input n_988;
input n_2796;
input n_2507;
input n_84;
input n_4534;
input n_1536;
input n_1204;
input n_1132;
input n_233;
input n_1327;
input n_955;
input n_246;
input n_2787;
input n_2969;
input n_2395;
input n_1554;
input n_4494;
input n_769;
input n_2380;
input n_4786;
input n_1120;
input n_555;
input n_4579;
input n_669;
input n_2290;
input n_4811;
input n_2048;
input n_176;
input n_114;
input n_2005;
input n_4857;
input n_3432;
input n_2736;
input n_2883;
input n_1408;
input n_4282;
input n_1196;
input n_3493;
input n_863;
input n_3774;
input n_2910;
input n_748;
input n_3268;
input n_1785;
input n_1147;
input n_1754;
input n_3057;
input n_3701;
input n_5148;
input n_2584;
input n_1812;
input n_866;
input n_2287;
input n_452;
input n_761;
input n_2492;
input n_3778;
input n_174;
input n_1173;
input n_4974;
input n_4911;
input n_4436;
input n_5119;
input n_4569;
input n_1174;
input n_3334;
input n_647;
input n_5097;
input n_844;
input n_17;
input n_4985;
input n_2117;
input n_2234;
input n_3823;
input n_4384;
input n_2741;
input n_3114;
input n_888;
input n_2203;
input n_2255;
input n_3584;
input n_236;
input n_4858;
input n_4678;
input n_2649;
input n_3556;
input n_3836;
input n_414;
input n_1922;
input n_4823;
input n_4309;
input n_4363;
input n_1215;
input n_93;
input n_839;
input n_5107;
input n_3456;
input n_5095;
input n_779;
input n_1537;
input n_2205;
input n_4243;
input n_4025;
input n_3404;
input n_1122;
input n_4059;
input n_1509;
input n_4121;
input n_3290;
input n_1109;
input n_4313;
input n_3309;
input n_3671;
input n_4142;
input n_2015;
input n_3982;
input n_2609;
input n_1161;
input n_3796;
input n_232;
input n_3840;
input n_46;
input n_3461;
input n_3408;
input n_4246;
input n_3513;
input n_3690;
input n_1184;
input n_2483;
input n_4532;
input n_228;
input n_1525;
input n_3995;
input n_4076;
input n_2594;
input n_4244;
input n_2147;
input n_592;
input n_2503;
input n_4049;
input n_1156;
input n_2600;
input n_984;
input n_3508;
input n_132;
input n_868;
input n_4353;
input n_735;
input n_4787;
input n_469;
input n_1218;
input n_3596;
input n_4537;
input n_4346;
input n_4351;
input n_357;
input n_2429;
input n_985;
input n_2440;
input n_3521;
input n_802;
input n_561;
input n_980;
input n_2681;
input n_1651;
input n_2360;
input n_3764;
input n_4784;
input n_4075;
input n_116;
input n_3947;
input n_1244;
input n_1685;
input n_3066;
input n_2844;
input n_2303;
input n_1619;
input n_2285;
input n_4451;
input n_4332;
input n_810;
input n_1194;
input n_4538;
input n_4506;
input n_2742;
input n_3695;
input n_3976;
input n_3563;
input n_2367;
input n_201;
input n_3198;
input n_3495;
input n_1034;
input n_2909;
input n_754;
input n_975;
input n_43;
input n_3359;
input n_467;
input n_3187;
input n_3218;
input n_582;
input n_861;
input n_857;
input n_2107;
input n_2040;
input n_2968;
input n_4201;
input n_4336;
input n_2221;
input n_588;
input n_4852;
input n_1010;
input n_4210;
input n_4981;
input n_1166;
input n_2891;
input n_2709;
input n_534;
input n_1578;
input n_1861;
input n_3955;
input n_1557;
input n_2280;
input n_3945;
input n_730;
input n_203;
input n_1898;
input n_2443;
input n_4936;
input n_4205;
input n_2162;
input n_1868;
input n_207;
input n_2079;
input n_4763;
input n_3587;
input n_4278;
input n_3433;
input n_4463;
input n_205;
input n_2185;
input n_1836;
input n_3833;
input n_2774;
input n_3162;
input n_1274;
input n_1486;
input n_3333;
input n_4129;
input n_81;
input n_5032;
input n_1899;
input n_784;
input n_4804;
input n_3965;
input n_4500;
input n_5065;
input n_862;
input n_2098;
input n_3085;
input n_4433;
input n_2813;
input n_1935;
input n_2027;
input n_2091;
input n_2991;
input n_5030;
input n_4194;
input n_1449;
input n_4703;
input n_361;
input n_2419;
input n_2677;
input n_3182;
input n_3283;
input n_1742;
input n_4030;

output n_18607;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_14428;
wire n_13611;
wire n_15214;
wire n_18318;
wire n_6566;
wire n_13045;
wire n_5172;
wire n_11173;
wire n_15268;
wire n_16218;
wire n_5315;
wire n_10487;
wire n_6872;
wire n_16664;
wire n_13998;
wire n_5254;
wire n_17347;
wire n_11926;
wire n_17825;
wire n_6441;
wire n_8668;
wire n_6806;
wire n_5362;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_10587;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_18540;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_13522;
wire n_10931;
wire n_6960;
wire n_15609;
wire n_8169;
wire n_12265;
wire n_9002;
wire n_16423;
wire n_16335;
wire n_14670;
wire n_9130;
wire n_7180;
wire n_5653;
wire n_11574;
wire n_13530;
wire n_8604;
wire n_15049;
wire n_16362;
wire n_5409;
wire n_5301;
wire n_17777;
wire n_7263;
wire n_13125;
wire n_15181;
wire n_8168;
wire n_7190;
wire n_7504;
wire n_8186;
wire n_5393;
wire n_6725;
wire n_6126;
wire n_12322;
wire n_14318;
wire n_17647;
wire n_8899;
wire n_14196;
wire n_15971;
wire n_5524;
wire n_10236;
wire n_17673;
wire n_5345;
wire n_11678;
wire n_11205;
wire n_11776;
wire n_17634;
wire n_17004;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_11650;
wire n_5818;
wire n_16307;
wire n_8005;
wire n_8130;
wire n_8534;
wire n_5963;
wire n_16911;
wire n_12179;
wire n_13942;
wire n_15294;
wire n_14439;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_18230;
wire n_11905;
wire n_10020;
wire n_14825;
wire n_16288;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_11536;
wire n_5950;
wire n_15295;
wire n_9104;
wire n_14914;
wire n_6999;
wire n_14741;
wire n_17050;
wire n_17992;
wire n_17991;
wire n_15665;
wire n_11046;
wire n_11079;
wire n_10283;
wire n_5548;
wire n_17408;
wire n_17735;
wire n_15581;
wire n_11065;
wire n_15445;
wire n_8339;
wire n_8272;
wire n_17624;
wire n_14215;
wire n_13997;
wire n_14402;
wire n_7161;
wire n_7868;
wire n_14882;
wire n_5838;
wire n_15764;
wire n_5725;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_16696;
wire n_17368;
wire n_11214;
wire n_18105;
wire n_7000;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_7398;
wire n_18335;
wire n_14341;
wire n_10392;
wire n_14232;
wire n_12882;
wire n_5900;
wire n_18057;
wire n_15074;
wire n_5545;
wire n_18104;
wire n_12617;
wire n_8411;
wire n_8499;
wire n_8236;
wire n_15253;
wire n_15356;
wire n_13137;
wire n_16733;
wire n_13221;
wire n_18525;
wire n_6882;
wire n_9626;
wire n_10775;
wire n_11163;
wire n_15933;
wire n_9526;
wire n_13657;
wire n_17188;
wire n_15571;
wire n_17511;
wire n_6325;
wire n_9840;
wire n_14099;
wire n_5598;
wire n_15632;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_15898;
wire n_18013;
wire n_16245;
wire n_7389;
wire n_10719;
wire n_11419;
wire n_9018;
wire n_12095;
wire n_8070;
wire n_13663;
wire n_13990;
wire n_16302;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_14939;
wire n_11740;
wire n_17471;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_17138;
wire n_17700;
wire n_10015;
wire n_13993;
wire n_16786;
wire n_18468;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_17227;
wire n_5819;
wire n_17118;
wire n_7008;
wire n_12392;
wire n_15353;
wire n_8366;
wire n_8102;
wire n_9362;
wire n_11979;
wire n_7516;
wire n_7401;
wire n_7596;
wire n_18087;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_15993;
wire n_18090;
wire n_5894;
wire n_16095;
wire n_18502;
wire n_10759;
wire n_17699;
wire n_8022;
wire n_17226;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_18211;
wire n_9658;
wire n_5239;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_17546;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_15797;
wire n_9962;
wire n_17279;
wire n_5908;
wire n_10373;
wire n_18183;
wire n_11104;
wire n_8913;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_11537;
wire n_16772;
wire n_14699;
wire n_13814;
wire n_12707;
wire n_14861;
wire n_7686;
wire n_6914;
wire n_10335;
wire n_5337;
wire n_15194;
wire n_15362;
wire n_11301;
wire n_12424;
wire n_13681;
wire n_14121;
wire n_15101;
wire n_5420;
wire n_15572;
wire n_17209;
wire n_10381;
wire n_18154;
wire n_6243;
wire n_6585;
wire n_11703;
wire n_16553;
wire n_11699;
wire n_18122;
wire n_6374;
wire n_7651;
wire n_11543;
wire n_17013;
wire n_10947;
wire n_6628;
wire n_16984;
wire n_8125;
wire n_13483;
wire n_6015;
wire n_14662;
wire n_11261;
wire n_14811;
wire n_17608;
wire n_10226;
wire n_16012;
wire n_13247;
wire n_16286;
wire n_6526;
wire n_13929;
wire n_16551;
wire n_7956;
wire n_17401;
wire n_17803;
wire n_7369;
wire n_6570;
wire n_16549;
wire n_8556;
wire n_7196;
wire n_10767;
wire n_15421;
wire n_17739;
wire n_8040;
wire n_14646;
wire n_15964;
wire n_11821;
wire n_14095;
wire n_5638;
wire n_13121;
wire n_13989;
wire n_9100;
wire n_14864;
wire n_15069;
wire n_6784;
wire n_17936;
wire n_16643;
wire n_12107;
wire n_14520;
wire n_10755;
wire n_14780;
wire n_18310;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_16998;
wire n_11447;
wire n_6323;
wire n_17847;
wire n_9614;
wire n_14431;
wire n_15200;
wire n_17349;
wire n_13515;
wire n_10682;
wire n_6110;
wire n_17478;
wire n_11684;
wire n_12652;
wire n_16024;
wire n_16324;
wire n_6371;
wire n_14410;
wire n_8079;
wire n_10699;
wire n_15507;
wire n_7846;
wire n_8595;
wire n_15800;
wire n_9400;
wire n_18352;
wire n_8142;
wire n_11627;
wire n_5684;
wire n_8598;
wire n_13139;
wire n_15887;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_13803;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_16078;
wire n_14066;
wire n_7856;
wire n_7774;
wire n_15600;
wire n_16267;
wire n_6674;
wire n_5680;
wire n_17883;
wire n_13606;
wire n_6951;
wire n_6148;
wire n_11659;
wire n_15899;
wire n_7625;
wire n_13501;
wire n_18317;
wire n_9106;
wire n_13509;
wire n_12775;
wire n_17637;
wire n_13729;
wire n_8869;
wire n_6989;
wire n_7863;
wire n_8381;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14813;
wire n_9520;
wire n_17149;
wire n_14791;
wire n_8958;
wire n_14485;
wire n_14931;
wire n_18002;
wire n_12833;
wire n_12090;
wire n_6896;
wire n_14628;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_13687;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_16268;
wire n_12371;
wire n_10114;
wire n_17854;
wire n_12203;
wire n_10357;
wire n_14540;
wire n_15762;
wire n_16784;
wire n_7147;
wire n_8115;
wire n_16351;
wire n_15883;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_11497;
wire n_14900;
wire n_17706;
wire n_15320;
wire n_12359;
wire n_12915;
wire n_6196;
wire n_9037;
wire n_15983;
wire n_13149;
wire n_13711;
wire n_15846;
wire n_13454;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_16721;
wire n_15874;
wire n_12742;
wire n_16662;
wire n_14091;
wire n_9042;
wire n_15755;
wire n_11768;
wire n_8412;
wire n_9267;
wire n_17329;
wire n_6485;
wire n_14478;
wire n_8987;
wire n_11805;
wire n_14461;
wire n_17848;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_16689;
wire n_5493;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_13958;
wire n_17619;
wire n_14935;
wire n_15332;
wire n_5346;
wire n_5252;
wire n_5309;
wire n_18445;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_12770;
wire n_10012;
wire n_14570;
wire n_15986;
wire n_16068;
wire n_13754;
wire n_12985;
wire n_13797;
wire n_13013;
wire n_13238;
wire n_7564;
wire n_11635;
wire n_16254;
wire n_14989;
wire n_15434;
wire n_16530;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_14171;
wire n_16191;
wire n_10204;
wire n_17564;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_8119;
wire n_10296;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_15212;
wire n_15977;
wire n_17136;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_9128;
wire n_10281;
wire n_13344;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_14380;
wire n_16004;
wire n_8748;
wire n_13984;
wire n_17766;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_14239;
wire n_6794;
wire n_6151;
wire n_15896;
wire n_16843;
wire n_8718;
wire n_7110;
wire n_5476;
wire n_17273;
wire n_12831;
wire n_13920;
wire n_9935;
wire n_6431;
wire n_18119;
wire n_6990;
wire n_8659;
wire n_14045;
wire n_14288;
wire n_14824;
wire n_10097;
wire n_8223;
wire n_15767;
wire n_18604;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_15635;
wire n_10018;
wire n_7297;
wire n_9866;
wire n_15183;
wire n_16509;
wire n_16800;
wire n_7298;
wire n_15118;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_12427;
wire n_7533;
wire n_14162;
wire n_13771;
wire n_7221;
wire n_13977;
wire n_10656;
wire n_15159;
wire n_16026;
wire n_6575;
wire n_8727;
wire n_6055;
wire n_8224;
wire n_11295;
wire n_18494;
wire n_16538;
wire n_11662;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_8952;
wire n_8246;
wire n_15679;
wire n_13014;
wire n_16992;
wire n_9070;
wire n_18065;
wire n_11708;
wire n_10266;
wire n_15629;
wire n_14401;
wire n_17949;
wire n_5609;
wire n_17721;
wire n_10897;
wire n_10827;
wire n_5922;
wire n_15154;
wire n_14922;
wire n_10449;
wire n_7569;
wire n_7861;
wire n_7734;
wire n_7062;
wire n_7823;
wire n_8955;
wire n_9477;
wire n_5658;
wire n_9680;
wire n_12172;
wire n_12147;
wire n_12923;
wire n_14769;
wire n_7039;
wire n_17781;
wire n_8577;
wire n_12384;
wire n_14961;
wire n_11349;
wire n_8594;
wire n_13227;
wire n_8428;
wire n_9829;
wire n_15438;
wire n_11260;
wire n_8848;
wire n_12825;
wire n_13341;
wire n_10685;
wire n_11351;
wire n_17139;
wire n_15185;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_14803;
wire n_5667;
wire n_8259;
wire n_12540;
wire n_15611;
wire n_10607;
wire n_14388;
wire n_16035;
wire n_15490;
wire n_5865;
wire n_15182;
wire n_12249;
wire n_8349;
wire n_18033;
wire n_6836;
wire n_5305;
wire n_14977;
wire n_11998;
wire n_8164;
wire n_13239;
wire n_10628;
wire n_13429;
wire n_15942;
wire n_5281;
wire n_7905;
wire n_8776;
wire n_11775;
wire n_15100;
wire n_9143;
wire n_8287;
wire n_10256;
wire n_7753;
wire n_10769;
wire n_6771;
wire n_10368;
wire n_14732;
wire n_7950;
wire n_9947;
wire n_16659;
wire n_13999;
wire n_9088;
wire n_8607;
wire n_14037;
wire n_10138;
wire n_12117;
wire n_17032;
wire n_11706;
wire n_6248;
wire n_16768;
wire n_11800;
wire n_16134;
wire n_10183;
wire n_10375;
wire n_18382;
wire n_17161;
wire n_6952;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_10452;
wire n_11464;
wire n_7806;
wire n_12960;
wire n_14878;
wire n_14094;
wire n_15928;
wire n_13033;
wire n_11642;
wire n_15046;
wire n_11143;
wire n_15703;
wire n_16092;
wire n_7595;
wire n_10383;
wire n_7648;
wire n_17103;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_16352;
wire n_12131;
wire n_6776;
wire n_12851;
wire n_5795;
wire n_18032;
wire n_11934;
wire n_12349;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_14282;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_6714;
wire n_15518;
wire n_11308;
wire n_13550;
wire n_16266;
wire n_17601;
wire n_14217;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_13348;
wire n_8416;
wire n_10396;
wire n_13919;
wire n_10724;
wire n_13642;
wire n_16398;
wire n_17596;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_15574;
wire n_11084;
wire n_14062;
wire n_9988;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_14167;
wire n_12740;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_15872;
wire n_10363;
wire n_13240;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_11553;
wire n_12578;
wire n_12795;
wire n_10517;
wire n_16889;
wire n_17580;
wire n_10323;
wire n_12194;
wire n_13623;
wire n_10842;
wire n_17620;
wire n_7519;
wire n_16465;
wire n_7400;
wire n_10876;
wire n_11511;
wire n_15833;
wire n_9137;
wire n_15649;
wire n_11180;
wire n_14043;
wire n_9724;
wire n_11146;
wire n_16046;
wire n_9281;
wire n_10883;
wire n_8995;
wire n_10101;
wire n_15863;
wire n_9393;
wire n_15974;
wire n_6581;
wire n_13845;
wire n_17785;
wire n_12709;
wire n_6010;
wire n_13432;
wire n_8711;
wire n_7013;
wire n_12771;
wire n_14150;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_18602;
wire n_7290;
wire n_12278;
wire n_13721;
wire n_17760;
wire n_18430;
wire n_10820;
wire n_13514;
wire n_9687;
wire n_17672;
wire n_14787;
wire n_18036;
wire n_7303;
wire n_17414;
wire n_6616;
wire n_8306;
wire n_17100;
wire n_10123;
wire n_10781;
wire n_18052;
wire n_7488;
wire n_7315;
wire n_13194;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_13244;
wire n_16183;
wire n_11866;
wire n_6185;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_5529;
wire n_15659;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_9102;
wire n_17191;
wire n_11526;
wire n_17483;
wire n_13404;
wire n_9578;
wire n_16115;
wire n_17689;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_14785;
wire n_7438;
wire n_17857;
wire n_16631;
wire n_14355;
wire n_14128;
wire n_7268;
wire n_7337;
wire n_11851;
wire n_17323;
wire n_9489;
wire n_12804;
wire n_14123;
wire n_6965;
wire n_5957;
wire n_12116;
wire n_10728;
wire n_6357;
wire n_10094;
wire n_9144;
wire n_6800;
wire n_10084;
wire n_10468;
wire n_14105;
wire n_14126;
wire n_18191;
wire n_7461;
wire n_8285;
wire n_13870;
wire n_10655;
wire n_13791;
wire n_9797;
wire n_15133;
wire n_6955;
wire n_8483;
wire n_16885;
wire n_9521;
wire n_17696;
wire n_15288;
wire n_8332;
wire n_9478;
wire n_9932;
wire n_13040;
wire n_7278;
wire n_11370;
wire n_6509;
wire n_13900;
wire n_16224;
wire n_16731;
wire n_7454;
wire n_11253;
wire n_14652;
wire n_17102;
wire n_11379;
wire n_15527;
wire n_16627;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_17443;
wire n_5787;
wire n_11981;
wire n_16146;
wire n_16654;
wire n_9895;
wire n_8741;
wire n_12918;
wire n_9351;
wire n_11585;
wire n_16452;
wire n_5445;
wire n_18332;
wire n_13140;
wire n_13962;
wire n_14556;
wire n_5501;
wire n_6839;
wire n_5342;
wire n_7377;
wire n_7232;
wire n_13753;
wire n_18145;
wire n_16132;
wire n_6646;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_9189;
wire n_16991;
wire n_18051;
wire n_15149;
wire n_16528;
wire n_15365;
wire n_13716;
wire n_17141;
wire n_14844;
wire n_16907;
wire n_14701;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_14391;
wire n_7904;
wire n_11691;
wire n_16587;
wire n_18171;
wire n_6033;
wire n_11541;
wire n_15495;
wire n_13610;
wire n_8851;
wire n_8921;
wire n_9410;
wire n_9801;
wire n_13332;
wire n_5748;
wire n_14408;
wire n_15293;
wire n_9356;
wire n_15880;
wire n_12865;
wire n_16499;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_8394;
wire n_11155;
wire n_5870;
wire n_18328;
wire n_9175;
wire n_7093;
wire n_6508;
wire n_7168;
wire n_17604;
wire n_12013;
wire n_11835;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_5636;
wire n_7840;
wire n_10972;
wire n_6359;
wire n_7782;
wire n_13213;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_8800;
wire n_16386;
wire n_17101;
wire n_13385;
wire n_15695;
wire n_10845;
wire n_7080;
wire n_17984;
wire n_6636;
wire n_5286;
wire n_8229;
wire n_17643;
wire n_16339;
wire n_8410;
wire n_14756;
wire n_14863;
wire n_5811;
wire n_14156;
wire n_13992;
wire n_17429;
wire n_18144;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_7624;
wire n_7629;
wire n_13790;
wire n_14384;
wire n_9735;
wire n_16185;
wire n_9186;
wire n_10818;
wire n_5530;
wire n_15905;
wire n_5397;
wire n_10624;
wire n_12552;
wire n_13304;
wire n_14633;
wire n_11069;
wire n_15178;
wire n_5595;
wire n_9941;
wire n_12222;
wire n_11951;
wire n_7003;
wire n_15699;
wire n_11900;
wire n_17131;
wire n_14711;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_17163;
wire n_11369;
wire n_10563;
wire n_14210;
wire n_8810;
wire n_5388;
wire n_9802;
wire n_15788;
wire n_5901;
wire n_13362;
wire n_6538;
wire n_14373;
wire n_5962;
wire n_7010;
wire n_5599;
wire n_8107;
wire n_11108;
wire n_12992;
wire n_9728;
wire n_12883;
wire n_11004;
wire n_16690;
wire n_5324;
wire n_6519;
wire n_15752;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_9818;
wire n_6530;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_15694;
wire n_8774;
wire n_14518;
wire n_16310;
wire n_10566;
wire n_17798;
wire n_16503;
wire n_16477;
wire n_13397;
wire n_16568;
wire n_10178;
wire n_17581;
wire n_7299;
wire n_12367;
wire n_17360;
wire n_12104;
wire n_17731;
wire n_15360;
wire n_17954;
wire n_6402;
wire n_12469;
wire n_13526;
wire n_9936;
wire n_12563;
wire n_15829;
wire n_6195;
wire n_18070;
wire n_13132;
wire n_7243;
wire n_7326;
wire n_9530;
wire n_6609;
wire n_10115;
wire n_13321;
wire n_17522;
wire n_14692;
wire n_15042;
wire n_17157;
wire n_5326;
wire n_7471;
wire n_16927;
wire n_7067;
wire n_10455;
wire n_11778;
wire n_12793;
wire n_14722;
wire n_13427;
wire n_15519;
wire n_15488;
wire n_14835;
wire n_5300;
wire n_15391;
wire n_9909;
wire n_11393;
wire n_14871;
wire n_16226;
wire n_8691;
wire n_8620;
wire n_12406;
wire n_14907;
wire n_6748;
wire n_15264;
wire n_7741;
wire n_9466;
wire n_13270;
wire n_16525;
wire n_7790;
wire n_11719;
wire n_16315;
wire n_6149;
wire n_16685;
wire n_10052;
wire n_17918;
wire n_10109;
wire n_18151;
wire n_7484;
wire n_7002;
wire n_16979;
wire n_16639;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_18282;
wire n_16239;
wire n_15358;
wire n_11963;
wire n_12428;
wire n_14636;
wire n_8424;
wire n_9571;
wire n_16334;
wire n_15814;
wire n_8026;
wire n_9638;
wire n_7528;
wire n_9470;
wire n_16003;
wire n_16069;
wire n_15516;
wire n_10265;
wire n_8174;
wire n_12655;
wire n_16676;
wire n_7941;
wire n_13524;
wire n_16096;
wire n_11175;
wire n_13792;
wire n_15756;
wire n_11483;
wire n_5352;
wire n_15067;
wire n_11995;
wire n_14378;
wire n_13356;
wire n_17897;
wire n_11371;
wire n_18299;
wire n_14912;
wire n_10040;
wire n_5394;
wire n_18229;
wire n_9405;
wire n_6264;
wire n_14191;
wire n_16546;
wire n_8861;
wire n_18252;
wire n_5359;
wire n_13480;
wire n_8644;
wire n_17426;
wire n_17454;
wire n_8907;
wire n_16144;
wire n_16669;
wire n_12304;
wire n_13571;
wire n_15156;
wire n_11080;
wire n_10984;
wire n_6902;
wire n_14079;
wire n_10100;
wire n_15168;
wire n_17557;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_15411;
wire n_15743;
wire n_18490;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7478;
wire n_7913;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_15144;
wire n_13600;
wire n_12692;
wire n_13715;
wire n_7939;
wire n_13602;
wire n_14224;
wire n_17436;
wire n_8503;
wire n_16675;
wire n_9612;
wire n_16785;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_16062;
wire n_14919;
wire n_6449;
wire n_17712;
wire n_7458;
wire n_6723;
wire n_9108;
wire n_16653;
wire n_16692;
wire n_9787;
wire n_7436;
wire n_6440;
wire n_10846;
wire n_13363;
wire n_15186;
wire n_16935;
wire n_14101;
wire n_6461;
wire n_18273;
wire n_9376;
wire n_8446;
wire n_9786;
wire n_5194;
wire n_14682;
wire n_14908;
wire n_18576;
wire n_9033;
wire n_13810;
wire n_14403;
wire n_12933;
wire n_7435;
wire n_12908;
wire n_15031;
wire n_15718;
wire n_9537;
wire n_17654;
wire n_11297;
wire n_14635;
wire n_6997;
wire n_10509;
wire n_17076;
wire n_5952;
wire n_13893;
wire n_17168;
wire n_12996;
wire n_15171;
wire n_14201;
wire n_5947;
wire n_8923;
wire n_13625;
wire n_12643;
wire n_13315;
wire n_13473;
wire n_6736;
wire n_7685;
wire n_6124;
wire n_7363;
wire n_8192;
wire n_14597;
wire n_5985;
wire n_8197;
wire n_18267;
wire n_15663;
wire n_14353;
wire n_15963;
wire n_16589;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_14950;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_12827;
wire n_12678;
wire n_13795;
wire n_9115;
wire n_17501;
wire n_12235;
wire n_14547;
wire n_15416;
wire n_5232;
wire n_11833;
wire n_7663;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_14386;
wire n_15868;
wire n_17249;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_16472;
wire n_17830;
wire n_9938;
wire n_11285;
wire n_8082;
wire n_12098;
wire n_8730;
wire n_7917;
wire n_7261;
wire n_15533;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_9203;
wire n_14415;
wire n_9977;
wire n_15073;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_15165;
wire n_5761;
wire n_13982;
wire n_13475;
wire n_16298;
wire n_9242;
wire n_15079;
wire n_6773;
wire n_12611;
wire n_13859;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_13569;
wire n_17040;
wire n_11262;
wire n_7968;
wire n_7455;
wire n_6382;
wire n_12713;
wire n_12880;
wire n_13144;
wire n_18042;
wire n_18542;
wire n_8651;
wire n_18129;
wire n_13959;
wire n_9141;
wire n_15867;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_6531;
wire n_10952;
wire n_10851;
wire n_11027;
wire n_13628;
wire n_11852;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_10221;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_11803;
wire n_15738;
wire n_18560;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_13685;
wire n_16749;
wire n_9286;
wire n_16301;
wire n_8015;
wire n_18507;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_8281;
wire n_10819;
wire n_14693;
wire n_15613;
wire n_8842;
wire n_14786;
wire n_14521;
wire n_9184;
wire n_9704;
wire n_16915;
wire n_13585;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_18418;
wire n_18472;
wire n_14486;
wire n_8024;
wire n_12562;
wire n_7730;
wire n_8814;
wire n_18396;
wire n_8530;
wire n_11428;
wire n_17553;
wire n_11592;
wire n_15090;
wire n_16531;
wire n_17626;
wire n_9193;
wire n_11677;
wire n_8467;
wire n_17043;
wire n_7281;
wire n_16882;
wire n_15385;
wire n_9717;
wire n_13577;
wire n_7711;
wire n_16094;
wire n_16181;
wire n_11090;
wire n_15948;
wire n_8984;
wire n_17123;
wire n_18523;
wire n_5688;
wire n_6417;
wire n_9290;
wire n_13281;
wire n_5740;
wire n_5820;
wire n_13769;
wire n_5648;
wire n_14870;
wire n_13266;
wire n_13957;
wire n_14580;
wire n_15627;
wire n_5745;
wire n_9403;
wire n_10996;
wire n_13672;
wire n_14028;
wire n_9875;
wire n_5180;
wire n_17600;
wire n_6763;
wire n_8956;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_14772;
wire n_8676;
wire n_5534;
wire n_8003;
wire n_13827;
wire n_8785;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_17170;
wire n_6542;
wire n_15681;
wire n_14542;
wire n_17826;
wire n_6556;
wire n_15048;
wire n_8692;
wire n_6889;
wire n_7230;
wire n_9183;
wire n_16142;
wire n_7989;
wire n_17135;
wire n_17552;
wire n_9778;
wire n_14326;
wire n_5196;
wire n_6199;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_15739;
wire n_16381;
wire n_16891;
wire n_18280;
wire n_18118;
wire n_10852;
wire n_15003;
wire n_14665;
wire n_6726;
wire n_12374;
wire n_13200;
wire n_9529;
wire n_5542;
wire n_7011;
wire n_8998;
wire n_10538;
wire n_16783;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_13342;
wire n_11066;
wire n_10315;
wire n_17327;
wire n_18321;
wire n_13886;
wire n_16887;
wire n_9123;
wire n_17374;
wire n_17187;
wire n_6576;
wire n_6471;
wire n_17031;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_15545;
wire n_14924;
wire n_12368;
wire n_17117;
wire n_5255;
wire n_8482;
wire n_17240;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_18477;
wire n_13193;
wire n_6100;
wire n_12796;
wire n_16242;
wire n_6516;
wire n_14489;
wire n_16053;
wire n_8462;
wire n_17845;
wire n_13774;
wire n_6977;
wire n_16854;
wire n_9380;
wire n_13847;
wire n_10062;
wire n_17542;
wire n_7660;
wire n_6915;
wire n_18235;
wire n_12529;
wire n_15708;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_17072;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_17889;
wire n_8979;
wire n_6522;
wire n_14053;
wire n_5906;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_16564;
wire n_17189;
wire n_14581;
wire n_5660;
wire n_7890;
wire n_12785;
wire n_17073;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_15312;
wire n_6675;
wire n_6270;
wire n_14155;
wire n_18111;
wire n_12461;
wire n_6808;
wire n_13603;
wire n_16091;
wire n_16395;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_7006;
wire n_6931;
wire n_5783;
wire n_6207;
wire n_5821;
wire n_15818;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_6079;
wire n_17231;
wire n_16481;
wire n_7948;
wire n_17809;
wire n_9082;
wire n_10925;
wire n_17900;
wire n_9879;
wire n_11158;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_15878;
wire n_16430;
wire n_17238;
wire n_11669;
wire n_16252;
wire n_14390;
wire n_8264;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_16160;
wire n_16715;
wire n_12078;
wire n_16565;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_10618;
wire n_8135;
wire n_18591;
wire n_15647;
wire n_9594;
wire n_7837;
wire n_16945;
wire n_9832;
wire n_16620;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_18187;
wire n_18462;
wire n_18260;
wire n_6427;
wire n_6580;
wire n_9898;
wire n_11739;
wire n_5500;
wire n_10497;
wire n_6412;
wire n_14561;
wire n_9445;
wire n_18410;
wire n_14978;
wire n_18405;
wire n_7627;
wire n_13301;
wire n_9803;
wire n_13293;
wire n_16698;
wire n_17041;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_6346;
wire n_14381;
wire n_15709;
wire n_5215;
wire n_7860;
wire n_18353;
wire n_15729;
wire n_8408;
wire n_12639;
wire n_17519;
wire n_18590;
wire n_14212;
wire n_5386;
wire n_10661;
wire n_7335;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_7811;
wire n_13158;
wire n_14737;
wire n_11676;
wire n_11044;
wire n_14649;
wire n_11771;
wire n_15967;
wire n_16870;
wire n_12266;
wire n_15940;
wire n_16949;
wire n_12175;
wire n_15530;
wire n_13536;
wire n_10512;
wire n_13833;
wire n_14714;
wire n_11384;
wire n_16518;
wire n_12287;
wire n_11679;
wire n_8450;
wire n_17665;
wire n_8273;
wire n_17799;
wire n_9867;
wire n_7499;
wire n_6059;
wire n_12353;
wire n_14441;
wire n_14129;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_16962;
wire n_7292;
wire n_12398;
wire n_17089;
wire n_10967;
wire n_13485;
wire n_9087;
wire n_7870;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_17832;
wire n_12991;
wire n_16264;
wire n_18377;
wire n_11134;
wire n_7397;
wire n_10789;
wire n_15333;
wire n_12705;
wire n_13735;
wire n_17020;
wire n_17316;
wire n_7977;
wire n_8886;
wire n_6117;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_5618;
wire n_8312;
wire n_6861;
wire n_6781;
wire n_11828;
wire n_14470;
wire n_12326;
wire n_15497;
wire n_14264;
wire n_7847;
wire n_8506;
wire n_14115;
wire n_16735;
wire n_15952;
wire n_16635;
wire n_6494;
wire n_13830;
wire n_13178;
wire n_18585;
wire n_6133;
wire n_16365;
wire n_11548;
wire n_13041;
wire n_17037;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_14184;
wire n_7822;
wire n_6453;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_5247;
wire n_6127;
wire n_14183;
wire n_10762;
wire n_11452;
wire n_11342;
wire n_11362;
wire n_17751;
wire n_15734;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_14200;
wire n_6006;
wire n_10797;
wire n_7289;
wire n_11266;
wire n_17656;
wire n_14110;
wire n_16558;
wire n_12309;
wire n_7926;
wire n_14806;
wire n_6598;
wire n_7399;
wire n_5338;
wire n_12479;
wire n_7354;
wire n_15568;
wire n_8352;
wire n_12502;
wire n_18312;
wire n_13824;
wire n_10360;
wire n_7960;
wire n_15620;
wire n_9450;
wire n_18053;
wire n_5689;
wire n_13953;
wire n_7482;
wire n_12912;
wire n_14847;
wire n_10312;
wire n_12211;
wire n_16777;
wire n_16859;
wire n_6115;
wire n_13377;
wire n_16703;
wire n_12454;
wire n_18308;
wire n_8143;
wire n_10480;
wire n_9223;
wire n_13191;
wire n_16493;
wire n_6048;
wire n_6416;
wire n_10131;
wire n_12537;
wire n_6838;
wire n_15464;
wire n_17741;
wire n_17183;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_17582;
wire n_11988;
wire n_17465;
wire n_12600;
wire n_12921;
wire n_14536;
wire n_13226;
wire n_6139;
wire n_5931;
wire n_15930;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_17943;
wire n_13686;
wire n_6256;
wire n_7965;
wire n_13645;
wire n_15645;
wire n_16433;
wire n_6613;
wire n_12919;
wire n_11438;
wire n_11244;
wire n_18577;
wire n_14432;
wire n_15965;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_16753;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_18473;
wire n_6361;
wire n_9880;
wire n_13253;
wire n_17485;
wire n_14321;
wire n_8183;
wire n_14981;
wire n_11348;
wire n_16098;
wire n_11245;
wire n_9685;
wire n_7474;
wire n_6085;
wire n_11169;
wire n_11685;
wire n_5731;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_8650;
wire n_12422;
wire n_17614;
wire n_6678;
wire n_11546;
wire n_15259;
wire n_16946;
wire n_17843;
wire n_14654;
wire n_15460;
wire n_8662;
wire n_10503;
wire n_14422;
wire n_15058;
wire n_9694;
wire n_7158;
wire n_14664;
wire n_16539;
wire n_16636;
wire n_13215;
wire n_13400;
wire n_14971;
wire n_9905;
wire n_16834;
wire n_10465;
wire n_9948;
wire n_14630;
wire n_16073;
wire n_12429;
wire n_10590;
wire n_17048;
wire n_13782;
wire n_14734;
wire n_15476;
wire n_14494;
wire n_8526;
wire n_13331;
wire n_14956;
wire n_7325;
wire n_13751;
wire n_10887;
wire n_14866;
wire n_9456;
wire n_16876;
wire n_7044;
wire n_17150;
wire n_14019;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_18593;
wire n_9923;
wire n_5883;
wire n_13743;
wire n_17769;
wire n_7166;
wire n_13812;
wire n_14970;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_13378;
wire n_6560;
wire n_14055;
wire n_11319;
wire n_7028;
wire n_7838;
wire n_9890;
wire n_11492;
wire n_5629;
wire n_12136;
wire n_16981;
wire n_16969;
wire n_7873;
wire n_6535;
wire n_16418;
wire n_12731;
wire n_17046;
wire n_16138;
wire n_12399;
wire n_16644;
wire n_17795;
wire n_7518;
wire n_12342;
wire n_12640;
wire n_7414;
wire n_9817;
wire n_9744;
wire n_6147;
wire n_10063;
wire n_9199;
wire n_13092;
wire n_14292;
wire n_9548;
wire n_8973;
wire n_11160;
wire n_6448;
wire n_13544;
wire n_7791;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_12533;
wire n_18172;
wire n_9862;
wire n_5934;
wire n_7431;
wire n_5434;
wire n_12616;
wire n_11385;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_18333;
wire n_12535;
wire n_12178;
wire n_14375;
wire n_17214;
wire n_12653;
wire n_6643;
wire n_12327;
wire n_17982;
wire n_7146;
wire n_9471;
wire n_16580;
wire n_18081;
wire n_11346;
wire n_18498;
wire n_17012;
wire n_10091;
wire n_11638;
wire n_17210;
wire n_6157;
wire n_14896;
wire n_9363;
wire n_12047;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_17181;
wire n_17440;
wire n_18206;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_14810;
wire n_9069;
wire n_13110;
wire n_15719;
wire n_14879;
wire n_16628;
wire n_16143;
wire n_18387;
wire n_17371;
wire n_5852;
wire n_14030;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_17274;
wire n_15164;
wire n_18344;
wire n_8249;
wire n_16660;
wire n_7052;
wire n_11343;
wire n_16755;
wire n_12348;
wire n_16929;
wire n_16099;
wire n_10496;
wire n_12257;
wire n_15590;
wire n_15770;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_14149;
wire n_13394;
wire n_16853;
wire n_10843;
wire n_13391;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_13384;
wire n_14680;
wire n_16869;
wire n_8234;
wire n_16048;
wire n_18225;
wire n_5321;
wire n_16835;
wire n_9960;
wire n_10997;
wire n_16262;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_18438;
wire n_17127;
wire n_10998;
wire n_15422;
wire n_9003;
wire n_9280;
wire n_16863;
wire n_18285;
wire n_6073;
wire n_7502;
wire n_12418;
wire n_14216;
wire n_6331;
wire n_5290;
wire n_16380;
wire n_14837;
wire n_13498;
wire n_7312;
wire n_13263;
wire n_7919;
wire n_14877;
wire n_15203;
wire n_11269;
wire n_10800;
wire n_17962;
wire n_7085;
wire n_11491;
wire n_16849;
wire n_12065;
wire n_13950;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_18289;
wire n_11408;
wire n_14048;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_14103;
wire n_16112;
wire n_5210;
wire n_13183;
wire n_6689;
wire n_13732;
wire n_14968;
wire n_16422;
wire n_10993;
wire n_15891;
wire n_7632;
wire n_12519;
wire n_14985;
wire n_9172;
wire n_12769;
wire n_15542;
wire n_15910;
wire n_14653;
wire n_17184;
wire n_6405;
wire n_7580;
wire n_17275;
wire n_14077;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_17573;
wire n_11311;
wire n_17734;
wire n_10112;
wire n_14443;
wire n_10765;
wire n_16136;
wire n_6698;
wire n_15263;
wire n_11792;
wire n_14285;
wire n_18553;
wire n_17345;
wire n_7304;
wire n_17770;
wire n_9734;
wire n_7288;
wire n_8558;
wire n_13242;
wire n_10489;
wire n_7707;
wire n_16325;
wire n_7223;
wire n_12421;
wire n_13282;
wire n_14436;
wire n_16842;
wire n_7833;
wire n_12113;
wire n_14868;
wire n_17355;
wire n_14599;
wire n_5512;
wire n_7274;
wire n_16087;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_14351;
wire n_6206;
wire n_9068;
wire n_13352;
wire n_8136;
wire n_9808;
wire n_17648;
wire n_18534;
wire n_6610;
wire n_17853;
wire n_18116;
wire n_7445;
wire n_14812;
wire n_10612;
wire n_11086;
wire n_7466;
wire n_6529;
wire n_10260;
wire n_11293;
wire n_14728;
wire n_17871;
wire n_6363;
wire n_6750;
wire n_12285;
wire n_13310;
wire n_11710;
wire n_8619;
wire n_11568;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_18217;
wire n_9150;
wire n_10134;
wire n_14508;
wire n_15122;
wire n_11603;
wire n_13798;
wire n_7277;
wire n_16894;
wire n_6455;
wire n_15277;
wire n_18435;
wire n_15092;
wire n_13804;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_14778;
wire n_17294;
wire n_15714;
wire n_17270;
wire n_16932;
wire n_18535;
wire n_15842;
wire n_13099;
wire n_12015;
wire n_8146;
wire n_13690;
wire n_14822;
wire n_18457;
wire n_8813;
wire n_18516;
wire n_5607;
wire n_11562;
wire n_7695;
wire n_10194;
wire n_14566;
wire n_17085;
wire n_7179;
wire n_10356;
wire n_17461;
wire n_7122;
wire n_18216;
wire n_10173;
wire n_12157;
wire n_7165;
wire n_7869;
wire n_5999;
wire n_13386;
wire n_13846;
wire n_8910;
wire n_12311;
wire n_6203;
wire n_6408;
wire n_14374;
wire n_15806;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_13064;
wire n_14815;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_16246;
wire n_13619;
wire n_16437;
wire n_8470;
wire n_9587;
wire n_18508;
wire n_12031;
wire n_5341;
wire n_16480;
wire n_8643;
wire n_17351;
wire n_15660;
wire n_9278;
wire n_10671;
wire n_15357;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_11718;
wire n_8565;
wire n_10821;
wire n_13648;
wire n_17657;
wire n_14831;
wire n_14996;
wire n_11170;
wire n_17683;
wire n_11758;
wire n_12126;
wire n_14383;
wire n_8550;
wire n_14543;
wire n_16695;
wire n_9396;
wire n_6892;
wire n_11094;
wire n_14450;
wire n_14747;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_15722;
wire n_14683;
wire n_10599;
wire n_9667;
wire n_14192;
wire n_17052;
wire n_14181;
wire n_6401;
wire n_7322;
wire n_17378;
wire n_15278;
wire n_9053;
wire n_11658;
wire n_15504;
wire n_11893;
wire n_18054;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_9739;
wire n_10573;
wire n_13492;
wire n_14358;
wire n_9480;
wire n_14001;
wire n_14213;
wire n_17320;
wire n_17885;
wire n_5562;
wire n_15397;
wire n_7051;
wire n_10850;
wire n_15840;
wire n_9185;
wire n_8477;
wire n_17886;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_12195;
wire n_13376;
wire n_14842;
wire n_13115;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_13864;
wire n_16855;
wire n_5911;
wire n_11601;
wire n_13289;
wire n_15279;
wire n_11971;
wire n_13182;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_16265;
wire n_16937;
wire n_5622;
wire n_9919;
wire n_12135;
wire n_16466;
wire n_6574;
wire n_11116;
wire n_13324;
wire n_12604;
wire n_6571;
wire n_13305;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_17484;
wire n_8876;
wire n_15215;
wire n_17092;
wire n_17748;
wire n_9151;
wire n_8829;
wire n_16379;
wire n_16728;
wire n_9359;
wire n_7824;
wire n_17202;
wire n_13381;
wire n_18080;
wire n_13236;
wire n_14189;
wire n_14299;
wire n_7094;
wire n_15761;
wire n_7097;
wire n_16320;
wire n_5413;
wire n_8140;
wire n_8971;
wire n_15111;
wire n_18076;
wire n_8060;
wire n_16667;
wire n_16897;
wire n_10558;
wire n_7036;
wire n_18563;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_17603;
wire n_15273;
wire n_6392;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_17470;
wire n_13777;
wire n_15301;
wire n_9049;
wire n_7351;
wire n_13718;
wire n_17621;
wire n_9352;
wire n_14775;
wire n_7608;
wire n_5779;
wire n_17053;
wire n_6260;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_13202;
wire n_7909;
wire n_15350;
wire n_7413;
wire n_13638;
wire n_16803;
wire n_6303;
wire n_16756;
wire n_17229;
wire n_8935;
wire n_14392;
wire n_17948;
wire n_11340;
wire n_15759;
wire n_10734;
wire n_6286;
wire n_16441;
wire n_16965;
wire n_7675;
wire n_8267;
wire n_15383;
wire n_11903;
wire n_7027;
wire n_7992;
wire n_13279;
wire n_13644;
wire n_6912;
wire n_11560;
wire n_10330;
wire n_10395;
wire n_7175;
wire n_8276;
wire n_13291;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_14966;
wire n_11465;
wire n_7524;
wire n_15255;
wire n_8027;
wire n_15897;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_17808;
wire n_11265;
wire n_16729;
wire n_9370;
wire n_11125;
wire n_9670;
wire n_13136;
wire n_13513;
wire n_17244;
wire n_12916;
wire n_18406;
wire n_18044;
wire n_9334;
wire n_7783;
wire n_13220;
wire n_15131;
wire n_6692;
wire n_10276;
wire n_14322;
wire n_12331;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_12531;
wire n_8245;
wire n_15072;
wire n_6036;
wire n_8471;
wire n_12521;
wire n_11302;
wire n_12910;
wire n_13349;
wire n_9956;
wire n_18215;
wire n_9800;
wire n_17007;
wire n_8454;
wire n_6552;
wire n_17096;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_15509;
wire n_10098;
wire n_11745;
wire n_17005;
wire n_8891;
wire n_15240;
wire n_11690;
wire n_16194;
wire n_9487;
wire n_11707;
wire n_5591;
wire n_11373;
wire n_7697;
wire n_16791;
wire n_14608;
wire n_6403;
wire n_15564;
wire n_7306;
wire n_13835;
wire n_16153;
wire n_16260;
wire n_7947;
wire n_10118;
wire n_16826;
wire n_17002;
wire n_14350;
wire n_7470;
wire n_7547;
wire n_7733;
wire n_6013;
wire n_13815;
wire n_13800;
wire n_7693;
wire n_17405;
wire n_9557;
wire n_15957;
wire n_6491;
wire n_16319;
wire n_16321;
wire n_17259;
wire n_14039;
wire n_14072;
wire n_15662;
wire n_17120;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_18578;
wire n_13039;
wire n_13773;
wire n_13130;
wire n_14109;
wire n_8582;
wire n_10441;
wire n_17237;
wire n_6982;
wire n_5518;
wire n_10002;
wire n_6293;
wire n_9124;
wire n_6661;
wire n_15671;
wire n_5847;
wire n_13719;
wire n_7345;
wire n_6049;
wire n_9762;
wire n_8847;
wire n_11242;
wire n_8957;
wire n_14136;
wire n_17526;
wire n_17974;
wire n_7385;
wire n_10923;
wire n_14548;
wire n_15793;
wire n_15923;
wire n_6558;
wire n_14176;
wire n_11149;
wire n_10841;
wire n_16076;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_13694;
wire n_18209;
wire n_12313;
wire n_8488;
wire n_9271;
wire n_18071;
wire n_17747;
wire n_17494;
wire n_9543;
wire n_13688;
wire n_14661;
wire n_11396;
wire n_8356;
wire n_6136;
wire n_9660;
wire n_15196;
wire n_16176;
wire n_16384;
wire n_16416;
wire n_11443;
wire n_9483;
wire n_15765;
wire n_6855;
wire n_15305;
wire n_15588;
wire n_14754;
wire n_10665;
wire n_18176;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_15020;
wire n_16233;
wire n_13467;
wire n_5357;
wire n_6091;
wire n_13093;
wire n_17344;
wire n_13062;
wire n_9328;
wire n_14252;
wire n_7857;
wire n_7481;
wire n_16511;
wire n_18374;
wire n_14130;
wire n_15830;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_14930;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_16596;
wire n_6312;
wire n_8747;
wire n_11532;
wire n_9539;
wire n_6668;
wire n_9415;
wire n_15274;
wire n_18548;
wire n_15548;
wire n_14343;
wire n_16410;
wire n_9385;
wire n_9147;
wire n_11209;
wire n_16714;
wire n_7653;
wire n_13462;
wire n_5381;
wire n_8354;
wire n_15918;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_14276;
wire n_6959;
wire n_5918;
wire n_16212;
wire n_8353;
wire n_13752;
wire n_8922;
wire n_6388;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_13185;
wire n_9027;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_18450;
wire n_13596;
wire n_6995;
wire n_10902;
wire n_12889;
wire n_13855;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_18092;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_18148;
wire n_16313;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_11304;
wire n_17957;
wire n_9642;
wire n_17058;
wire n_18309;
wire n_16363;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_15232;
wire n_7475;
wire n_10485;
wire n_14231;
wire n_18448;
wire n_12105;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_13219;
wire n_14329;
wire n_5673;
wire n_5443;
wire n_17449;
wire n_6351;
wire n_16895;
wire n_9079;
wire n_15544;
wire n_15721;
wire n_9382;
wire n_16392;
wire n_10282;
wire n_7668;
wire n_6212;
wire n_16145;
wire n_17602;
wire n_9775;
wire n_10444;
wire n_17512;
wire n_11377;
wire n_8653;
wire n_8018;
wire n_13295;
wire n_15142;
wire n_8920;
wire n_16906;
wire n_18194;
wire n_18557;
wire n_17693;
wire n_10913;
wire n_7937;
wire n_18409;
wire n_17521;
wire n_9176;
wire n_6829;
wire n_17838;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_15991;
wire n_5823;
wire n_17981;
wire n_7305;
wire n_13388;
wire n_13160;
wire n_13731;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_15249;
wire n_6682;
wire n_17337;
wire n_17477;
wire n_6334;
wire n_6823;
wire n_14550;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_14503;
wire n_16780;
wire n_12248;
wire n_13818;
wire n_15024;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_15346;
wire n_13477;
wire n_17754;
wire n_8884;
wire n_8803;
wire n_14886;
wire n_18200;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_10978;
wire n_5537;
wire n_8222;
wire n_13808;
wire n_14644;
wire n_6822;
wire n_11715;
wire n_18478;
wire n_8553;
wire n_7071;
wire n_9706;
wire n_15174;
wire n_15454;
wire n_10642;
wire n_15213;
wire n_17068;
wire n_17904;
wire n_18428;
wire n_12181;
wire n_10187;
wire n_10387;
wire n_11014;
wire n_13764;
wire n_14560;
wire n_17508;
wire n_15033;
wire n_17257;
wire n_8751;
wire n_17789;
wire n_11864;
wire n_14829;
wire n_11007;
wire n_11224;
wire n_15473;
wire n_11006;
wire n_15584;
wire n_9564;
wire n_15018;
wire n_7391;
wire n_8790;
wire n_15569;
wire n_9230;
wire n_6617;
wire n_10219;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_15193;
wire n_14067;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_18386;
wire n_16515;
wire n_14108;
wire n_6389;
wire n_6137;
wire n_15903;
wire n_14833;
wire n_17914;
wire n_10364;
wire n_15439;
wire n_10479;
wire n_11422;
wire n_16049;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_13660;
wire n_8398;
wire n_14480;
wire n_13970;
wire n_8178;
wire n_6801;
wire n_15247;
wire n_16656;
wire n_12489;
wire n_8491;
wire n_14000;
wire n_14372;
wire n_18099;
wire n_5630;
wire n_10065;
wire n_17911;
wire n_12046;
wire n_10212;
wire n_16610;
wire n_9283;
wire n_8700;
wire n_12030;
wire n_12738;
wire n_13408;
wire n_15062;
wire n_17585;
wire n_18566;
wire n_15248;
wire n_13727;
wire n_17500;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_10268;
wire n_15236;
wire n_14801;
wire n_14098;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_12601;
wire n_14482;
wire n_15399;
wire n_16178;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_13641;
wire n_17174;
wire n_17549;
wire n_14223;
wire n_15962;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_17473;
wire n_14947;
wire n_17746;
wire n_17304;
wire n_5505;
wire n_5868;
wire n_18393;
wire n_10305;
wire n_8560;
wire n_14983;
wire n_17332;
wire n_14748;
wire n_10559;
wire n_13173;
wire n_8439;
wire n_16862;
wire n_18434;
wire n_9641;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_15355;
wire n_15669;
wire n_18466;
wire n_18522;
wire n_12059;
wire n_12488;
wire n_15945;
wire n_18018;
wire n_18541;
wire n_7321;
wire n_18257;
wire n_14848;
wire n_5289;
wire n_8200;
wire n_15845;
wire n_16055;
wire n_11110;
wire n_7154;
wire n_6129;
wire n_16232;
wire n_17338;
wire n_6518;
wire n_18179;
wire n_18564;
wire n_16211;
wire n_15001;
wire n_8304;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_18072;
wire n_5401;
wire n_18048;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_14544;
wire n_13328;
wire n_7537;
wire n_10516;
wire n_8675;
wire n_10892;
wire n_6254;
wire n_5989;
wire n_15924;
wire n_18556;
wire n_10493;
wire n_17906;
wire n_13542;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_5769;
wire n_10405;
wire n_15037;
wire n_15130;
wire n_16122;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_17386;
wire n_14604;
wire n_14735;
wire n_7964;
wire n_17091;
wire n_9016;
wire n_14426;
wire n_13101;
wire n_11887;
wire n_15456;
wire n_14349;
wire n_6278;
wire n_17442;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_17852;
wire n_11545;
wire n_9729;
wire n_12691;
wire n_8846;
wire n_8315;
wire n_16446;
wire n_12471;
wire n_11033;
wire n_15885;
wire n_17528;
wire n_12451;
wire n_11040;
wire n_12665;
wire n_16367;
wire n_16526;
wire n_17243;
wire n_16397;
wire n_11754;
wire n_11850;
wire n_14916;
wire n_15740;
wire n_18203;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_14356;
wire n_17467;
wire n_5581;
wire n_13748;
wire n_9029;
wire n_9411;
wire n_11672;
wire n_16926;
wire n_6837;
wire n_10353;
wire n_16006;
wire n_17418;
wire n_10847;
wire n_12651;
wire n_10451;
wire n_11043;
wire n_15801;
wire n_17778;
wire n_5303;
wire n_16476;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_16373;
wire n_9414;
wire n_18539;
wire n_16719;
wire n_7023;
wire n_12003;
wire n_9615;
wire n_14205;
wire n_14564;
wire n_7496;
wire n_11277;
wire n_12165;
wire n_18532;
wire n_18416;
wire n_10866;
wire n_17606;
wire n_14190;
wire n_7410;
wire n_18127;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_14600;
wire n_8777;
wire n_17223;
wire n_11061;
wire n_11763;
wire n_16495;
wire n_15546;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_8535;
wire n_10653;
wire n_11587;
wire n_6373;
wire n_5375;
wire n_11534;
wire n_12280;
wire n_9221;
wire n_12492;
wire n_13581;
wire n_13461;
wire n_14344;
wire n_15742;
wire n_16686;
wire n_12972;
wire n_16282;
wire n_16347;
wire n_5370;
wire n_17011;
wire n_13789;
wire n_5601;
wire n_9811;
wire n_5784;
wire n_7899;
wire n_8631;
wire n_13188;
wire n_14511;
wire n_7906;
wire n_16385;
wire n_13286;
wire n_17639;
wire n_5248;
wire n_9951;
wire n_7131;
wire n_14723;
wire n_6411;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_8909;
wire n_14488;
wire n_11032;
wire n_13582;
wire n_10507;
wire n_16356;
wire n_17950;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_18162;
wire n_11843;
wire n_17437;
wire n_10045;
wire n_11174;
wire n_14614;
wire n_13531;
wire n_18574;
wire n_7797;
wire n_11335;
wire n_11629;
wire n_15147;
wire n_6381;
wire n_7030;
wire n_18606;
wire n_6656;
wire n_9730;
wire n_13880;
wire n_18544;
wire n_7687;
wire n_9554;
wire n_10294;
wire n_13988;
wire n_18246;
wire n_10106;
wire n_18251;
wire n_5635;
wire n_17865;
wire n_7582;
wire n_17180;
wire n_15272;
wire n_9934;
wire n_10541;
wire n_17169;
wire n_13609;
wire n_14587;
wire n_6546;
wire n_5528;
wire n_9234;
wire n_10674;
wire n_8959;
wire n_16886;
wire n_6534;
wire n_17326;
wire n_10614;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_13679;
wire n_10417;
wire n_15927;
wire n_16011;
wire n_16877;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_18169;
wire n_5778;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_17370;
wire n_18185;
wire n_8087;
wire n_15834;
wire n_13276;
wire n_9910;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_14458;
wire n_8938;
wire n_5665;
wire n_16790;
wire n_16058;
wire n_11801;
wire n_17255;
wire n_17540;
wire n_13217;
wire n_16519;
wire n_12073;
wire n_13655;
wire n_16994;
wire n_6898;
wire n_6596;
wire n_5363;
wire n_17810;
wire n_10743;
wire n_13424;
wire n_16332;
wire n_14658;
wire n_15066;
wire n_14830;
wire n_14397;
wire n_17971;
wire n_10853;
wire n_7867;
wire n_9651;
wire n_13565;
wire n_14281;
wire n_13755;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_6135;
wire n_13802;
wire n_14594;
wire n_15474;
wire n_17303;
wire n_18213;
wire n_18559;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_15316;
wire n_10270;
wire n_6814;
wire n_10557;
wire n_11115;
wire n_8669;
wire n_12978;
wire n_13784;
wire n_8001;
wire n_7525;
wire n_13468;
wire n_7257;
wire n_12363;
wire n_18201;
wire n_9372;
wire n_7553;
wire n_17417;
wire n_7529;
wire n_15668;
wire n_6791;
wire n_15137;
wire n_14233;
wire n_8496;
wire n_11915;
wire n_13704;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_11788;
wire n_12544;
wire n_13036;
wire n_14146;
wire n_7650;
wire n_12476;
wire n_13199;
wire n_17297;
wire n_8568;
wire n_6903;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_18423;
wire n_12023;
wire n_17655;
wire n_8637;
wire n_6168;
wire n_16225;
wire n_6881;
wire n_16677;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_17260;
wire n_13413;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_13002;
wire n_15153;
wire n_17324;
wire n_12632;
wire n_12620;
wire n_7520;
wire n_9831;
wire n_13203;
wire n_13868;
wire n_6309;
wire n_7903;
wire n_18245;
wire n_9697;
wire n_18596;
wire n_11303;
wire n_11877;
wire n_6733;
wire n_14462;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_13285;
wire n_5430;
wire n_5942;
wire n_8610;
wire n_7894;
wire n_7137;
wire n_9902;
wire n_18414;
wire n_14933;
wire n_8362;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_17367;
wire n_8256;
wire n_15521;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_18415;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_12598;
wire n_9039;
wire n_13374;
wire n_11854;
wire n_16458;
wire n_12416;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_8704;
wire n_8265;
wire n_7639;
wire n_16520;
wire n_5762;
wire n_17589;
wire n_6132;
wire n_5211;
wire n_5336;
wire n_11609;
wire n_18287;
wire n_5447;
wire n_16464;
wire n_17493;
wire n_17389;
wire n_7743;
wire n_13230;
wire n_9294;
wire n_12811;
wire n_12494;
wire n_12186;
wire n_11747;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_13032;
wire n_13826;
wire n_7054;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_10021;
wire n_5327;
wire n_13684;
wire n_14199;
wire n_16673;
wire n_17858;
wire n_9146;
wire n_9125;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_14027;
wire n_15108;
wire n_15753;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_17941;
wire n_8941;
wire n_16316;
wire n_17093;
wire n_5747;
wire n_17685;
wire n_16898;
wire n_18331;
wire n_9073;
wire n_10075;
wire n_16357;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_18325;
wire n_17762;
wire n_6171;
wire n_13750;
wire n_17291;
wire n_8775;
wire n_14104;
wire n_12272;
wire n_17895;
wire n_9302;
wire n_5519;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_14684;
wire n_11895;
wire n_13458;
wire n_6269;
wire n_7092;
wire n_5753;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_15713;
wire n_9171;
wire n_10886;
wire n_14857;
wire n_5233;
wire n_18124;
wire n_8279;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_12191;
wire n_17432;
wire n_9580;
wire n_8019;
wire n_14572;
wire n_13963;
wire n_9972;
wire n_13091;
wire n_13003;
wire n_6083;
wire n_17707;
wire n_12909;
wire n_6434;
wire n_6387;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_9465;
wire n_16417;
wire n_17880;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_13811;
wire n_14316;
wire n_17242;
wire n_7726;
wire n_8807;
wire n_18120;
wire n_5436;
wire n_17026;
wire n_13839;
wire n_5231;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_14011;
wire n_13954;
wire n_10436;
wire n_18300;
wire n_8464;
wire n_15701;
wire n_6547;
wire n_8799;
wire n_12794;
wire n_5193;
wire n_6423;
wire n_15496;
wire n_9442;
wire n_6342;
wire n_18571;
wire n_6641;
wire n_17744;
wire n_15260;
wire n_6984;
wire n_18394;
wire n_15612;
wire n_17392;
wire n_5789;
wire n_15104;
wire n_10763;
wire n_7441;
wire n_9957;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_16374;
wire n_7106;
wire n_18173;
wire n_7213;
wire n_17251;
wire n_12112;
wire n_13060;
wire n_14689;
wire n_16187;
wire n_10245;
wire n_17586;
wire n_5961;
wire n_10905;
wire n_14132;
wire n_11235;
wire n_9449;
wire n_14817;
wire n_5866;
wire n_9050;
wire n_6507;
wire n_9313;
wire n_6399;
wire n_6687;
wire n_5822;
wire n_9173;
wire n_17381;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_15055;
wire n_5726;
wire n_11015;
wire n_9563;
wire n_14087;
wire n_9160;
wire n_17077;
wire n_5364;
wire n_9974;
wire n_17702;
wire n_12129;
wire n_14753;
wire n_11166;
wire n_15980;
wire n_7031;
wire n_9285;
wire n_13658;
wire n_18093;
wire n_5533;
wire n_16595;
wire n_7763;
wire n_9631;
wire n_14671;
wire n_8033;
wire n_15172;
wire n_14751;
wire n_6194;
wire n_14438;
wire n_16454;
wire n_17977;
wire n_8393;
wire n_16253;
wire n_7133;
wire n_16561;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_10784;
wire n_12202;
wire n_18441;
wire n_14674;
wire n_13836;
wire n_8463;
wire n_18313;
wire n_8153;
wire n_12815;
wire n_15913;
wire n_6524;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_18554;
wire n_9945;
wire n_18077;
wire n_8661;
wire n_16089;
wire n_12431;
wire n_7424;
wire n_7523;
wire n_17694;
wire n_8654;
wire n_16314;
wire n_11855;
wire n_14229;
wire n_15060;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_15115;
wire n_16671;
wire n_15520;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_17628;
wire n_11156;
wire n_8531;
wire n_14188;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_13799;
wire n_5718;
wire n_16084;
wire n_6459;
wire n_6505;
wire n_16139;
wire n_12333;
wire n_12636;
wire n_8379;
wire n_8609;
wire n_13854;
wire n_17666;
wire n_18250;
wire n_17219;
wire n_11227;
wire n_7626;
wire n_13576;
wire n_15380;
wire n_13100;
wire n_7310;
wire n_16154;
wire n_12334;
wire n_17451;
wire n_6686;
wire n_15956;
wire n_18397;
wire n_9209;
wire n_7311;
wire n_6001;
wire n_18234;
wire n_7669;
wire n_11218;
wire n_12119;
wire n_12618;
wire n_11787;
wire n_5958;
wire n_8793;
wire n_16059;
wire n_12355;
wire n_8103;
wire n_15052;
wire n_9767;
wire n_10195;
wire n_9838;
wire n_13722;
wire n_9300;
wire n_16093;
wire n_11500;
wire n_12943;
wire n_17266;
wire n_17598;
wire n_15129;
wire n_17146;
wire n_7327;
wire n_14306;
wire n_16209;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_8367;
wire n_11891;
wire n_16276;
wire n_17956;
wire n_7367;
wire n_14752;
wire n_18427;
wire n_5792;
wire n_11021;
wire n_12401;
wire n_16439;
wire n_8543;
wire n_16502;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_14897;
wire n_15447;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_6905;
wire n_16688;
wire n_18600;
wire n_10243;
wire n_9700;
wire n_10564;
wire n_17520;
wire n_17633;
wire n_18114;
wire n_8682;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_17815;
wire n_7655;
wire n_5554;
wire n_7244;
wire n_15925;
wire n_10745;
wire n_7368;
wire n_18255;
wire n_17958;
wire n_10596;
wire n_18276;
wire n_5553;
wire n_8011;
wire n_7633;
wire n_13937;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_10263;
wire n_5790;
wire n_11509;
wire n_8640;
wire n_14359;
wire n_8063;
wire n_15141;
wire n_11960;
wire n_12599;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_12411;
wire n_16933;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_12465;
wire n_7427;
wire n_10605;
wire n_13532;
wire n_11029;
wire n_14013;
wire n_14419;
wire n_13250;
wire n_13118;
wire n_5404;
wire n_9933;
wire n_17390;
wire n_11449;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_9892;
wire n_15251;
wire n_8570;
wire n_6163;
wire n_16727;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_5549;
wire n_9408;
wire n_6785;
wire n_6553;
wire n_15854;
wire n_10163;
wire n_10454;
wire n_17409;
wire n_17630;
wire n_15401;
wire n_13339;
wire n_5444;
wire n_12568;
wire n_16163;
wire n_13478;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_18256;
wire n_12970;
wire n_8916;
wire n_8902;
wire n_14295;
wire n_7557;
wire n_10087;
wire n_17518;
wire n_16544;
wire n_8843;
wire n_10146;
wire n_9891;
wire n_7128;
wire n_9946;
wire n_12959;
wire n_17529;
wire n_15810;
wire n_14367;
wire n_9885;
wire n_6849;
wire n_7594;
wire n_12330;
wire n_13915;
wire n_8129;
wire n_8162;
wire n_14890;
wire n_14819;
wire n_15057;
wire n_15871;
wire n_13906;
wire n_7457;
wire n_18263;
wire n_10643;
wire n_16974;
wire n_16300;
wire n_8744;
wire n_18288;
wire n_10504;
wire n_5824;
wire n_7788;
wire n_10872;
wire n_5488;
wire n_13783;
wire n_6760;
wire n_10701;
wire n_14265;
wire n_13987;
wire n_13664;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_13566;
wire n_15626;
wire n_12591;
wire n_12466;
wire n_18060;
wire n_15775;
wire n_9509;
wire n_8286;
wire n_17346;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_5329;
wire n_9015;
wire n_9925;
wire n_9757;
wire n_5637;
wire n_16066;
wire n_10874;
wire n_6825;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_11831;
wire n_13726;
wire n_9628;
wire n_14399;
wire n_7767;
wire n_14412;
wire n_16213;
wire n_16408;
wire n_8294;
wire n_17587;
wire n_9419;
wire n_12243;
wire n_12279;
wire n_16402;
wire n_6611;
wire n_8562;
wire n_13705;
wire n_18279;
wire n_12614;
wire n_17986;
wire n_11378;
wire n_10250;
wire n_14631;
wire n_5728;
wire n_17771;
wire n_5471;
wire n_10032;
wire n_11433;
wire n_10592;
wire n_9277;
wire n_9257;
wire n_17773;
wire n_14063;
wire n_18130;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_13425;
wire n_17070;
wire n_16657;
wire n_17105;
wire n_8170;
wire n_9159;
wire n_5843;
wire n_11558;
wire n_17978;
wire n_17233;
wire n_18515;
wire n_7744;
wire n_7021;
wire n_10595;
wire n_13591;
wire n_7748;
wire n_8537;
wire n_10126;
wire n_6827;
wire n_14421;
wire n_17584;
wire n_18296;
wire n_12041;
wire n_15890;
wire n_11713;
wire n_13653;
wire n_11073;
wire n_15586;
wire n_16972;
wire n_16734;
wire n_5484;
wire n_6355;
wire n_12566;
wire n_17821;
wire n_12931;
wire n_15525;
wire n_17783;
wire n_6227;
wire n_13680;
wire n_7215;
wire n_15157;
wire n_17790;
wire n_7485;
wire n_13074;
wire n_16077;
wire n_9066;
wire n_17566;
wire n_5523;
wire n_14332;
wire n_18379;
wire n_10302;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_14716;
wire n_10645;
wire n_13058;
wire n_15313;
wire n_18342;
wire n_10604;
wire n_11096;
wire n_17398;
wire n_12036;
wire n_12876;
wire n_15286;
wire n_6564;
wire n_11161;
wire n_17650;
wire n_9671;
wire n_8709;
wire n_8782;
wire n_14698;
wire n_12911;
wire n_15715;
wire n_6468;
wire n_12491;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_11216;
wire n_14368;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_18390;
wire n_9857;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_14323;
wire n_12929;
wire n_10882;
wire n_16065;
wire n_18565;
wire n_9338;
wire n_13071;
wire n_6857;
wire n_8144;
wire n_15075;
wire n_12261;
wire n_10435;
wire n_9542;
wire n_12536;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_16333;
wire n_18007;
wire n_6442;
wire n_12106;
wire n_12061;
wire n_18359;
wire n_15116;
wire n_16200;
wire n_14585;
wire n_11085;
wire n_8049;
wire n_16041;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_16541;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_10609;
wire n_11157;
wire n_13739;
wire n_13649;
wire n_14804;
wire n_5594;
wire n_15126;
wire n_12291;
wire n_14510;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_12124;
wire n_11755;
wire n_16497;
wire n_16846;
wire n_9783;
wire n_13806;
wire n_14364;
wire n_9510;
wire n_15472;
wire n_9389;
wire n_18055;
wire n_12074;
wire n_13497;
wire n_9404;
wire n_15406;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_14396;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_13234;
wire n_5292;
wire n_18351;
wire n_9314;
wire n_11918;
wire n_16198;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_14466;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5403;
wire n_14473;
wire n_12887;
wire n_16718;
wire n_5551;
wire n_7652;
wire n_10220;
wire n_10341;
wire n_8701;
wire n_11347;
wire n_16810;
wire n_17635;
wire n_6499;
wire n_10550;
wire n_7830;
wire n_14673;
wire n_15816;
wire n_18158;
wire n_18314;
wire n_12217;
wire n_12365;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_15922;
wire n_8097;
wire n_13738;
wire n_13851;
wire n_9679;
wire n_17341;
wire n_17380;
wire n_14972;
wire n_8084;
wire n_16996;
wire n_9306;
wire n_8645;
wire n_14138;
wire n_13272;
wire n_8712;
wire n_10232;
wire n_14113;
wire n_10461;
wire n_14586;
wire n_8289;
wire n_11178;
wire n_7966;
wire n_8591;
wire n_16411;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_16717;
wire n_16428;
wire n_17652;
wire n_8824;
wire n_11673;
wire n_14938;
wire n_14784;
wire n_11432;
wire n_14641;
wire n_14179;
wire n_17755;
wire n_14031;
wire n_7191;
wire n_16506;
wire n_14979;
wire n_7712;
wire n_10412;
wire n_17543;
wire n_5242;
wire n_15433;
wire n_10326;
wire n_12650;
wire n_15953;
wire n_5219;
wire n_8417;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_10499;
wire n_8340;
wire n_6008;
wire n_12658;
wire n_12487;
wire n_14324;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_5460;
wire n_18425;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_17300;
wire n_13613;
wire n_14740;
wire n_9210;
wire n_12185;
wire n_17763;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_6893;
wire n_5686;
wire n_7406;
wire n_8681;
wire n_5899;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_16044;
wire n_16299;
wire n_17176;
wire n_10617;
wire n_12271;
wire n_12704;
wire n_7807;
wire n_9592;
wire n_18126;
wire n_14198;
wire n_7680;
wire n_9180;
wire n_14846;
wire n_15190;
wire n_10922;
wire n_10544;
wire n_16524;
wire n_17507;
wire n_16909;
wire n_12958;
wire n_13030;
wire n_8172;
wire n_17819;
wire n_9917;
wire n_10718;
wire n_18475;
wire n_12056;
wire n_14539;
wire n_15094;
wire n_8106;
wire n_16880;
wire n_9502;
wire n_13821;
wire n_6447;
wire n_13712;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_9625;
wire n_5937;
wire n_6422;
wire n_13896;
wire n_14761;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_15243;
wire n_16473;
wire n_14420;
wire n_18562;
wire n_11087;
wire n_15041;
wire n_11477;
wire n_17262;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_13299;
wire n_15393;
wire n_13243;
wire n_14314;
wire n_8612;
wire n_13042;
wire n_14144;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_16642;
wire n_15658;
wire n_10095;
wire n_14227;
wire n_13725;
wire n_10309;
wire n_15873;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_8974;
wire n_8268;
wire n_14164;
wire n_9871;
wire n_6160;
wire n_10050;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_17551;
wire n_7066;
wire n_15595;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_18128;
wire n_7789;
wire n_13197;
wire n_10306;
wire n_15081;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_6368;
wire n_10056;
wire n_18408;
wire n_7140;
wire n_16597;
wire n_17627;
wire n_7193;
wire n_6039;
wire n_18180;
wire n_16474;
wire n_11919;
wire n_14860;
wire n_6583;
wire n_10450;
wire n_5721;
wire n_11414;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_16940;
wire n_17419;
wire n_18142;
wire n_12520;
wire n_8515;
wire n_10529;
wire n_17705;
wire n_13632;
wire n_5719;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_17728;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_17134;
wire n_9392;
wire n_13148;
wire n_10429;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_14531;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_17618;
wire n_11538;
wire n_16344;
wire n_10037;
wire n_12808;
wire n_13871;
wire n_18029;
wire n_6707;
wire n_9698;
wire n_13435;
wire n_15408;
wire n_18275;
wire n_12744;
wire n_6064;
wire n_15173;
wire n_11136;
wire n_9903;
wire n_17208;
wire n_13801;
wire n_5793;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_15480;
wire n_10179;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_9499;
wire n_12143;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_13879;
wire n_6647;
wire n_6275;
wire n_14038;
wire n_14771;
wire n_9522;
wire n_5578;
wire n_15617;
wire n_15463;
wire n_18064;
wire n_11215;
wire n_5296;
wire n_11076;
wire n_14339;
wire n_11890;
wire n_9366;
wire n_14253;
wire n_7915;
wire n_7750;
wire n_5893;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_16005;
wire n_9148;
wire n_11806;
wire n_11054;
wire n_15902;
wire n_8406;
wire n_6277;
wire n_15919;
wire n_10754;
wire n_5742;
wire n_11050;
wire n_5207;
wire n_16652;
wire n_12443;
wire n_17714;
wire n_6463;
wire n_5676;
wire n_11683;
wire n_8554;
wire n_10920;
wire n_9275;
wire n_10223;
wire n_8896;
wire n_6051;
wire n_14398;
wire n_11484;
wire n_7206;
wire n_11126;
wire n_7538;
wire n_5674;
wire n_12934;
wire n_18453;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_5282;
wire n_10295;
wire n_9409;
wire n_5464;
wire n_6799;
wire n_17979;
wire n_10336;
wire n_10228;
wire n_17814;
wire n_12555;
wire n_11646;
wire n_7716;
wire n_6487;
wire n_17903;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_8818;
wire n_16648;
wire n_8617;
wire n_16724;
wire n_17953;
wire n_12980;
wire n_13966;
wire n_9881;
wire n_12530;
wire n_8954;
wire n_6807;
wire n_9463;
wire n_12212;
wire n_7251;
wire n_7254;
wire n_10466;
wire n_18178;
wire n_12973;
wire n_7540;
wire n_17313;
wire n_11953;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_13231;
wire n_12624;
wire n_7882;
wire n_16309;
wire n_8552;
wire n_16348;
wire n_16514;
wire n_10425;
wire n_7554;
wire n_8069;
wire n_7558;
wire n_8373;
wire n_10848;
wire n_13165;
wire n_17412;
wire n_17704;
wire n_6481;
wire n_15926;
wire n_5628;
wire n_7765;
wire n_11482;
wire n_7816;
wire n_12151;
wire n_16943;
wire n_15201;
wire n_17407;
wire n_11089;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_13422;
wire n_15809;
wire n_15204;
wire n_6384;
wire n_7421;
wire n_15579;
wire n_18549;
wire n_13828;
wire n_10166;
wire n_7489;
wire n_7541;
wire n_6906;
wire n_18084;
wire n_14702;
wire n_13179;
wire n_14562;
wire n_15585;
wire n_5251;
wire n_15844;
wire n_12033;
wire n_11839;
wire n_18039;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_14376;
wire n_13834;
wire n_18277;
wire n_10366;
wire n_18284;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_17800;
wire n_11365;
wire n_18138;
wire n_17016;
wire n_17613;
wire n_9595;
wire n_7188;
wire n_15015;
wire n_16081;
wire n_5475;
wire n_11217;
wire n_15651;
wire n_15555;
wire n_15341;
wire n_7334;
wire n_17759;
wire n_6923;
wire n_5807;
wire n_13923;
wire n_9287;
wire n_7991;
wire n_15477;
wire n_13051;
wire n_16376;
wire n_6233;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_16737;
wire n_17220;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_14991;
wire n_17959;
wire n_14686;
wire n_12214;
wire n_10225;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_16259;
wire n_8926;
wire n_6257;
wire n_11228;
wire n_10361;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_8383;
wire n_10086;
wire n_5439;
wire n_7143;
wire n_18286;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_13924;
wire n_8965;
wire n_11290;
wire n_17080;
wire n_5936;
wire n_12518;
wire n_9608;
wire n_7646;
wire n_14047;
wire n_9052;
wire n_13476;
wire n_18454;
wire n_8817;
wire n_8190;
wire n_11488;
wire n_17447;
wire n_18399;
wire n_13671;
wire n_12162;
wire n_17537;
wire n_17678;
wire n_6587;
wire n_14627;
wire n_14876;
wire n_6987;
wire n_7781;
wire n_18265;
wire n_7360;
wire n_11037;
wire n_14568;
wire n_16925;
wire n_11702;
wire n_6069;
wire n_13699;
wire n_14319;
wire n_16970;
wire n_7497;
wire n_17087;
wire n_11372;
wire n_5706;
wire n_7665;
wire n_16763;
wire n_9354;
wire n_10817;
wire n_10501;
wire n_11829;
wire n_14026;
wire n_15324;
wire n_18437;
wire n_11517;
wire n_17782;
wire n_7793;
wire n_16102;
wire n_17462;
wire n_16274;
wire n_8355;
wire n_6991;
wire n_10556;
wire n_15287;
wire n_17098;
wire n_12741;
wire n_18041;
wire n_7101;
wire n_7671;
wire n_9436;
wire n_7530;
wire n_8489;
wire n_13150;
wire n_15006;
wire n_18157;
wire n_13776;
wire n_5431;
wire n_15103;
wire n_15619;
wire n_7248;
wire n_10350;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_15835;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_14818;
wire n_13343;
wire n_7654;
wire n_16123;
wire n_13152;
wire n_8303;
wire n_17221;
wire n_6153;
wire n_6637;
wire n_8369;
wire n_9238;
wire n_9022;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_18364;
wire n_17339;
wire n_6633;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_9103;
wire n_11665;
wire n_5774;
wire n_6579;
wire n_11031;
wire n_13590;
wire n_13907;
wire n_17142;
wire n_16747;
wire n_5798;
wire n_11138;
wire n_11731;
wire n_17365;
wire n_5875;
wire n_5187;
wire n_9839;
wire n_12821;
wire n_14782;
wire n_18479;
wire n_16257;
wire n_8831;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_15704;
wire n_6569;
wire n_7120;
wire n_8728;
wire n_6335;
wire n_10807;
wire n_12837;
wire n_12478;
wire n_12233;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_17265;
wire n_8853;
wire n_14070;
wire n_14330;
wire n_15327;
wire n_17718;
wire n_13491;
wire n_6252;
wire n_13545;
wire n_13471;
wire n_13760;
wire n_17615;
wire n_18403;
wire n_13883;
wire n_6211;
wire n_15716;
wire n_10511;
wire n_5844;
wire n_8862;
wire n_15748;
wire n_17499;
wire n_16161;
wire n_10580;
wire n_17287;
wire n_14235;
wire n_17172;
wire n_17898;
wire n_17995;
wire n_6164;
wire n_13261;
wire n_7576;
wire n_8081;
wire n_6173;
wire n_9675;
wire n_14851;
wire n_16608;
wire n_17310;
wire n_18012;
wire n_7786;
wire n_11023;
wire n_7313;
wire n_10058;
wire n_16471;
wire n_16923;
wire n_10873;
wire n_14484;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_11454;
wire n_13442;
wire n_8900;
wire n_12523;
wire n_14444;
wire n_17539;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_10484;
wire n_18531;
wire n_6737;
wire n_11744;
wire n_17247;
wire n_18388;
wire n_15726;
wire n_8396;
wire n_16560;
wire n_6612;
wire n_14307;
wire n_8478;
wire n_6606;
wire n_13450;
wire n_16988;
wire n_6695;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_15302;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_14178;
wire n_11626;
wire n_12148;
wire n_15299;
wire n_11072;
wire n_5867;
wire n_17475;
wire n_16872;
wire n_5508;
wire n_17363;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_12907;
wire n_16312;
wire n_15500;
wire n_8497;
wire n_10770;
wire n_16204;
wire n_8820;
wire n_6410;
wire n_14891;
wire n_16793;
wire n_17051;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_5597;
wire n_9028;
wire n_13944;
wire n_17217;
wire n_17873;
wire n_9492;
wire n_15592;
wire n_8020;
wire n_6090;
wire n_6413;
wire n_16064;
wire n_16443;
wire n_18524;
wire n_9374;
wire n_7419;
wire n_15319;
wire n_6506;
wire n_18456;
wire n_18476;
wire n_5515;
wire n_5662;
wire n_18123;
wire n_13634;
wire n_18281;
wire n_12132;
wire n_17086;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_18027;
wire n_10593;
wire n_13019;
wire n_14452;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_16801;
wire n_17894;
wire n_13464;
wire n_18343;
wire n_12670;
wire n_12182;
wire n_10636;
wire n_12043;
wire n_16817;
wire n_18336;
wire n_17786;
wire n_7667;
wire n_16478;
wire n_5697;
wire n_18489;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_15369;
wire n_8992;
wire n_15134;
wire n_17835;
wire n_12708;
wire n_16110;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_6234;
wire n_6821;
wire n_17459;
wire n_5462;
wire n_9983;
wire n_9375;
wire n_10082;
wire n_17715;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_7182;
wire n_15453;
wire n_5318;
wire n_7365;
wire n_13573;
wire n_6608;
wire n_10467;
wire n_9109;
wire n_9849;
wire n_13622;
wire n_6105;
wire n_6022;
wire n_11207;
wire n_17476;
wire n_9856;
wire n_10964;
wire n_18449;
wire n_16951;
wire n_5498;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_17591;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_14794;
wire n_17684;
wire n_9237;
wire n_13931;
wire n_11668;
wire n_7885;
wire n_15208;
wire n_15684;
wire n_6860;
wire n_6557;
wire n_14404;
wire n_8466;
wire n_18302;
wire n_6753;
wire n_12137;
wire n_18164;
wire n_6527;
wire n_16720;
wire n_17151;
wire n_7341;
wire n_11328;
wire n_9349;
wire n_12306;
wire n_15275;
wire n_17423;
wire n_11200;
wire n_12088;
wire n_14442;
wire n_15210;
wire n_15423;
wire n_11091;
wire n_8094;
wire n_10940;
wire n_14377;
wire n_16463;
wire n_15976;
wire n_16536;
wire n_6639;
wire n_12096;
wire n_12508;
wire n_6430;
wire n_13418;
wire n_18100;
wire n_18268;
wire n_8832;
wire n_10987;
wire n_17723;
wire n_5477;
wire n_12684;
wire n_8839;
wire n_5175;
wire n_7996;
wire n_12891;
wire n_11098;
wire n_15815;
wire n_11615;
wire n_10533;
wire n_11059;
wire n_5987;
wire n_16403;
wire n_5179;
wire n_7957;
wire n_14616;
wire n_11965;
wire n_16799;
wire n_10938;
wire n_16681;
wire n_10176;
wire n_7517;
wire n_6627;
wire n_8080;
wire n_14696;
wire n_17147;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_17965;
wire n_7745;
wire n_12941;
wire n_14006;
wire n_13551;
wire n_6666;
wire n_18019;
wire n_10927;
wire n_14258;
wire n_12200;
wire n_8321;
wire n_16060;
wire n_14024;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_11722;
wire n_8592;
wire n_8786;
wire n_15597;
wire n_17212;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_13682;
wire n_6249;
wire n_16920;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_9805;
wire n_10155;
wire n_5480;
wire n_16199;
wire n_13593;
wire n_8157;
wire n_7095;
wire n_11461;
wire n_13902;
wire n_10714;
wire n_11701;
wire n_16672;
wire n_6969;
wire n_7459;
wire n_6615;
wire n_6161;
wire n_17331;
wire n_7294;
wire n_8206;
wire n_9110;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_8622;
wire n_18338;
wire n_18010;
wire n_18358;
wire n_5904;
wire n_13917;
wire n_15367;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_9335;
wire n_13546;
wire n_14595;
wire n_17001;
wire n_14468;
wire n_7908;
wire n_6062;
wire n_12550;
wire n_9452;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_13350;
wire n_13861;
wire n_10051;
wire n_8104;
wire n_10414;
wire n_11255;
wire n_8344;
wire n_17597;
wire n_13592;
wire n_17428;
wire n_17224;
wire n_5284;
wire n_11720;
wire n_18511;
wire n_12673;
wire n_14694;
wire n_8120;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_9075;
wire n_12961;
wire n_13874;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_10746;
wire n_12225;
wire n_17817;
wire n_9188;
wire n_6294;
wire n_16407;
wire n_18009;
wire n_9611;
wire n_15506;
wire n_18371;
wire n_9021;
wire n_8779;
wire n_9810;
wire n_14469;
wire n_16269;
wire n_8621;
wire n_5503;
wire n_9250;
wire n_5845;
wire n_5945;
wire n_11212;
wire n_9550;
wire n_12884;
wire n_13145;
wire n_16591;
wire n_10697;
wire n_11714;
wire n_16201;
wire n_16179;
wire n_11263;
wire n_10641;
wire n_6246;
wire n_8868;
wire n_15070;
wire n_17690;
wire n_8134;
wire n_12207;
wire n_9975;
wire n_7250;
wire n_5755;
wire n_5600;
wire n_16566;
wire n_8762;
wire n_12011;
wire n_13195;
wire n_8043;
wire n_8694;
wire n_16377;
wire n_17503;
wire n_14492;
wire n_13965;
wire n_18365;
wire n_17358;
wire n_6053;
wire n_11994;
wire n_7252;
wire n_13419;
wire n_9207;
wire n_13358;
wire n_14134;
wire n_11860;
wire n_17057;
wire n_11990;
wire n_16693;
wire n_10103;
wire n_5245;
wire n_6843;
wire n_10926;
wire n_14519;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_16125;
wire n_10626;
wire n_15457;
wire n_6901;
wire n_14345;
wire n_13273;
wire n_11503;
wire n_16847;
wire n_8191;
wire n_17104;
wire n_10325;
wire n_6841;
wire n_10153;
wire n_17622;
wire n_16354;
wire n_17952;
wire n_8101;
wire n_10298;
wire n_8376;
wire n_8171;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_18271;
wire n_16701;
wire n_7698;
wire n_5749;
wire n_6774;
wire n_12854;
wire n_15640;
wire n_6271;
wire n_16964;
wire n_6489;
wire n_8600;
wire n_16427;
wire n_7402;
wire n_8431;
wire n_14816;
wire n_8710;
wire n_15683;
wire n_12806;
wire n_16336;
wire n_16202;
wire n_16248;
wire n_14302;
wire n_8599;
wire n_8549;
wire n_13460;
wire n_15451;
wire n_10172;
wire n_8054;
wire n_5993;
wire n_11273;
wire n_13904;
wire n_16614;
wire n_10400;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_6020;
wire n_16954;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_14035;
wire n_17045;
wire n_14496;
wire n_14467;
wire n_13218;
wire n_9096;
wire n_9081;
wire n_13952;
wire n_11697;
wire n_14789;
wire n_15784;
wire n_13076;
wire n_15526;
wire n_11762;
wire n_9236;
wire n_6844;
wire n_11969;
wire n_12950;
wire n_16963;
wire n_7914;
wire n_8628;
wire n_16388;
wire n_6521;
wire n_7891;
wire n_18074;
wire n_13028;
wire n_14413;
wire n_15150;
wire n_8857;
wire n_8517;
wire n_14243;
wire n_8547;
wire n_10156;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_6162;
wire n_10433;
wire n_6779;
wire n_8010;
wire n_6432;
wire n_9116;
wire n_14096;
wire n_10774;
wire n_12332;
wire n_10901;
wire n_11034;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_7216;
wire n_12762;
wire n_13574;
wire n_15990;
wire n_11499;
wire n_15364;
wire n_10825;
wire n_14583;
wire n_14893;
wire n_16740;
wire n_8275;
wire n_6198;
wire n_17292;
wire n_5418;
wire n_6543;
wire n_18270;
wire n_9830;
wire n_6762;
wire n_18023;
wire n_6178;
wire n_9621;
wire n_5685;
wire n_10761;
wire n_14777;
wire n_18075;
wire n_16117;
wire n_14057;
wire n_5459;
wire n_9035;
wire n_11579;
wire n_10398;
wire n_15303;
wire n_17788;
wire n_8291;
wire n_18017;
wire n_16960;
wire n_17947;
wire n_16459;
wire n_11535;
wire n_17987;
wire n_17942;
wire n_15661;
wire n_16406;
wire n_18165;
wire n_12558;
wire n_14915;
wire n_17932;
wire n_17780;
wire n_18400;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_7477;
wire n_5173;
wire n_17028;
wire n_15654;
wire n_17075;
wire n_12975;
wire n_17289;
wire n_11402;
wire n_6458;
wire n_7642;
wire n_9678;
wire n_11401;
wire n_17828;
wire n_8247;
wire n_17820;
wire n_6577;
wire n_12506;
wire n_16291;
wire n_18356;
wire n_13850;
wire n_6740;
wire n_12718;
wire n_12956;
wire n_17373;
wire n_11510;
wire n_6315;
wire n_10581;
wire n_12638;
wire n_14116;
wire n_14856;
wire n_15235;
wire n_14949;
wire n_17487;
wire n_17866;
wire n_9284;
wire n_12736;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_9163;
wire n_18372;
wire n_15461;
wire n_12086;
wire n_15711;
wire n_16453;
wire n_16645;
wire n_5170;
wire n_6910;
wire n_7604;
wire n_6262;
wire n_14800;
wire n_16952;
wire n_7703;
wire n_9606;
wire n_6319;
wire n_17352;
wire n_17018;
wire n_13459;
wire n_10470;
wire n_16449;
wire n_14268;
wire n_11589;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_14888;
wire n_15034;
wire n_12350;
wire n_16775;
wire n_12542;
wire n_13860;
wire n_5839;
wire n_14240;
wire n_14504;
wire n_18266;
wire n_13449;
wire n_14127;
wire n_6536;
wire n_12747;
wire n_6175;
wire n_7040;
wire n_8827;
wire n_10625;
wire n_16606;
wire n_8280;
wire n_12561;
wire n_12390;
wire n_14460;
wire n_5514;
wire n_13216;
wire n_18420;
wire n_8388;
wire n_18469;
wire n_12849;
wire n_14730;
wire n_10235;
wire n_11312;
wire n_6978;
wire n_17937;
wire n_13786;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_10445;
wire n_15110;
wire n_16306;
wire n_7378;
wire n_10738;
wire n_14894;
wire n_12866;
wire n_17801;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_15491;
wire n_15025;
wire n_18485;
wire n_9190;
wire n_14925;
wire n_6947;
wire n_11612;
wire n_9482;
wire n_14918;
wire n_5293;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_18161;
wire n_12900;
wire n_13414;
wire n_8569;
wire n_5400;
wire n_14598;
wire n_6140;
wire n_8877;
wire n_15489;
wire n_9412;
wire n_7498;
wire n_10679;
wire n_11323;
wire n_10799;
wire n_15561;
wire n_6321;
wire n_12914;
wire n_17159;
wire n_11916;
wire n_6819;
wire n_7501;
wire n_9506;
wire n_5201;
wire n_10136;
wire n_18440;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_17228;
wire n_10585;
wire n_18519;
wire n_12764;
wire n_13696;
wire n_15148;
wire n_15325;
wire n_11356;
wire n_16457;
wire n_16542;
wire n_15955;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_13322;
wire n_15158;
wire n_14238;
wire n_9092;
wire n_10034;
wire n_16918;
wire n_9451;
wire n_11148;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_13934;
wire n_6899;
wire n_15389;
wire n_7549;
wire n_10692;
wire n_17054;
wire n_17308;
wire n_7373;
wire n_17425;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_14826;
wire n_15331;
wire n_15776;
wire n_16019;
wire n_16421;
wire n_17109;
wire n_17732;
wire n_6592;
wire n_11280;
wire n_12337;
wire n_13254;
wire n_14987;
wire n_13466;
wire n_15082;
wire n_15191;
wire n_18520;
wire n_8686;
wire n_17617;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_11114;
wire n_15676;
wire n_9011;
wire n_17044;
wire n_16023;
wire n_17641;
wire n_8418;
wire n_7740;
wire n_8403;
wire n_5891;
wire n_13050;
wire n_14042;
wire n_7613;
wire n_11493;
wire n_9220;
wire n_6101;
wire n_17312;
wire n_14440;
wire n_17742;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_10860;
wire n_18259;
wire n_12763;
wire n_17517;
wire n_16208;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_5623;
wire n_15209;
wire n_15269;
wire n_18460;
wire n_12273;
wire n_13875;
wire n_17272;
wire n_17319;
wire n_16394;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_17774;
wire n_15310;
wire n_17989;
wire n_12712;
wire n_14076;
wire n_11220;
wire n_17709;
wire n_9012;
wire n_15078;
wire n_13012;
wire n_8698;
wire n_8924;
wire n_12584;
wire n_14435;
wire n_14638;
wire n_18150;
wire n_14946;
wire n_10376;
wire n_15510;
wire n_12752;
wire n_15674;
wire n_7515;
wire n_6928;
wire n_10880;
wire n_15511;
wire n_17567;
wire n_7238;
wire n_9994;
wire n_14226;
wire n_17933;
wire n_8780;
wire n_7309;
wire n_15811;
wire n_17384;
wire n_14936;
wire n_7958;
wire n_16469;
wire n_18037;
wire n_8047;
wire n_11596;
wire n_18204;
wire n_8559;
wire n_5693;
wire n_6273;
wire n_14278;
wire n_11885;
wire n_17670;
wire n_15618;
wire n_7572;
wire n_5663;
wire n_11955;
wire n_8214;
wire n_10224;
wire n_12777;
wire n_14706;
wire n_15849;
wire n_5990;
wire n_7043;
wire n_10777;
wire n_11462;
wire n_11732;
wire n_16490;
wire n_16156;
wire n_9391;
wire n_7760;
wire n_16105;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_13306;
wire n_12819;
wire n_14159;
wire n_14515;
wire n_18137;
wire n_8722;
wire n_16489;
wire n_11654;
wire n_12268;
wire n_16900;
wire n_10214;
wire n_8589;
wire n_8241;
wire n_18361;
wire n_12077;
wire n_12982;
wire n_7573;
wire n_8442;
wire n_15321;
wire n_6281;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_14757;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_6311;
wire n_10469;
wire n_9229;
wire n_11194;
wire n_11480;
wire n_15282;
wire n_16812;
wire n_16038;
wire n_7590;
wire n_9342;
wire n_18062;
wire n_12237;
wire n_13271;
wire n_18350;
wire n_6134;
wire n_9329;
wire n_5426;
wire n_10175;
wire n_11481;
wire n_5803;
wire n_13372;
wire n_15812;
wire n_16292;
wire n_9868;
wire n_11375;
wire n_17119;
wire n_5285;
wire n_18458;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_9311;
wire n_12275;
wire n_6593;
wire n_13742;
wire n_8630;
wire n_17019;
wire n_15177;
wire n_16491;
wire n_12376;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_8145;
wire n_8405;
wire n_10447;
wire n_9260;
wire n_15063;
wire n_7176;
wire n_14534;
wire n_8928;
wire n_17638;
wire n_13630;
wire n_7682;
wire n_15223;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_16535;
wire n_11925;
wire n_13700;
wire n_18584;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_10406;
wire n_5715;
wire n_12509;
wire n_14902;
wire n_16033;
wire n_8295;
wire n_6932;
wire n_17859;
wire n_6746;
wire n_11985;
wire n_13527;
wire n_8447;
wire n_7901;
wire n_5395;
wire n_10522;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_6446;
wire n_16618;
wire n_10278;
wire n_14290;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_6996;
wire n_7218;
wire n_8828;
wire n_9430;
wire n_15935;
wire n_17674;
wire n_15384;
wire n_17687;
wire n_11407;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_12710;
wire n_15686;
wire n_6749;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_7005;
wire n_15950;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_18098;
wire n_10798;
wire n_10965;
wire n_17182;
wire n_7732;
wire n_13325;
wire n_6337;
wire n_14850;
wire n_6181;
wire n_15135;
wire n_16196;
wire n_7447;
wire n_9776;
wire n_18212;
wire n_17998;
wire n_16736;
wire n_11911;
wire n_6777;
wire n_18156;
wire n_11987;
wire n_18208;
wire n_11442;
wire n_8227;
wire n_12936;
wire n_12721;
wire n_18301;
wire n_5634;
wire n_18424;
wire n_5672;
wire n_16008;
wire n_8475;
wire n_11730;
wire n_10482;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_18527;
wire n_14064;
wire n_14524;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_16883;
wire n_7405;
wire n_12039;
wire n_11651;
wire n_11388;
wire n_14151;
wire n_8314;
wire n_9386;
wire n_15120;
wire n_10154;
wire n_5617;
wire n_17946;
wire n_7922;
wire n_13089;
wire n_17469;
wire n_15826;
wire n_15459;
wire n_15192;
wire n_10377;
wire n_5266;
wire n_5580;
wire n_18360;
wire n_9926;
wire n_10033;
wire n_11121;
wire n_13167;
wire n_16836;
wire n_11270;
wire n_17877;
wire n_12329;
wire n_6310;
wire n_15161;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_8311;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_5310;
wire n_9661;
wire n_16303;
wire n_9843;
wire n_15013;
wire n_9877;
wire n_8764;
wire n_14284;
wire n_6953;
wire n_16710;
wire n_14945;
wire n_16559;
wire n_5722;
wire n_13001;
wire n_5390;
wire n_13232;
wire n_9901;
wire n_16167;
wire n_17377;
wire n_17334;
wire n_13320;
wire n_5593;
wire n_12990;
wire n_18348;
wire n_14246;
wire n_6683;
wire n_10683;
wire n_18487;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_16353;
wire n_6365;
wire n_6920;
wire n_9921;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_8567;
wire n_11817;
wire n_13278;
wire n_15455;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_5237;
wire n_13597;
wire n_14957;
wire n_13488;
wire n_11042;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_13447;
wire n_15907;
wire n_7089;
wire n_7144;
wire n_16534;
wire n_7286;
wire n_16579;
wire n_18232;
wire n_11479;
wire n_11737;
wire n_8048;
wire n_14681;
wire n_12028;
wire n_13668;
wire n_7072;
wire n_13016;
wire n_11272;
wire n_14230;
wire n_13095;
wire n_8253;
wire n_6177;
wire n_16961;
wire n_14708;
wire n_6332;
wire n_17293;
wire n_5853;
wire n_12048;
wire n_18592;
wire n_15032;
wire n_8283;
wire n_5982;
wire n_10930;
wire n_11600;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_17972;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_17855;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_14546;
wire n_18264;
wire n_7129;
wire n_13938;
wire n_12057;
wire n_6696;
wire n_15440;
wire n_13251;
wire n_17590;
wire n_9882;
wire n_9527;
wire n_16484;
wire n_8566;
wire n_16450;
wire n_7343;
wire n_14875;
wire n_12766;
wire n_15860;
wire n_8516;
wire n_10637;
wire n_8302;
wire n_15056;
wire n_8317;
wire n_17288;
wire n_17717;
wire n_5376;
wire n_15610;
wire n_12229;
wire n_14003;
wire n_16197;
wire n_9205;
wire n_6116;
wire n_9511;
wire n_8167;
wire n_15329;
wire n_7859;
wire n_14315;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_17822;
wire n_13670;
wire n_17464;
wire n_7972;
wire n_11254;
wire n_13319;
wire n_15023;
wire n_11617;
wire n_13858;
wire n_13512;
wire n_9071;
wire n_7916;
wire n_17913;
wire n_9368;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_10415;
wire n_13069;
wire n_18184;
wire n_11711;
wire n_5410;
wire n_12362;
wire n_8944;
wire n_6167;
wire n_15666;
wire n_16255;
wire n_13233;
wire n_11931;
wire n_8008;
wire n_18495;
wire n_10023;
wire n_18436;
wire n_10999;
wire n_6170;
wire n_8109;
wire n_13297;
wire n_9459;
wire n_14185;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_6307;
wire n_10410;
wire n_6094;
wire n_9098;
wire n_7987;
wire n_7483;
wire n_14953;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_14873;
wire n_15604;
wire n_7434;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_9504;
wire n_15359;
wire n_16983;
wire n_14840;
wire n_8975;
wire n_16556;
wire n_6267;
wire n_16000;
wire n_9063;
wire n_7787;
wire n_12360;
wire n_5998;
wire n_9268;
wire n_17116;
wire n_15431;
wire n_5304;
wire n_17861;
wire n_17009;
wire n_6568;
wire n_15035;
wire n_18500;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_18038;
wire n_17668;
wire n_18536;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_10456;
wire n_15631;
wire n_16072;
wire n_6261;
wire n_14083;
wire n_13186;
wire n_5916;
wire n_11907;
wire n_15655;
wire n_10096;
wire n_13617;
wire n_10627;
wire n_10025;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_14755;
wire n_6299;
wire n_6813;
wire n_8825;
wire n_12969;
wire n_15430;
wire n_11753;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_15732;
wire n_8266;
wire n_5691;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_8981;
wire n_8420;
wire n_17082;
wire n_17616;
wire n_8297;
wire n_11150;
wire n_18199;
wire n_8771;
wire n_17772;
wire n_10881;
wire n_13519;
wire n_16111;
wire n_15750;
wire n_14170;
wire n_16583;
wire n_15641;
wire n_13496;
wire n_16007;
wire n_12939;
wire n_17129;
wire n_6316;
wire n_15038;
wire n_6292;
wire n_17925;
wire n_9726;
wire n_13884;
wire n_10404;
wire n_8639;
wire n_8138;
wire n_8058;
wire n_9308;
wire n_6638;
wire n_12779;
wire n_16796;
wire n_11838;
wire n_10508;
wire n_16510;
wire n_17125;
wire n_17505;
wire n_18008;
wire n_7719;
wire n_15892;
wire n_10811;
wire n_14049;
wire n_8333;
wire n_17199;
wire n_5615;
wire n_6220;
wire n_7562;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_7619;
wire n_6985;
wire n_17152;
wire n_12783;
wire n_7170;
wire n_13853;
wire n_9211;
wire n_12019;
wire n_8176;
wire n_8124;
wire n_14529;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_16106;
wire n_5269;
wire n_10891;
wire n_17348;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_15284;
wire n_10803;
wire n_8147;
wire n_13190;
wire n_5468;
wire n_6188;
wire n_17671;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_14195;
wire n_18363;
wire n_5262;
wire n_10700;
wire n_17743;
wire n_7938;
wire n_10968;
wire n_11695;
wire n_17595;
wire n_7935;
wire n_8458;
wire n_5421;
wire n_14247;
wire n_6772;
wire n_16902;
wire n_8113;
wire n_9716;
wire n_16646;
wire n_15877;
wire n_14300;
wire n_11453;
wire n_16155;
wire n_15443;
wire n_5206;
wire n_17901;
wire n_6077;
wire n_17896;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_6318;
wire n_15418;
wire n_16445;
wire n_11970;
wire n_16997;
wire n_18228;
wire n_17090;
wire n_14678;
wire n_17833;
wire n_7918;
wire n_13599;
wire n_17282;
wire n_18471;
wire n_13354;
wire n_14690;
wire n_17356;
wire n_15008;
wire n_16852;
wire n_5188;
wire n_13647;
wire n_6916;
wire n_15524;
wire n_13683;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_10783;
wire n_10147;
wire n_11862;
wire n_12163;
wire n_17921;
wire n_14839;
wire n_10725;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_17197;
wire n_18354;
wire n_12944;
wire n_15409;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_16207;
wire n_18503;
wire n_9433;
wire n_9737;
wire n_18568;
wire n_9298;
wire n_11660;
wire n_18058;
wire n_10812;
wire n_14709;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_14249;
wire n_16939;
wire n_18152;
wire n_6230;
wire n_14241;
wire n_6604;
wire n_14497;
wire n_16108;
wire n_5373;
wire n_10001;
wire n_16101;
wire n_11107;
wire n_14280;
wire n_13724;
wire n_13280;
wire n_9301;
wire n_12145;
wire n_11088;
wire n_5573;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_8160;
wire n_6391;
wire n_10284;
wire n_12757;
wire n_12054;
wire n_15827;
wire n_14379;
wire n_5659;
wire n_8099;
wire n_14446;
wire n_17256;
wire n_11595;
wire n_8840;
wire n_16284;
wire n_11405;
wire n_14719;
wire n_16001;
wire n_15575;
wire n_17806;
wire n_13768;
wire n_13189;
wire n_5881;
wire n_16707;
wire n_8522;
wire n_12971;
wire n_7222;
wire n_7942;
wire n_8578;
wire n_6473;
wire n_13103;
wire n_13838;
wire n_15630;
wire n_16599;
wire n_18385;
wire n_10046;
wire n_15696;
wire n_12328;
wire n_14558;
wire n_11318;
wire n_9083;
wire n_7725;
wire n_10977;
wire n_16950;
wire n_17198;
wire n_11299;
wire n_10397;
wire n_6483;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_14004;
wire n_17023;
wire n_5863;
wire n_7647;
wire n_8626;
wire n_10936;
wire n_12442;
wire n_16221;
wire n_8611;
wire n_8036;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_17927;
wire n_16222;
wire n_15123;
wire n_9835;
wire n_15068;
wire n_15442;
wire n_7300;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_14666;
wire n_13605;
wire n_17387;
wire n_10532;
wire n_17776;
wire n_5466;
wire n_13995;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_13441;
wire n_6728;
wire n_6729;
wire n_14237;
wire n_16082;
wire n_15095;
wire n_11240;
wire n_10207;
wire n_13857;
wire n_13841;
wire n_16029;
wire n_13556;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_13367;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_17737;
wire n_10771;
wire n_17166;
wire n_13816;
wire n_11487;
wire n_18355;
wire n_11441;
wire n_8441;
wire n_16119;
wire n_14203;
wire n_6076;
wire n_8933;
wire n_17269;
wire n_15876;
wire n_17215;
wire n_7778;
wire n_15231;
wire n_12844;
wire n_5851;
wire n_14736;
wire n_7073;
wire n_9755;
wire n_11287;
wire n_9774;
wire n_8397;
wire n_6390;
wire n_10139;
wire n_13409;
wire n_13246;
wire n_14061;
wire n_5796;
wire n_10104;
wire n_8726;
wire n_17916;
wire n_12986;
wire n_11381;
wire n_6665;
wire n_16378;
wire n_17250;
wire n_16109;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_9117;
wire n_16172;
wire n_9720;
wire n_16611;
wire n_7746;
wire n_9381;
wire n_10169;
wire n_15727;
wire n_6958;
wire n_16277;
wire n_16598;
wire n_12049;
wire n_12690;
wire n_14498;
wire n_15417;
wire n_7563;
wire n_12475;
wire n_17588;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_6653;
wire n_16806;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_14713;
wire n_15512;
wire n_7853;
wire n_12526;
wire n_14414;
wire n_15565;
wire n_7531;
wire n_12377;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_18486;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_16575;
wire n_13650;
wire n_16789;
wire n_7721;
wire n_7192;
wire n_14202;
wire n_15636;
wire n_15859;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_14554;
wire n_9887;
wire n_9149;
wire n_15946;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_15807;
wire n_13211;
wire n_18063;
wire n_8316;
wire n_16858;
wire n_16980;
wire n_9990;
wire n_5829;
wire n_10005;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_5191;
wire n_14874;
wire n_15311;
wire n_8505;
wire n_15113;
wire n_17258;
wire n_9273;
wire n_18198;
wire n_17667;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_15498;
wire n_8970;
wire n_17315;
wire n_16910;
wire n_7527;
wire n_7417;
wire n_13061;
wire n_9682;
wire n_18550;
wire n_18097;
wire n_12513;
wire n_17719;
wire n_10640;
wire n_16824;
wire n_6582;
wire n_5734;
wire n_15098;
wire n_13395;
wire n_10729;
wire n_12545;
wire n_18432;
wire n_14656;
wire n_16832;
wire n_7388;
wire n_16052;
wire n_18320;
wire n_11657;
wire n_18078;
wire n_9924;
wire n_14745;
wire n_8717;
wire n_14744;
wire n_13336;
wire n_5770;
wire n_5705;
wire n_16074;
wire n_15091;
wire n_9064;
wire n_7635;
wire n_17420;
wire n_5525;
wire n_13102;
wire n_11268;
wire n_17121;
wire n_12753;
wire n_17527;
wire n_14760;
wire n_18108;
wire n_7090;
wire n_9254;
wire n_12894;
wire n_14135;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_16482;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_13390;
wire n_13691;
wire n_13375;
wire n_15769;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_8030;
wire n_18526;
wire n_9247;
wire n_17340;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_16809;
wire n_16913;
wire n_14194;
wire n_10526;
wire n_8725;
wire n_5575;
wire n_12010;
wire n_9738;
wire n_5675;
wire n_9570;
wire n_12026;
wire n_16663;
wire n_12356;
wire n_11857;
wire n_13825;
wire n_11077;
wire n_6240;
wire n_8243;
wire n_17481;
wire n_8633;
wire n_6347;
wire n_9593;
wire n_9846;
wire n_7689;
wire n_13262;
wire n_13482;
wire n_17645;
wire n_6511;
wire n_18069;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_18470;
wire n_9469;
wire n_10764;
wire n_15869;
wire n_18005;
wire n_18429;
wire n_13398;
wire n_9677;
wire n_15598;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_14676;
wire n_8449;
wire n_17605;
wire n_6358;
wire n_13204;
wire n_14331;
wire n_6603;
wire n_17812;
wire n_16604;
wire n_13873;
wire n_15805;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_8201;
wire n_8967;
wire n_6986;
wire n_8801;
wire n_9322;
wire n_10438;
wire n_15017;
wire n_5959;
wire n_11201;
wire n_16485;
wire n_10531;
wire n_14964;
wire n_8918;
wire n_8031;
wire n_15591;
wire n_12878;
wire n_9348;
wire n_14262;
wire n_16438;
wire n_12188;
wire n_8219;
wire n_15373;
wire n_16609;
wire n_8696;
wire n_18580;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_15167;
wire n_12630;
wire n_17756;
wire n_6890;
wire n_11028;
wire n_12171;
wire n_12299;
wire n_16739;
wire n_16603;
wire n_15706;
wire n_12022;
wire n_9249;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_17271;
wire n_8180;
wire n_10741;
wire n_15211;
wire n_18207;
wire n_6109;
wire n_14727;
wire n_10760;
wire n_15580;
wire n_12425;
wire n_14762;
wire n_9444;
wire n_15334;
wire n_7731;
wire n_10772;
wire n_11527;
wire n_7114;
wire n_13507;
wire n_18404;
wire n_16486;
wire n_11327;
wire n_10915;
wire n_9535;
wire n_18290;
wire n_15984;
wire n_6770;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_15900;
wire n_12199;
wire n_17133;
wire n_5302;
wire n_12000;
wire n_17730;
wire n_17729;
wire n_15410;
wire n_9707;
wire n_12490;
wire n_15151;
wire n_16002;
wire n_16626;
wire n_16258;
wire n_13594;
wire n_17281;
wire n_5639;
wire n_5781;
wire n_17547;
wire n_14182;
wire n_8943;
wire n_8486;
wire n_14767;
wire n_10279;
wire n_18463;
wire n_15853;
wire n_5299;
wire n_12829;
wire n_14352;
wire n_13889;
wire n_14773;
wire n_10680;
wire n_10127;
wire n_5543;
wire n_17864;
wire n_13654;
wire n_5361;
wire n_11610;
wire n_7081;
wire n_7132;
wire n_11814;
wire n_12255;
wire n_12739;
wire n_13015;
wire n_17021;
wire n_5885;
wire n_6663;
wire n_17710;
wire n_14228;
wire n_12609;
wire n_9723;
wire n_5356;
wire n_7319;
wire n_18248;
wire n_15831;
wire n_5458;
wire n_7644;
wire n_11176;
wire n_16131;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_11360;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5330;
wire n_7199;
wire n_10039;
wire n_11726;
wire n_10854;
wire n_11358;
wire n_5463;
wire n_15944;
wire n_13366;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_12904;
wire n_8833;
wire n_9191;
wire n_5489;
wire n_7828;
wire n_5892;
wire n_10142;
wire n_14623;
wire n_7940;
wire n_17791;
wire n_9918;
wire n_15932;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_16467;
wire n_6009;
wire n_18202;
wire n_9034;
wire n_16345;
wire n_17669;
wire n_6503;
wire n_6376;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_9390;
wire n_18141;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_17325;
wire n_5714;
wire n_8541;
wire n_17357;
wire n_8074;
wire n_15381;
wire n_18233;
wire n_8485;
wire n_13639;
wire n_14852;
wire n_8860;
wire n_15989;
wire n_5510;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_16103;
wire n_7001;
wire n_9650;
wire n_13070;
wire n_8271;
wire n_15514;
wire n_5692;
wire n_16460;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_9266;
wire n_14491;
wire n_12728;
wire n_5555;
wire n_15011;
wire n_10027;
wire n_16210;
wire n_12784;
wire n_17607;
wire n_16651;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_13678;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_14582;
wire n_8699;
wire n_16305;
wire n_14261;
wire n_14677;
wire n_6897;
wire n_13523;
wire n_18020;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_5366;
wire n_14928;
wire n_15550;
wire n_16016;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_15861;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_16297;
wire n_13778;
wire n_14250;
wire n_16896;
wire n_16818;
wire n_16573;
wire n_9931;
wire n_13198;
wire n_16419;
wire n_16470;
wire n_16562;
wire n_15914;
wire n_16956;
wire n_9187;
wire n_6296;
wire n_13741;
wire n_13819;
wire n_7708;
wire n_16621;
wire n_15777;
wire n_12610;
wire n_14634;
wire n_11671;
wire n_10328;
wire n_14416;
wire n_5968;
wire n_11251;
wire n_14424;
wire n_18398;
wire n_14523;
wire n_12293;
wire n_11063;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_13174;
wire n_15705;
wire n_7108;
wire n_14455;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_16816;
wire n_8368;
wire n_15691;
wire n_9259;
wire n_17560;
wire n_8322;
wire n_7333;
wire n_17164;
wire n_11879;
wire n_16127;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_15376;
wire n_16555;
wire n_17175;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_8300;
wire n_15336;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_15050;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_14161;
wire n_6573;
wire n_17767;
wire n_18112;
wire n_16760;
wire n_9656;
wire n_7634;
wire n_17488;
wire n_17427;
wire n_8148;
wire n_11400;
wire n_13290;
wire n_8150;
wire n_13500;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_15848;
wire n_15398;
wire n_10483;
wire n_15593;
wire n_16844;
wire n_18175;
wire n_17758;
wire n_12160;
wire n_11563;
wire n_9620;
wire n_16424;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_18586;
wire n_16409;
wire n_5419;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_14513;
wire n_7260;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_6409;
wire n_11939;
wire n_17145;
wire n_7954;
wire n_11119;
wire n_9824;
wire n_14347;
wire n_15089;
wire n_7951;
wire n_7552;
wire n_8096;
wire n_14602;
wire n_11468;
wire n_15995;
wire n_16150;
wire n_17969;
wire n_13901;
wire n_12166;
wire n_8233;
wire n_6130;
wire n_7273;
wire n_9683;
wire n_10646;
wire n_17403;
wire n_14750;
wire n_17939;
wire n_7231;
wire n_15725;
wire n_5976;
wire n_11704;
wire n_14074;
wire n_15252;
wire n_18043;
wire n_15132;
wire n_17506;
wire n_5732;
wire n_5372;
wire n_16238;
wire n_14050;
wire n_11878;
wire n_15843;
wire n_15763;
wire n_16666;
wire n_17983;
wire n_15749;
wire n_15317;
wire n_18050;
wire n_7449;
wire n_7772;
wire n_8763;
wire n_12800;
wire n_5208;
wire n_14197;
wire n_15638;
wire n_8679;
wire n_16547;
wire n_7239;
wire n_14289;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_16479;
wire n_16574;
wire n_11962;
wire n_15145;
wire n_5690;
wire n_9227;
wire n_17516;
wire n_18159;
wire n_8187;
wire n_10751;
wire n_16967;
wire n_7050;
wire n_10240;
wire n_17137;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_15838;
wire n_15297;
wire n_6623;
wire n_9561;
wire n_13968;
wire n_13951;
wire n_10378;
wire n_13979;
wire n_12070;
wire n_16104;
wire n_9714;
wire n_16924;
wire n_9740;
wire n_9773;
wire n_13316;
wire n_10313;
wire n_14898;
wire n_15672;
wire n_12947;
wire n_5371;
wire n_9745;
wire n_13689;
wire n_17178;
wire n_15413;
wire n_10216;
wire n_15628;
wire n_15920;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_17733;
wire n_15160;
wire n_17268;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_12354;
wire n_12666;
wire n_14395;
wire n_14297;
wire n_13528;
wire n_17388;
wire n_6047;
wire n_12581;
wire n_18000;
wire n_8292;
wire n_16368;
wire n_17395;
wire n_12631;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_8601;
wire n_10773;
wire n_18210;
wire n_18426;
wire n_6652;
wire n_9377;
wire n_11932;
wire n_10971;
wire n_18073;
wire n_8830;
wire n_6921;
wire n_6970;
wire n_5347;
wire n_14836;
wire n_13027;
wire n_18506;
wire n_12867;
wire n_7674;
wire n_14675;
wire n_9826;
wire n_12607;
wire n_14516;
wire n_15960;
wire n_7568;
wire n_15343;
wire n_6354;
wire n_7272;
wire n_18484;
wire n_15782;
wire n_12075;
wire n_11942;
wire n_15998;
wire n_6344;
wire n_12305;
wire n_13489;
wire n_12123;
wire n_9772;
wire n_12170;
wire n_15370;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_9630;
wire n_6624;
wire n_6956;
wire n_13313;
wire n_13927;
wire n_18001;
wire n_12966;
wire n_13877;
wire n_15851;
wire n_15308;
wire n_17025;
wire n_9255;
wire n_6305;
wire n_6209;
wire n_8310;
wire n_10231;
wire n_12547;
wire n_9758;
wire n_16148;
wire n_15577;
wire n_16500;
wire n_16550;
wire n_15884;
wire n_11922;
wire n_14020;
wire n_15175;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_18413;
wire n_5857;
wire n_12358;
wire n_7329;
wire n_14502;
wire n_15206;
wire n_8646;
wire n_7408;
wire n_13415;
wire n_9691;
wire n_12997;
wire n_14533;
wire n_10259;
wire n_14005;
wire n_7107;
wire n_14293;
wire n_5652;
wire n_17111;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_14334;
wire n_17951;
wire n_17379;
wire n_7690;
wire n_8969;
wire n_14187;
wire n_15245;
wire n_7123;
wire n_17935;
wire n_10752;
wire n_11577;
wire n_17840;
wire n_15225;
wire n_5499;
wire n_8117;
wire n_10067;
wire n_15169;
wire n_16914;
wire n_18021;
wire n_18513;
wire n_18528;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_13562;
wire n_14537;
wire n_12498;
wire n_17907;
wire n_13888;
wire n_16592;
wire n_11475;
wire n_6950;
wire n_8208;
wire n_17583;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_17794;
wire n_11010;
wire n_10274;
wire n_15614;
wire n_9590;
wire n_16017;
wire n_11588;
wire n_16346;
wire n_6694;
wire n_13956;
wire n_15318;
wire n_6880;
wire n_7418;
wire n_9168;
wire n_18101;
wire n_14220;
wire n_11221;
wire n_13837;
wire n_12387;
wire n_9497;
wire n_15772;
wire n_8536;
wire n_17252;
wire n_13255;
wire n_15911;
wire n_9435;
wire n_7229;
wire n_14245;
wire n_18570;
wire n_8350;
wire n_16475;
wire n_17659;
wire n_11448;
wire n_17321;
wire n_18272;
wire n_9219;
wire n_5507;
wire n_17376;
wire n_5569;
wire n_8028;
wire n_8328;
wire n_15559;
wire n_8914;
wire n_15076;
wire n_12576;
wire n_15502;
wire n_16871;
wire n_7258;
wire n_15276;
wire n_5190;
wire n_13892;
wire n_8391;
wire n_16361;
wire n_14221;
wire n_16343;
wire n_10579;
wire n_10832;
wire n_13345;
wire n_13964;
wire n_13749;
wire n_8336;
wire n_6856;
wire n_6466;
wire n_14559;
wire n_16039;
wire n_7864;
wire n_15552;
wire n_16831;
wire n_17722;
wire n_17492;
wire n_18295;
wire n_16228;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_5392;
wire n_17110;
wire n_12862;
wire n_11445;
wire n_13151;
wire n_13601;
wire n_13621;
wire n_14052;
wire n_14311;
wire n_8216;
wire n_11552;
wire n_13765;
wire n_10332;
wire n_17457;
wire n_7709;
wire n_17115;
wire n_15290;
wire n_15102;
wire n_14733;
wire n_16953;
wire n_11874;
wire n_13926;
wire n_9982;
wire n_10171;
wire n_15184;
wire n_14157;
wire n_5455;
wire n_18131;
wire n_5442;
wire n_6386;
wire n_14317;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_18155;
wire n_12656;
wire n_16220;
wire n_9852;
wire n_6820;
wire n_11623;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_5511;
wire n_6208;
wire n_5295;
wire n_17083;
wire n_6739;
wire n_15779;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_18599;
wire n_10540;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_11936;
wire n_15366;
wire n_16993;
wire n_17931;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_10200;
wire n_13392;
wire n_7332;
wire n_12734;
wire n_10382;
wire n_13164;
wire n_18247;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_17563;
wire n_11489;
wire n_13662;
wire n_10269;
wire n_8374;
wire n_12262;
wire n_13223;
wire n_16275;
wire n_17062;
wire n_13340;
wire n_9169;
wire n_14910;
wire n_13451;
wire n_13939;
wire n_5834;
wire n_10229;
wire n_17887;
wire n_17192;
wire n_5584;
wire n_13728;
wire n_7512;
wire n_14385;
wire n_7386;
wire n_17824;
wire n_9939;
wire n_7766;
wire n_10981;
wire n_8738;
wire n_11018;
wire n_14499;
wire n_18401;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_15368;
wire n_16014;
wire n_12797;
wire n_11376;
wire n_6223;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_18433;
wire n_7808;
wire n_8798;
wire n_9481;
wire n_6544;
wire n_13379;
wire n_9600;
wire n_13781;
wire n_9122;
wire n_14731;
wire n_8085;
wire n_11274;
wire n_17513;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_17081;
wire n_5707;
wire n_12012;
wire n_17997;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_16337;
wire n_9927;
wire n_14613;
wire n_5497;
wire n_10076;
wire n_17691;
wire n_11515;
wire n_17466;
wire n_8721;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_16973;
wire n_13558;
wire n_11554;
wire n_15657;
wire n_15881;
wire n_7637;
wire n_10148;
wire n_17571;
wire n_16577;
wire n_10318;
wire n_18422;
wire n_7127;
wire n_18091;
wire n_9635;
wire n_16890;
wire n_13890;
wire n_5481;
wire n_12890;
wire n_8666;
wire n_15513;
wire n_5344;
wire n_9264;
wire n_13994;
wire n_14483;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_17060;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_15724;
wire n_14308;
wire n_18322;
wire n_5408;
wire n_7801;
wire n_13484;
wire n_9155;
wire n_10234;
wire n_17298;
wire n_8460;
wire n_10416;
wire n_15837;
wire n_14370;
wire n_17468;
wire n_14593;
wire n_8836;
wire n_7959;
wire n_13430;
wire n_7019;
wire n_8181;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_8254;
wire n_13452;
wire n_13521;
wire n_8071;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_16013;
wire n_6667;
wire n_14926;
wire n_7409;
wire n_5271;
wire n_17480;
wire n_10735;
wire n_10731;
wire n_10583;
wire n_17153;
wire n_9878;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_13807;
wire n_14591;
wire n_14363;
wire n_9825;
wire n_7444;
wire n_5494;
wire n_11628;
wire n_16942;
wire n_14576;
wire n_5234;
wire n_7546;
wire n_17569;
wire n_6272;
wire n_14274;
wire n_6588;
wire n_11549;
wire n_17797;
wire n_17162;
wire n_18125;
wire n_14033;
wire n_12286;
wire n_9001;
wire n_10393;
wire n_15403;
wire n_11498;
wire n_13081;
wire n_15221;
wire n_16107;
wire n_15602;
wire n_10513;
wire n_12252;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_14545;
wire n_16090;
wire n_12627;
wire n_16743;
wire n_18031;
wire n_18467;
wire n_7575;
wire n_16730;
wire n_9045;
wire n_7083;
wire n_12281;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_9373;
wire n_15012;
wire n_14337;
wire n_6268;
wire n_16683;
wire n_17804;
wire n_5827;
wire n_12347;
wire n_14551;
wire n_5199;
wire n_17424;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_15720;
wire n_16823;
wire n_17994;
wire n_11181;
wire n_16966;
wire n_13651;
wire n_9967;
wire n_13553;
wire n_7521;
wire n_14088;
wire n_5992;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_13817;
wire n_9971;
wire n_7187;
wire n_17926;
wire n_15517;
wire n_10894;
wire n_14118;
wire n_17063;
wire n_17818;
wire n_13974;
wire n_18082;
wire n_9524;
wire n_12277;
wire n_14917;
wire n_12698;
wire n_5312;
wire n_6467;
wire n_9243;
wire n_9182;
wire n_9282;
wire n_16075;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_15680;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_9224;
wire n_10347;
wire n_16086;
wire n_5513;
wire n_5614;
wire n_17383;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_17441;
wire n_12410;
wire n_16857;
wire n_13225;
wire n_14855;
wire n_16757;
wire n_16327;
wire n_5225;
wire n_17006;
wire n_14707;
wire n_15326;
wire n_17555;
wire n_16043;
wire n_10208;
wire n_7722;
wire n_8487;
wire n_9240;
wire n_18601;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_14726;
wire n_8141;
wire n_14612;
wire n_12294;
wire n_14180;
wire n_17246;
wire n_7603;
wire n_17167;
wire n_18357;
wire n_10667;
wire n_14058;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_13355;
wire n_12957;
wire n_13141;
wire n_11616;
wire n_16461;
wire n_17688;
wire n_18160;
wire n_14065;
wire n_8791;
wire n_11920;
wire n_10793;
wire n_8288;
wire n_17299;
wire n_14672;
wire n_14366;
wire n_15127;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_12786;
wire n_16022;
wire n_13382;
wire n_12711;
wire n_11675;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_17752;
wire n_9573;
wire n_15543;
wire n_5846;
wire n_8323;
wire n_10440;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_10391;
wire n_7636;
wire n_9799;
wire n_9695;
wire n_17235;
wire n_11306;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_7866;
wire n_11083;
wire n_13176;
wire n_15143;
wire n_9784;
wire n_11198;
wire n_18346;
wire n_7205;
wire n_18238;
wire n_18283;
wire n_8757;
wire n_7990;
wire n_7020;
wire n_13035;
wire n_10036;
wire n_18368;
wire n_13021;
wire n_17631;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_14905;
wire n_8596;
wire n_15128;
wire n_11840;
wire n_11698;
wire n_9556;
wire n_11292;
wire n_13157;
wire n_8590;
wire n_8720;
wire n_10261;
wire n_16682;
wire n_5708;
wire n_13502;
wire n_17038;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_5474;
wire n_14084;
wire n_15798;
wire n_12289;
wire n_16912;
wire n_10813;
wire n_10757;
wire n_13046;
wire n_5649;
wire n_11326;
wire n_6421;
wire n_13935;
wire n_11870;
wire n_16215;
wire n_7407;
wire n_9827;
wire n_14009;
wire n_16670;
wire n_13334;
wire n_10907;
wire n_5704;
wire n_15787;
wire n_11431;
wire n_7148;
wire n_14002;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_13646;
wire n_6236;
wire n_9417;
wire n_11834;
wire n_13361;
wire n_12020;
wire n_17286;
wire n_7214;
wire n_15061;
wire n_6007;
wire n_6144;
wire n_11506;
wire n_16205;
wire n_10135;
wire n_13161;
wire n_18186;
wire n_6197;
wire n_6658;
wire n_6835;
wire n_8834;
wire n_11624;
wire n_13399;
wire n_14010;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_15262;
wire n_16429;
wire n_16413;
wire n_5516;
wire n_7075;
wire n_6247;
wire n_10822;
wire n_11234;
wire n_14697;
wire n_15030;
wire n_10919;
wire n_18205;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_13967;
wire n_12099;
wire n_12858;
wire n_7467;
wire n_14609;
wire n_16451;
wire n_15351;
wire n_7799;
wire n_8364;
wire n_5698;
wire n_11092;
wire n_9534;
wire n_14310;
wire n_15228;
wire n_13380;
wire n_18170;
wire n_5771;
wire n_7544;
wire n_15832;
wire n_17369;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_11836;
wire n_17629;
wire n_6602;
wire n_17536;
wire n_10924;
wire n_15281;
wire n_15792;
wire n_17421;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_15675;
wire n_9647;
wire n_15515;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_16177;
wire n_10885;
wire n_15106;
wire n_6484;
wire n_13201;
wire n_18529;
wire n_6242;
wire n_12527;
wire n_14759;
wire n_13274;
wire n_12379;
wire n_9312;
wire n_9019;
wire n_13891;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_18222;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_12477;
wire n_7469;
wire n_5538;
wire n_14325;
wire n_15503;
wire n_14078;
wire n_17030;
wire n_7776;
wire n_10418;
wire n_14309;
wire n_10895;
wire n_10875;
wire n_11977;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_15576;
wire n_16256;
wire n_14222;
wire n_11696;
wire n_16741;
wire n_17416;
wire n_12400;
wire n_16990;
wire n_11734;
wire n_12114;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_11507;
wire n_16861;
wire n_14430;
wire n_9145;
wire n_15337;
wire n_17290;
wire n_13996;
wire n_17276;
wire n_7082;
wire n_12092;
wire n_14749;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_17944;
wire n_18483;
wire n_11837;
wire n_5428;
wire n_16545;
wire n_13709;
wire n_7451;
wire n_8260;
wire n_17713;
wire n_13898;
wire n_17679;
wire n_9000;
wire n_16507;
wire n_5677;
wire n_9454;
wire n_18442;
wire n_18505;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_16543;
wire n_18412;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_14704;
wire n_17003;
wire n_8307;
wire n_11967;
wire n_9383;
wire n_18096;
wire n_9253;
wire n_15084;
wire n_13559;
wire n_10571;
wire n_17692;
wire n_8874;
wire n_15258;
wire n_5927;
wire n_15071;
wire n_7495;
wire n_7392;
wire n_9566;
wire n_11338;
wire n_11996;
wire n_5435;
wire n_13426;
wire n_12174;
wire n_9765;
wire n_16322;
wire n_9807;
wire n_9057;
wire n_5200;
wire n_8706;
wire n_15220;
wire n_6400;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_16304;
wire n_6941;
wire n_12053;
wire n_15947;
wire n_17738;
wire n_5566;
wire n_12619;
wire n_11250;
wire n_7829;
wire n_18417;
wire n_7543;
wire n_13504;
wire n_16787;
wire n_15328;
wire n_8680;
wire n_11289;
wire n_13169;
wire n_7877;
wire n_7963;
wire n_13555;
wire n_9672;
wire n_12582;
wire n_16522;
wire n_5487;
wire n_15291;
wire n_8855;
wire n_18375;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_5486;
wire n_9503;
wire n_15345;
wire n_12423;
wire n_11391;
wire n_15462;
wire n_15426;
wire n_5244;
wire n_14721;
wire n_14137;
wire n_13265;
wire n_8270;
wire n_12714;
wire n_16051;
wire n_16779;
wire n_12153;
wire n_5889;
wire n_11738;
wire n_7284;
wire n_16905;
wire n_7264;
wire n_18196;
wire n_5391;
wire n_11522;
wire n_17765;
wire n_9763;
wire n_14163;
wire n_7737;
wire n_17851;
wire n_13666;
wire n_15523;
wire n_6537;
wire n_16569;
wire n_8614;
wire n_11070;
wire n_7328;
wire n_10702;
wire n_13337;
wire n_18459;
wire n_10958;
wire n_15682;
wire n_15112;
wire n_18146;
wire n_9479;
wire n_15556;
wire n_9162;
wire n_9568;
wire n_13730;
wire n_14849;
wire n_15621;
wire n_18411;
wire n_12405;
wire n_8816;
wire n_14041;
wire n_9119;
wire n_10319;
wire n_5849;
wire n_16661;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_10322;
wire n_7135;
wire n_13529;
wire n_6224;
wire n_8802;
wire n_6578;
wire n_9859;
wire n_14763;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_18293;
wire n_6092;
wire n_15912;
wire n_10879;
wire n_16206;
wire n_17686;
wire n_5951;
wire n_18381;
wire n_6241;
wire n_6589;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_18395;
wire n_10639;
wire n_16359;
wire n_17448;
wire n_16037;
wire n_16529;
wire n_8121;
wire n_8207;
wire n_12554;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_13351;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_17445;
wire n_7754;
wire n_15549;
wire n_10491;
wire n_12037;
wire n_15371;
wire n_17572;
wire n_13453;
wire n_15080;
wire n_5265;
wire n_16805;
wire n_12792;
wire n_15937;
wire n_11717;
wire n_9943;
wire n_16141;
wire n_5574;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_9821;
wire n_11112;
wire n_7152;
wire n_11723;
wire n_15246;
wire n_9575;
wire n_16647;
wire n_14940;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_18219;
wire n_11822;
wire n_18231;
wire n_10521;
wire n_9610;
wire n_15889;
wire n_12438;
wire n_11830;
wire n_15395;
wire n_5469;
wire n_14393;
wire n_8766;
wire n_12364;
wire n_12420;
wire n_12838;
wire n_16173;
wire n_9165;
wire n_6567;
wire n_16483;
wire n_16665;
wire n_13505;
wire n_14016;
wire n_12323;
wire n_5910;
wire n_15566;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_16231;
wire n_18461;
wire n_14369;
wire n_7240;
wire n_7570;
wire n_7033;
wire n_15354;
wire n_10476;
wire n_9966;
wire n_13156;
wire n_17805;
wire n_7817;
wire n_5682;
wire n_17318;
wire n_15529;
wire n_10710;
wire n_5387;
wire n_5557;
wire n_11394;
wire n_8850;
wire n_16794;
wire n_11906;
wire n_9928;
wire n_11820;
wire n_14647;
wire n_18384;
wire n_14298;
wire n_8002;
wire n_9741;
wire n_13897;
wire n_11486;
wire n_14792;
wire n_15280;
wire n_15999;
wire n_16290;
wire n_12677;
wire n_10180;
wire n_14248;
wire n_14112;
wire n_8370;
wire n_7237;
wire n_17867;
wire n_13300;
wire n_16296;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_16722;
wire n_9090;
wire n_16412;
wire n_16456;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_16364;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_9217;
wire n_9261;
wire n_17283;
wire n_9166;
wire n_12901;
wire n_17036;
wire n_10518;
wire n_8301;
wire n_12895;
wire n_17453;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_15170;
wire n_16936;
wire n_9771;
wire n_13401;
wire n_15774;
wire n_5316;
wire n_7718;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_13844;
wire n_14122;
wire n_16758;
wire n_7396;
wire n_10942;
wire n_12668;
wire n_12726;
wire n_17565;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_15437;
wire n_18543;
wire n_13010;
wire n_6320;
wire n_8126;
wire n_11239;
wire n_15819;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_12432;
wire n_10953;
wire n_7561;
wire n_15603;
wire n_18349;
wire n_6810;
wire n_7842;
wire n_12352;
wire n_17267;
wire n_17010;
wire n_9969;
wire n_6202;
wire n_10099;
wire n_11437;
wire n_12898;
wire n_9961;
wire n_14068;
wire n_16130;
wire n_17831;
wire n_12879;
wire n_14853;
wire n_16833;
wire n_5564;
wire n_11869;
wire n_13746;
wire n_14895;
wire n_12559;
wire n_13508;
wire n_5620;
wire n_14660;
wire n_15540;
wire n_7163;
wire n_16582;
wire n_10343;
wire n_18028;
wire n_10836;
wire n_15270;
wire n_17964;
wire n_9899;
wire n_9258;
wire n_16375;
wire n_13004;
wire n_10181;
wire n_15670;
wire n_18035;
wire n_10286;
wire n_5406;
wire n_13479;
wire n_8072;
wire n_10371;
wire n_14990;
wire n_16691;
wire n_8277;
wire n_7236;
wire n_16295;
wire n_18014;
wire n_13117;
wire n_10257;
wire n_7130;
wire n_5724;
wire n_14437;
wire n_7201;
wire n_11219;
wire n_10047;
wire n_14541;
wire n_16825;
wire n_13759;
wire n_16186;
wire n_10949;
wire n_5806;
wire n_13766;
wire n_10486;
wire n_11282;
wire n_11226;
wire n_16613;
wire n_8724;
wire n_5738;
wire n_18197;
wire n_15938;
wire n_17720;
wire n_17216;
wire n_16989;
wire n_11413;
wire n_14700;
wire n_15146;
wire n_5355;
wire n_16617;
wire n_5320;
wire n_16382;
wire n_7491;
wire n_13969;
wire n_5353;
wire n_9995;
wire n_13710;
wire n_16548;
wire n_5710;
wire n_5186;
wire n_9076;
wire n_11232;
wire n_12351;
wire n_18474;
wire n_12693;
wire n_9105;
wire n_6792;
wire n_16360;
wire n_12080;
wire n_16261;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_13359;
wire n_9668;
wire n_10372;
wire n_14867;
wire n_7559;
wire n_5438;
wire n_8867;
wire n_6044;
wire n_9491;
wire n_13259;
wire n_13335;
wire n_14022;
wire n_12702;
wire n_17811;
wire n_15188;
wire n_5517;
wire n_13175;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_14954;
wire n_10744;
wire n_12648;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_6125;
wire n_7314;
wire n_9095;
wire n_7678;
wire n_11334;
wire n_5907;
wire n_15757;
wire n_15979;
wire n_18465;
wire n_6045;
wire n_13075;
wire n_13129;
wire n_13736;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_14186;
wire n_7526;
wire n_14023;
wire n_17816;
wire n_17890;
wire n_6063;
wire n_16118;
wire n_10736;
wire n_10917;
wire n_16050;
wire n_6504;
wire n_11575;
wire n_18006;
wire n_7004;
wire n_7821;
wire n_14418;
wire n_12407;
wire n_13586;
wire n_8308;
wire n_6154;
wire n_15813;
wire n_11284;
wire n_6943;
wire n_10597;
wire n_14668;
wire n_16281;
wire n_17382;
wire n_11827;
wire n_13049;
wire n_8165;
wire n_13961;
wire n_14283;
wire n_12038;
wire n_17413;
wire n_14776;
wire n_8400;
wire n_10458;
wire n_15745;
wire n_8210;
wire n_11656;
wire n_12644;
wire n_18177;
wire n_5977;
wire n_10446;
wire n_13134;
wire n_11826;
wire n_7879;
wire n_18241;
wire n_10271;
wire n_16372;
wire n_10888;
wire n_15958;
wire n_10116;
wire n_15415;
wire n_16764;
wire n_14808;
wire n_7696;
wire n_18135;
wire n_11570;
wire n_16567;
wire n_6003;
wire n_12952;
wire n_16808;
wire n_6684;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_14795;
wire n_5451;
wire n_9323;
wire n_14140;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_9331;
wire n_6031;
wire n_9922;
wire n_10170;
wire n_13252;
wire n_11909;
wire n_8331;
wire n_12024;
wire n_13084;
wire n_14479;
wire n_16425;
wire n_16769;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_12004;
wire n_16622;
wire n_15374;
wire n_12830;
wire n_12637;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_7929;
wire n_10255;
wire n_16440;
wire n_16821;
wire n_18109;
wire n_10572;
wire n_14172;
wire n_16431;
wire n_12009;
wire n_13612;
wire n_7270;
wire n_13985;
wire n_11490;
wire n_17594;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_14124;
wire n_10113;
wire n_7550;
wire n_17498;
wire n_15077;
wire n_15086;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_6853;
wire n_6742;
wire n_10188;
wire n_13525;
wire n_17658;
wire n_18117;
wire n_5864;
wire n_10686;
wire n_15733;
wire n_15864;
wire n_9841;
wire n_14997;
wire n_15931;
wire n_13552;
wire n_6691;
wire n_8743;
wire n_18086;
wire n_7087;
wire n_12681;
wire n_14207;
wire n_8753;
wire n_14799;
wire n_6191;
wire n_16838;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_12634;
wire n_18419;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_13863;
wire n_8627;
wire n_17047;
wire n_18583;
wire n_14305;
wire n_9513;
wire n_16447;
wire n_14774;
wire n_9863;
wire n_12680;
wire n_15330;
wire n_11613;
wire n_13659;
wire n_16124;
wire n_10233;
wire n_12034;
wire n_10500;
wire n_16586;
wire n_15446;
wire n_10555;
wire n_5432;
wire n_15261;
wire n_15492;
wire n_18443;
wire n_10314;
wire n_6988;
wire n_17343;
wire n_11929;
wire n_10810;
wire n_11075;
wire n_16056;
wire n_7851;
wire n_6894;
wire n_13303;
wire n_13346;
wire n_12176;
wire n_9791;
wire n_13702;
wire n_16605;
wire n_10311;
wire n_9179;
wire n_15894;
wire n_5453;
wire n_13656;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_18237;
wire n_18533;
wire n_11177;
wire n_13667;
wire n_18056;
wire n_6817;
wire n_5842;
wire n_10937;
wire n_18367;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_12449;
wire n_5814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_16841;
wire n_10857;
wire n_15470;
wire n_18491;
wire n_11310;
wire n_13275;
wire n_12094;
wire n_6215;
wire n_16399;
wire n_11165;
wire n_9736;
wire n_5699;
wire n_5531;
wire n_14411;
wire n_5765;
wire n_12823;
wire n_15412;
wire n_12517;
wire n_6517;
wire n_15754;
wire n_6284;
wire n_18431;
wire n_5943;
wire n_15441;
wire n_17375;
wire n_10167;
wire n_7862;
wire n_16708;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_17353;
wire n_11923;
wire n_12071;
wire n_17439;
wire n_13832;
wire n_10630;
wire n_8105;
wire n_9031;
wire n_6088;
wire n_5777;
wire n_17955;
wire n_18113;
wire n_6883;
wire n_8808;
wire n_10061;
wire n_15257;
wire n_12963;
wire n_10428;
wire n_16860;
wire n_17869;
wire n_13087;
wire n_13972;
wire n_15599;
wire n_11865;
wire n_15436;
wire n_17920;
wire n_12366;
wire n_15633;
wire n_8528;
wire n_8204;
wire n_13024;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_14951;
wire n_5495;
wire n_10694;
wire n_15646;
wire n_12339;
wire n_10602;
wire n_18214;
wire n_16630;
wire n_7100;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_11041;
wire n_14632;
wire n_9420;
wire n_14490;
wire n_16995;
wire n_18347;
wire n_5655;
wire n_6393;
wire n_15969;
wire n_9708;
wire n_14336;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_14738;
wire n_15479;
wire n_7119;
wire n_8154;
wire n_7212;
wire n_5610;
wire n_6966;
wire n_8889;
wire n_13986;
wire n_9790;
wire n_13849;
wire n_13796;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_15522;
wire n_17577;
wire n_5759;
wire n_10778;
wire n_17874;
wire n_17961;
wire n_6722;
wire n_17892;
wire n_13258;
wire n_7874;
wire n_6035;
wire n_13329;
wire n_8490;
wire n_7622;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_13166;
wire n_15435;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_13946;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_14464;
wire n_6364;
wire n_15028;
wire n_16754;
wire n_8635;
wire n_7420;
wire n_7102;
wire n_15482;
wire n_12605;
wire n_13618;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_16217;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_15535;
wire n_18132;
wire n_16633;
wire n_7831;
wire n_6253;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_8532;
wire n_17534;
wire n_14993;
wire n_14327;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_14097;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_11140;
wire n_16323;
wire n_5377;
wire n_17882;
wire n_6201;
wire n_8796;
wire n_12218;
wire n_5737;
wire n_12343;
wire n_17829;
wire n_10733;
wire n_17677;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_17014;
wire n_12597;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_13744;
wire n_11478;
wire n_12834;
wire n_16067;
wire n_18226;
wire n_15650;
wire n_10066;
wire n_13017;
wire n_17239;
wire n_12236;
wire n_14335;
wire n_12902;
wire n_6419;
wire n_8372;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_16230;
wire n_17042;
wire n_10088;
wire n_16884;
wire n_14887;
wire n_13038;
wire n_7225;
wire n_15199;
wire n_15087;
wire n_18153;
wire n_8077;
wire n_12892;
wire n_17768;
wire n_11294;
wire n_15667;
wire n_18530;
wire n_6244;
wire n_9812;
wire n_6900;
wire n_9337;
wire n_15419;
wire n_15219;
wire n_6755;
wire n_16948;
wire n_7361;
wire n_9432;
wire n_6565;
wire n_9949;
wire n_10289;
wire n_17295;
wire n_6942;
wire n_7705;
wire n_11819;
wire n_14889;
wire n_7228;
wire n_13762;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_7932;
wire n_11573;
wire n_9576;
wire n_13420;
wire n_7509;
wire n_10145;
wire n_5872;
wire n_6862;
wire n_14225;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_17200;
wire n_15053;
wire n_6255;
wire n_6840;
wire n_13005;
wire n_14805;
wire n_6338;
wire n_15267;
wire n_17675;
wire n_15009;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_7981;
wire n_6037;
wire n_9577;
wire n_9874;
wire n_12588;
wire n_17203;
wire n_15648;
wire n_12589;
wire n_17548;
wire n_5874;
wire n_6266;
wire n_14796;
wire n_14143;
wire n_6488;
wire n_8337;
wire n_7164;
wire n_9231;
wire n_11844;
wire n_15390;
wire n_14044;
wire n_17431;
wire n_17792;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_11364;
wire n_9569;
wire n_13184;
wire n_14823;
wire n_15634;
wire n_18249;
wire n_12790;
wire n_18561;
wire n_8632;
wire n_18134;
wire n_14691;
wire n_17000;
wire n_13535;
wire n_14982;
wire n_17397;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_16508;
wire n_16908;
wire n_8358;
wire n_10009;
wire n_14770;
wire n_9552;
wire n_12927;
wire n_11100;
wire n_13822;
wire n_9279;
wire n_14948;
wire n_11902;
wire n_16588;
wire n_6317;
wire n_8199;
wire n_16782;
wire n_5588;
wire n_11993;
wire n_17456;
wire n_10443;
wire n_17317;
wire n_8656;
wire n_7167;
wire n_10756;
wire n_12813;
wire n_14909;
wire n_6480;
wire n_15105;
wire n_17099;
wire n_14387;
wire n_10918;
wire n_13122;
wire n_13534;
wire n_16572;
wire n_11797;
wire n_18383;
wire n_12765;
wire n_14106;
wire n_7865;
wire n_15553;
wire n_13616;
wire n_15690;
wire n_12663;
wire n_10384;
wire n_9289;
wire n_11315;
wire n_16349;
wire n_17165;
wire n_5736;
wire n_15841;
wire n_17623;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_18083;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_7134;
wire n_9633;
wire n_15468;
wire n_17422;
wire n_11153;
wire n_12312;
wire n_17128;
wire n_10074;
wire n_9547;
wire n_13097;
wire n_6875;
wire n_13627;
wire n_17850;
wire n_10934;
wire n_10197;
wire n_15786;
wire n_16350;
wire n_8346;
wire n_8761;
wire n_13112;
wire n_15458;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_13734;
wire n_8226;
wire n_11949;
wire n_17532;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_16581;
wire n_9084;
wire n_18597;
wire n_5928;
wire n_12256;
wire n_5478;
wire n_6016;
wire n_11746;
wire n_11812;
wire n_9371;
wire n_14051;
wire n_13163;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_16968;
wire n_14650;
wire n_16837;
wire n_7267;
wire n_10367;
wire n_14610;
wire n_18068;
wire n_17680;
wire n_12315;
wire n_11505;
wire n_18551;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_14100;
wire n_17938;
wire n_12556;
wire n_12375;
wire n_12998;
wire n_7812;
wire n_7103;
wire n_13723;
wire n_13143;
wire n_9080;
wire n_14601;
wire n_14549;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_9519;
wire n_14717;
wire n_14814;
wire n_6367;
wire n_11363;
wire n_12156;
wire n_13564;
wire n_15794;
wire n_14459;
wire n_16426;
wire n_13128;
wire n_13490;
wire n_11530;
wire n_17663;
wire n_12671;
wire n_17066;
wire n_10621;
wire n_14913;
wire n_13411;
wire n_7056;
wire n_14645;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_13260;
wire n_17302;
wire n_10085;
wire n_7813;
wire n_15382;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_16031;
wire n_17823;
wire n_6080;
wire n_8182;
wire n_8387;
wire n_12525;
wire n_16116;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_12076;
wire n_14090;
wire n_15825;
wire n_6717;
wire n_6056;
wire n_15823;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_13758;
wire n_7200;
wire n_11359;
wire n_7688;
wire n_15997;
wire n_16820;
wire n_8707;
wire n_12357;
wire n_15424;
wire n_10561;
wire n_17301;
wire n_11434;
wire n_9208;
wire n_11791;
wire n_14695;
wire n_15554;
wire n_7611;
wire n_15836;
wire n_6873;
wire n_15966;
wire n_16251;
wire n_16009;
wire n_15309;
wire n_13212;
wire n_14463;
wire n_8494;
wire n_16978;
wire n_15166;
wire n_17218;
wire n_5812;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_15216;
wire n_8544;
wire n_18304;
wire n_11848;
wire n_13503;
wire n_11152;
wire n_15138;
wire n_10749;
wire n_16516;
wire n_16318;
wire n_18517;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_14166;
wire n_12180;
wire n_8788;
wire n_15608;
wire n_17533;
wire n_14405;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_14081;
wire n_7723;
wire n_11621;
wire n_10560;
wire n_10160;
wire n_9327;
wire n_7404;
wire n_16175;
wire n_12857;
wire n_13171;
wire n_5368;
wire n_8177;
wire n_9854;
wire n_14271;
wire n_16171;
wire n_7059;
wire n_7450;
wire n_11667;
wire n_12025;
wire n_14854;
wire n_8962;
wire n_17311;
wire n_9538;
wire n_14254;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_16137;
wire n_12208;
wire n_6145;
wire n_11964;
wire n_17455;
wire n_6539;
wire n_6926;
wire n_15266;
wire n_13421;
wire n_7271;
wire n_7826;
wire n_9713;
wire n_14565;
wire n_17248;
wire n_11298;
wire n_15796;
wire n_5933;
wire n_13495;
wire n_16501;
wire n_8993;
wire n_6204;
wire n_7076;
wire n_13474;
wire n_10300;
wire n_13949;
wire n_13314;
wire n_9588;
wire n_11403;
wire n_14903;
wire n_14218;
wire n_11741;
wire n_15107;
wire n_12383;
wire n_11912;
wire n_15537;
wire n_6842;
wire n_12773;
wire n_14967;
wire n_6866;
wire n_13876;
wire n_17108;
wire n_9044;
wire n_9423;
wire n_16619;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_18174;
wire n_14487;
wire n_14883;
wire n_12962;
wire n_17024;
wire n_6451;
wire n_9813;
wire n_9127;
wire n_14596;
wire n_6514;
wire n_16263;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_18482;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_16767;
wire n_12612;
wire n_9244;
wire n_16387;
wire n_17322;
wire n_9869;
wire n_11142;
wire n_16369;
wire n_15304;
wire n_7049;
wire n_5903;
wire n_14449;
wire n_17094;
wire n_17213;
wire n_17434;
wire n_15271;
wire n_5986;
wire n_16795;
wire n_17509;
wire n_6710;
wire n_8278;
wire n_12885;
wire n_14865;
wire n_11644;
wire n_15539;
wire n_6345;
wire n_16165;
wire n_9715;
wire n_15893;
wire n_17112;
wire n_8618;
wire n_18326;
wire n_12108;
wire n_9094;
wire n_17664;
wire n_15432;
wire n_13108;
wire n_5782;
wire n_7535;
wire n_13170;
wire n_10862;
wire n_11531;
wire n_8911;
wire n_8248;
wire n_9056;
wire n_11357;
wire n_14471;
wire n_9407;
wire n_11476;
wire n_15906;
wire n_14476;
wire n_13633;
wire n_9985;
wire n_15244;
wire n_12089;
wire n_12496;
wire n_14538;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_17999;
wire n_17888;
wire n_11959;
wire n_11367;
wire n_15478;
wire n_6957;
wire n_9361;
wire n_15943;
wire n_16797;
wire n_11921;
wire n_8495;
wire n_14532;
wire n_12676;
wire n_13976;
wire n_16578;
wire n_8783;
wire n_12987;
wire n_13579;
wire n_14557;
wire n_11566;
wire n_17452;
wire n_16650;
wire n_13913;
wire n_8529;
wire n_8733;
wire n_14639;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_17067;
wire n_15392;
wire n_10254;
wire n_14340;
wire n_18444;
wire n_14032;
wire n_14715;
wire n_7944;
wire n_15970;
wire n_16944;
wire n_13080;
wire n_11208;
wire n_15702;
wire n_18049;
wire n_7262;
wire n_11374;
wire n_8647;
wire n_12967;
wire n_13403;
wire n_12452;
wire n_15978;
wire n_15857;
wire n_14899;
wire n_15961;
wire n_8574;
wire n_17444;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_13557;
wire n_12232;
wire n_18115;
wire n_14952;
wire n_11859;
wire n_12818;
wire n_15616;
wire n_15773;
wire n_10386;
wire n_16709;
wire n_12128;
wire n_6379;
wire n_14060;
wire n_15589;
wire n_17491;
wire n_14018;
wire n_17757;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_15959;
wire n_5563;
wire n_15307;
wire n_13583;
wire n_11026;
wire n_14111;
wire n_8044;
wire n_13309;
wire n_16330;
wire n_5840;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9439;
wire n_9553;
wire n_11633;
wire n_15292;
wire n_11467;
wire n_17333;
wire n_15239;
wire n_7506;
wire n_12672;
wire n_17749;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_14361;
wire n_8330;
wire n_12760;
wire n_16658;
wire n_18291;
wire n_15444;
wire n_13455;
wire n_15560;
wire n_15065;
wire n_6232;
wire n_15289;
wire n_9132;
wire n_13172;
wire n_5717;
wire n_16234;
wire n_6017;
wire n_9696;
wire n_14943;
wire n_10861;
wire n_17035;
wire n_9120;
wire n_17335;
wire n_8879;
wire n_15771;
wire n_15508;
wire n_17610;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_12168;
wire n_6362;
wire n_17990;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_14148;
wire n_16496;
wire n_17097;
wire n_8903;
wire n_16765;
wire n_11030;
wire n_12590;
wire n_15605;
wire n_5871;
wire n_12924;
wire n_16331;
wire n_7142;
wire n_12577;
wire n_17711;
wire n_10182;
wire n_12732;
wire n_16813;
wire n_13928;
wire n_17171;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_17458;
wire n_16057;
wire n_7125;
wire n_16401;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_10073;
wire n_14619;
wire n_11655;
wire n_15781;
wire n_11017;
wire n_12843;
wire n_14448;
wire n_7241;
wire n_7247;
wire n_14279;
wire n_12069;
wire n_10419;
wire n_7172;
wire n_15656;
wire n_16899;
wire n_18455;
wire n_16957;
wire n_15427;
wire n_17364;
wire n_14622;
wire n_10333;
wire n_12430;
wire n_10317;
wire n_17856;
wire n_7893;
wire n_6213;
wire n_14739;
wire n_16649;
wire n_18330;
wire n_15687;
wire n_7235;
wire n_8540;
wire n_11248;
wire n_12613;
wire n_6239;
wire n_12270;
wire n_14365;
wire n_9915;
wire n_9325;
wire n_16021;
wire n_9196;
wire n_16448;
wire n_13407;
wire n_5896;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_17173;
wire n_13676;
wire n_18480;
wire n_9384;
wire n_18391;
wire n_16694;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_13788;
wire n_14555;
wire n_11141;
wire n_12695;
wire n_15467;
wire n_10893;
wire n_11093;
wire n_16537;
wire n_14219;
wire n_9251;
wire n_18227;
wire n_11576;
wire n_8939;
wire n_13584;
wire n_17716;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_15471;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_8468;
wire n_15968;
wire n_9665;
wire n_13181;
wire n_10201;
wire n_17893;
wire n_7096;
wire n_18303;
wire n_12210;
wire n_13327;
wire n_8778;
wire n_11197;
wire n_16487;
wire n_17592;
wire n_7442;
wire n_15047;
wire n_10093;
wire n_15428;
wire n_5567;
wire n_8343;
wire n_15014;
wire n_6174;
wire n_12006;
wire n_17106;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_14168;
wire n_6087;
wire n_7593;
wire n_17156;
wire n_17908;
wire n_16311;
wire n_12246;
wire n_18319;
wire n_5249;
wire n_14085;
wire n_18220;
wire n_8068;
wire n_15342;
wire n_9955;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_17402;
wire n_10107;
wire n_13975;
wire n_5969;
wire n_10196;
wire n_10121;
wire n_8198;
wire n_14573;
wire n_17433;
wire n_17884;
wire n_13085;
wire n_15536;
wire n_7780;
wire n_6828;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_13224;
wire n_11469;
wire n_6454;
wire n_12625;
wire n_9270;
wire n_14046;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_14142;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_14512;
wire n_8557;
wire n_6918;
wire n_6041;
wire n_9099;
wire n_12389;
wire n_16214;
wire n_13761;
wire n_9309;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_10814;
wire n_5276;
wire n_16034;
wire n_9627;
wire n_16219;
wire n_13971;
wire n_17008;
wire n_11252;
wire n_17017;
wire n_16563;
wire n_16750;
wire n_8012;
wire n_14456;
wire n_13364;
wire n_7672;
wire n_11494;
wire n_6664;
wire n_14743;
wire n_17055;
wire n_7318;
wire n_17575;
wire n_6472;
wire n_10218;
wire n_18067;
wire n_8114;
wire n_18492;
wire n_13131;
wire n_14941;
wire n_12995;
wire n_18261;
wire n_14406;
wire n_13209;
wire n_11154;
wire n_11700;
wire n_14859;
wire n_16227;
wire n_5879;
wire n_14563;
wire n_8062;
wire n_11883;
wire n_5238;
wire n_16329;
wire n_11256;
wire n_11832;
wire n_14959;
wire n_6166;
wire n_5855;
wire n_12370;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_15387;
wire n_16128;
wire n_16278;
wire n_10975;
wire n_11901;
wire n_17404;
wire n_6352;
wire n_12974;
wire n_9460;
wire n_15973;
wire n_17698;
wire n_8542;
wire n_10859;
wire n_13078;
wire n_18446;
wire n_7063;
wire n_7047;
wire n_11652;
wire n_14768;
wire n_14320;
wire n_6632;
wire n_11056;
wire n_17241;
wire n_8576;
wire n_14807;
wire n_13885;
wire n_6238;
wire n_15795;
wire n_10542;
wire n_16814;
wire n_8038;
wire n_13631;
wire n_13932;
wire n_16804;
wire n_18103;
wire n_15162;
wire n_10681;
wire n_15606;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_16494;
wire n_11572;
wire n_13370;
wire n_11894;
wire n_16746;
wire n_15929;
wire n_14493;
wire n_10222;
wire n_6724;
wire n_18306;
wire n_13113;
wire n_13387;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_8716;
wire n_11336;
wire n_6705;
wire n_15866;
wire n_17988;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_17410;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_14764;
wire n_7074;
wire n_8734;
wire n_9204;
wire n_9476;
wire n_11849;
wire n_9689;
wire n_12142;
wire n_16807;
wire n_15237;
wire n_16711;
wire n_15862;
wire n_10659;
wire n_6591;
wire n_7585;
wire n_12564;
wire n_5268;
wire n_13643;
wire n_9780;
wire n_6946;
wire n_18538;
wire n_6002;
wire n_17576;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_13607;
wire n_12983;
wire n_15538;
wire n_7037;
wire n_6289;
wire n_13697;
wire n_11784;
wire n_6424;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_14244;
wire n_17578;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_16271;
wire n_15541;
wire n_8768;
wire n_10884;
wire n_12886;
wire n_14114;
wire n_15870;
wire n_13980;
wire n_6532;
wire n_7293;
wire n_13000;
wire n_16366;
wire n_12035;
wire n_14362;
wire n_13006;
wire n_5640;
wire n_17807;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_14742;
wire n_15996;
wire n_6778;
wire n_14904;
wire n_17359;
wire n_6721;
wire n_5560;
wire n_13205;
wire n_6644;
wire n_6512;
wire n_17878;
wire n_5544;
wire n_12810;
wire n_8258;
wire n_6108;
wire n_10370;
wire n_16930;
wire n_18537;
wire n_9597;
wire n_13820;
wire n_13947;
wire n_11322;
wire n_5744;
wire n_6703;
wire n_12122;
wire n_11892;
wire n_17562;
wire n_5384;
wire n_15283;
wire n_13428;
wire n_5841;
wire n_12241;
wire n_12396;
wire n_15407;
wire n_7614;
wire n_9343;
wire n_15731;
wire n_15895;
wire n_16554;
wire n_17194;
wire n_7839;
wire n_17779;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_6086;
wire n_9837;
wire n_11421;
wire n_11057;
wire n_16668;
wire n_10969;
wire n_10896;
wire n_14474;
wire n_11966;
wire n_17450;
wire n_17761;
wire n_18011;
wire n_18139;
wire n_12748;
wire n_7383;
wire n_6805;
wire n_8863;
wire n_10562;
wire n_16829;
wire n_16042;
wire n_5941;
wire n_18501;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_14417;
wire n_5611;
wire n_6340;
wire n_10054;
wire n_10355;
wire n_11551;
wire n_6219;
wire n_7479;
wire n_6706;
wire n_12571;
wire n_16893;
wire n_11853;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_10598;
wire n_13034;
wire n_16770;
wire n_8947;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_15494;
wire n_17305;
wire n_18047;
wire n_18579;
wire n_7078;
wire n_8188;
wire n_13831;
wire n_16828;
wire n_6761;
wire n_8972;
wire n_10007;
wire n_11751;
wire n_16792;
wire n_18572;
wire n_17550;
wire n_11725;
wire n_11423;
wire n_5701;
wire n_13635;
wire n_6067;
wire n_10801;
wire n_18378;
wire n_9206;
wire n_12674;
wire n_17727;
wire n_17839;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_17185;
wire n_18488;
wire n_15698;
wire n_9567;
wire n_14637;
wire n_6811;
wire n_9061;
wire n_11495;
wire n_16865;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_17122;
wire n_17015;
wire n_7372;
wire n_17154;
wire n_16922;
wire n_5367;
wire n_16778;
wire n_12220;
wire n_17980;
wire n_6868;
wire n_8664;
wire n_16822;
wire n_10704;
wire n_17535;
wire n_11520;
wire n_11622;
wire n_16552;
wire n_5970;
wire n_16867;
wire n_16133;
wire n_12169;
wire n_16788;
wire n_12283;
wire n_12336;
wire n_16638;
wire n_7174;
wire n_14783;
wire n_13268;
wire n_18345;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_16338;
wire n_13383;
wire n_10457;
wire n_12543;
wire n_15088;
wire n_16129;
wire n_17079;
wire n_17976;
wire n_16383;
wire n_8021;
wire n_17968;
wire n_9705;
wire n_16585;
wire n_17538;
wire n_7803;
wire n_15124;
wire n_17490;
wire n_11012;
wire n_6111;
wire n_14158;
wire n_12595;
wire n_9624;
wire n_17836;
wire n_9701;
wire n_11502;
wire n_14236;
wire n_15348;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_10389;
wire n_11631;
wire n_16745;
wire n_13588;
wire n_13510;
wire n_13570;
wire n_14640;
wire n_6659;
wire n_15688;
wire n_9709;
wire n_13677;
wire n_13983;
wire n_6011;
wire n_9295;
wire n_9416;
wire n_14036;
wire n_13757;
wire n_6225;
wire n_11842;
wire n_14710;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_5502;
wire n_6218;
wire n_8982;
wire n_17899;
wire n_17489;
wire n_16678;
wire n_9929;
wire n_13317;
wire n_10264;
wire n_5850;
wire n_12920;
wire n_13910;
wire n_15029;
wire n_9953;
wire n_13737;
wire n_7086;
wire n_16590;
wire n_18188;
wire n_6648;
wire n_14286;
wire n_15578;
wire n_16640;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_17640;
wire n_7226;
wire n_7927;
wire n_9013;
wire n_6182;
wire n_12717;
wire n_18373;
wire n_6520;
wire n_12660;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_17846;
wire n_5876;
wire n_9998;
wire n_18195;
wire n_11795;
wire n_5521;
wire n_9850;
wire n_17662;
wire n_6601;
wire n_10916;
wire n_16247;
wire n_12141;
wire n_8584;
wire n_17651;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_13196;
wire n_17113;
wire n_13520;
wire n_16748;
wire n_15363;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_10301;
wire n_17399;
wire n_17482;
wire n_14955;
wire n_8034;
wire n_13018;
wire n_7025;
wire n_9364;
wire n_15886;
wire n_8228;
wire n_18240;
wire n_15139;
wire n_8076;
wire n_17022;
wire n_6826;
wire n_15856;
wire n_16015;
wire n_15824;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_15642;
wire n_9836;
wire n_10929;
wire n_14357;
wire n_9107;
wire n_11279;
wire n_18370;
wire n_11724;
wire n_16393;
wire n_13044;
wire n_11789;
wire n_14152;
wire n_13228;
wire n_11525;
wire n_13862;
wire n_13518;
wire n_8100;
wire n_11999;
wire n_13446;
wire n_13086;
wire n_10837;
wire n_14869;
wire n_14008;
wire n_17069;
wire n_10554;
wire n_8014;
wire n_8994;
wire n_17827;
wire n_8091;
wire n_8413;
wire n_12746;
wire n_5837;
wire n_10149;
wire n_16162;
wire n_17155;
wire n_10970;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_5825;
wire n_14651;
wire n_16285;
wire n_5491;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_7982;
wire n_15791;
wire n_12190;
wire n_14927;
wire n_12787;
wire n_8804;
wire n_13881;
wire n_15484;
wire n_15152;
wire n_11383;
wire n_12799;
wire n_11847;
wire n_11976;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_17205;
wire n_9769;
wire n_5547;
wire n_15205;
wire n_15882;
wire n_13747;
wire n_8158;
wire n_12511;
wire n_17740;
wire n_11167;
wire n_12532;
wire n_6879;
wire n_17059;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_8433;
wire n_10102;
wire n_8931;
wire n_5596;
wire n_18481;
wire n_6074;
wire n_8213;
wire n_5983;
wire n_14472;
wire n_10534;
wire n_11825;
wire n_10932;
wire n_10619;
wire n_7684;
wire n_11049;
wire n_14354;
wire n_14974;
wire n_15532;
wire n_8451;
wire n_5604;
wire n_5411;
wire n_8334;
wire n_12743;
wire n_16523;
wire n_16083;
wire n_17263;
wire n_8731;
wire n_10589;
wire n_11681;
wire n_11611;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_16113;
wire n_11202;
wire n_16848;
wire n_15587;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_10552;
wire n_10248;
wire n_5815;
wire n_7370;
wire n_9748;
wire n_13365;
wire n_15254;
wire n_7771;
wire n_6595;
wire n_15322;
wire n_18221;
wire n_13539;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_18324;
wire n_16287;
wire n_16169;
wire n_17917;
wire n_8539;
wire n_5695;
wire n_6027;
wire n_16289;
wire n_10205;
wire n_16947;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_14618;
wire n_16342;
wire n_17556;
wire n_15747;
wire n_17278;
wire n_9226;
wire n_5235;
wire n_10110;
wire n_13899;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_16355;
wire n_11688;
wire n_6888;
wire n_7173;
wire n_7042;
wire n_12715;
wire n_12434;
wire n_11709;
wire n_14328;
wire n_12628;
wire n_8122;
wire n_6095;
wire n_13444;
wire n_16235;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_16504;
wire n_17095;
wire n_17915;
wire n_7592;
wire n_17049;
wire n_16540;
wire n_14209;
wire n_11331;
wire n_14429;
wire n_5311;
wire n_12979;
wire n_16774;
wire n_16436;
wire n_9528;
wire n_16901;
wire n_6590;
wire n_14348;
wire n_10638;
wire n_17923;
wire n_7583;
wire n_12201;
wire n_14086;
wire n_12499;
wire n_6559;
wire n_9112;
wire n_15799;
wire n_18582;
wire n_12448;
wire n_17195;
wire n_18243;
wire n_11876;
wire n_5797;
wire n_9235;
wire n_16570;
wire n_10610;
wire n_11187;
wire n_12761;
wire n_5572;
wire n_13852;
wire n_16455;
wire n_9333;
wire n_7151;
wire n_15004;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_8950;
wire n_17813;
wire n_14089;
wire n_10758;
wire n_16625;
wire n_13431;
wire n_10190;
wire n_16025;
wire n_5520;
wire n_15758;
wire n_11804;
wire n_14234;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_6287;
wire n_12809;
wire n_13614;
wire n_8347;
wire n_17703;
wire n_14552;
wire n_7353;
wire n_9330;
wire n_12538;
wire n_14208;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_9490;
wire n_15693;
wire n_12029;
wire n_18140;
wire n_11052;
wire n_9355;
wire n_15954;
wire n_9523;
wire n_14584;
wire n_17350;
wire n_15386;
wire n_14620;
wire n_5888;
wire n_5669;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_15349;
wire n_18598;
wire n_7571;
wire n_9582;
wire n_10060;
wire n_5884;
wire n_6671;
wire n_13470;
wire n_16249;
wire n_11009;
wire n_18192;
wire n_6812;
wire n_12361;
wire n_9288;
wire n_9686;
wire n_16435;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_13068;
wire n_6308;
wire n_16723;
wire n_7897;
wire n_17130;
wire n_11446;
wire n_10910;
wire n_17701;
wire n_10162;
wire n_18552;
wire n_8242;
wire n_7118;
wire n_15002;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_13248;
wire n_7792;
wire n_15985;
wire n_17296;
wire n_17515;
wire n_13842;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_15338;
wire n_15378;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_14501;
wire n_17881;
wire n_6738;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_8703;
wire n_10014;
wire n_15723;
wire n_7109;
wire n_12642;
wire n_15839;
wire n_16840;
wire n_12484;
wire n_16135;
wire n_6128;
wire n_13549;
wire n_8822;
wire n_6029;
wire n_14790;
wire n_17361;
wire n_14999;
wire n_17661;
wire n_10677;
wire n_17204;
wire n_12187;
wire n_18269;
wire n_5751;
wire n_15852;
wire n_5264;
wire n_16080;
wire n_12321;
wire n_5924;
wire n_9992;
wire n_11247;
wire n_15180;
wire n_15692;
wire n_18581;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_12669;
wire n_13106;
wire n_18079;
wire n_17201;
wire n_8476;
wire n_14296;
wire n_14294;
wire n_6702;
wire n_11927;
wire n_17745;
wire n_16674;
wire n_17609;
wire n_13720;
wire n_11179;
wire n_16326;
wire n_6701;
wire n_16571;
wire n_17074;
wire n_7339;
wire n_14862;
wire n_13706;
wire n_8359;
wire n_7380;
wire n_13903;
wire n_15808;
wire n_9051;
wire n_8736;
wire n_8545;
wire n_10385;
wire n_7749;
wire n_10078;
wire n_10105;
wire n_11514;
wire n_12470;
wire n_12994;
wire n_11321;
wire n_14313;
wire n_15785;
wire n_9500;
wire n_16752;
wire n_18496;
wire n_8705;
wire n_14574;
wire n_10215;
wire n_14451;
wire n_11779;
wire n_14059;
wire n_7508;
wire n_17114;
wire n_5694;
wire n_9455;
wire n_10251;
wire n_8708;
wire n_14211;
wire n_15234;
wire n_10834;
wire n_7574;
wire n_17632;
wire n_14092;
wire n_17611;
wire n_17524;
wire n_9980;
wire n_14509;
wire n_14394;
wire n_11882;
wire n_13516;
wire n_17649;
wire n_11647;
wire n_15027;
wire n_12064;
wire n_14273;
wire n_15404;
wire n_10706;
wire n_12462;
wire n_6005;
wire n_8872;
wire n_12696;
wire n_17261;
wire n_9555;
wire n_15735;
wire n_18024;
wire n_11133;
wire n_5449;
wire n_16462;
wire n_14845;
wire n_6169;
wire n_8238;
wire n_15230;
wire n_17143;
wire n_12735;
wire n_7713;
wire n_15465;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_16182;
wire n_10709;
wire n_12646;
wire n_10871;
wire n_15858;
wire n_15875;
wire n_18341;
wire n_7352;
wire n_16405;
wire n_5926;
wire n_10304;
wire n_5398;
wire n_5860;
wire n_6936;
wire n_14624;
wire n_10244;
wire n_15934;
wire n_16600;
wire n_15036;
wire n_16827;
wire n_17695;
wire n_18193;
wire n_14765;
wire n_16121;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_16170;
wire n_14120;
wire n_14995;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_13794;
wire n_7641;
wire n_17479;
wire n_18512;
wire n_6106;
wire n_7203;
wire n_12999;
wire n_13537;
wire n_14407;
wire n_14260;
wire n_9397;
wire n_16845;
wire n_17307;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_18258;
wire n_12682;
wire n_16010;
wire n_14802;
wire n_9673;
wire n_14434;
wire n_14175;
wire n_17574;
wire n_6848;
wire n_17415;
wire n_8642;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11941;
wire n_11875;
wire n_5919;
wire n_8159;
wire n_14834;
wire n_18567;
wire n_12111;
wire n_15780;
wire n_8912;
wire n_14346;
wire n_18085;
wire n_16955;
wire n_13463;
wire n_7439;
wire n_9496;
wire n_16241;
wire n_15189;
wire n_17653;
wire n_8110;
wire n_14275;
wire n_5319;
wire n_10796;
wire n_14506;
wire n_10016;
wire n_12903;
wire n_9008;
wire n_12079;
wire n_15335;
wire n_6343;
wire n_12593;
wire n_16018;
wire n_14615;
wire n_5270;
wire n_10030;
wire n_15227;
wire n_15222;
wire n_8805;
wire n_6850;
wire n_17922;
wire n_12864;
wire n_17849;
wire n_15285;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_13294;
wire n_15689;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_7209;
wire n_6014;
wire n_7112;
wire n_15026;
wire n_17474;
wire n_13895;
wire n_11307;
wire n_5181;
wire n_13936;
wire n_17860;
wire n_13933;
wire n_18274;
wire n_6979;
wire n_7815;
wire n_13222;
wire n_7934;
wire n_9545;
wire n_13813;
wire n_16190;
wire n_8111;
wire n_18315;
wire n_9629;
wire n_9603;
wire n_11578;
wire n_6865;
wire n_18003;
wire n_10432;
wire n_12719;
wire n_16888;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_18376;
wire n_15361;
wire n_18595;
wire n_8739;
wire n_17078;
wire n_6747;
wire n_9674;
wire n_13714;
wire n_16244;
wire n_17284;
wire n_5583;
wire n_13438;
wire n_6433;
wire n_17862;
wire n_15987;
wire n_10462;
wire n_18253;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_15850;
wire n_15469;
wire n_11769;
wire n_8856;
wire n_6142;
wire n_9930;
wire n_16079;
wire n_11908;
wire n_14371;
wire n_12925;
wire n_18166;
wire n_5775;
wire n_17140;
wire n_14901;
wire n_6462;
wire n_17372;
wire n_7769;
wire n_14988;
wire n_18407;
wire n_6034;
wire n_17034;
wire n_9781;
wire n_10291;
wire n_13159;
wire n_9659;
wire n_18575;
wire n_17502;
wire n_14333;
wire n_16293;
wire n_7233;
wire n_8732;
wire n_13636;
wire n_13506;
wire n_13287;
wire n_11913;
wire n_14788;
wire n_7602;
wire n_9296;
wire n_18587;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_14590;
wire n_11341;
wire n_7390;
wire n_10787;
wire n_13389;
wire n_10669;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_14603;
wire n_8231;
wire n_17726;
wire n_16308;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_13905;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_16986;
wire n_13717;
wire n_17872;
wire n_12317;
wire n_13302;
wire n_6071;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_15119;
wire n_15821;
wire n_8908;
wire n_10185;
wire n_11182;
wire n_10092;
wire n_16085;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_16766;
wire n_17834;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_12782;
wire n_15256;
wire n_11231;
wire n_14145;
wire n_18366;
wire n_8090;
wire n_13740;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_17966;
wire n_12875;
wire n_15982;
wire n_15064;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_17796;
wire n_13918;
wire n_8137;
wire n_7045;
wire n_13775;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_10983;
wire n_9987;
wire n_15218;
wire n_15452;
wire n_17366;
wire n_7984;
wire n_11727;
wire n_13615;
wire n_15625;
wire n_17514;
wire n_6788;
wire n_18307;
wire n_7014;
wire n_17975;
wire n_12633;
wire n_12192;
wire n_10430;
wire n_14779;
wire n_16697;
wire n_15114;
wire n_18110;
wire n_8305;
wire n_14973;
wire n_10277;
wire n_16751;
wire n_18147;
wire n_17934;
wire n_8163;
wire n_7220;
wire n_18015;
wire n_17342;
wire n_6709;
wire n_16632;
wire n_14465;
wire n_13412;
wire n_16028;
wire n_17525;
wire n_10948;
wire n_11749;
wire n_18242;
wire n_6712;
wire n_6550;
wire n_10525;
wire n_9507;
wire n_14287;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_15296;
wire n_15828;
wire n_18107;
wire n_8841;
wire n_14553;
wire n_16126;
wire n_13457;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_16594;
wire n_18102;
wire n_16370;
wire n_18066;
wire n_18545;
wire n_15136;
wire n_6743;
wire n_12497;
wire n_15043;
wire n_10354;
wire n_16223;
wire n_12412;
wire n_16168;
wire n_11880;
wire n_5785;
wire n_16602;
wire n_15915;
wire n_7465;
wire n_14528;
wire n_13177;
wire n_5967;
wire n_10049;
wire n_12724;
wire n_16864;
wire n_14958;
wire n_15551;
wire n_16761;
wire n_6672;
wire n_9457;
wire n_9485;
wire n_5780;
wire n_7679;
wire n_13940;
wire n_16738;
wire n_18133;
wire n_7936;
wire n_8966;
wire n_6084;
wire n_11249;
wire n_16744;
wire n_17876;
wire n_15449;
wire n_10287;
wire n_15992;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_14342;
wire n_12101;
wire n_10119;
wire n_13693;
wire n_11145;
wire n_12606;
wire n_17406;
wire n_11986;
wire n_16684;
wire n_8395;
wire n_10900;
wire n_14798;
wire n_5966;
wire n_10349;
wire n_6634;
wire n_14107;
wire n_14758;
wire n_18392;
wire n_5213;
wire n_8961;
wire n_14781;
wire n_17579;
wire n_10849;
wire n_7462;
wire n_13333;
wire n_16802;
wire n_13229;
wire n_5735;
wire n_12118;
wire n_17909;
wire n_18439;
wire n_17336;
wire n_13311;
wire n_14409;
wire n_14724;
wire n_16340;
wire n_18451;
wire n_7490;
wire n_11380;
wire n_15737;
wire n_14291;
wire n_7545;
wire n_10792;
wire n_15573;
wire n_11513;
wire n_8625;
wire n_13296;
wire n_16020;
wire n_7464;
wire n_7160;
wire n_9809;
wire n_8937;
wire n_6919;
wire n_14611;
wire n_10750;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_7295;
wire n_7115;
wire n_12087;
wire n_13675;
wire n_9192;
wire n_15022;
wire n_17863;
wire n_14338;
wire n_7348;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_17554;
wire n_6104;
wire n_16071;
wire n_8179;
wire n_10537;
wire n_17088;
wire n_11861;
wire n_15051;
wire n_6548;
wire n_15394;
wire n_6082;
wire n_6993;
wire n_8511;
wire n_15916;
wire n_6973;
wire n_16875;
wire n_12081;
wire n_18305;
wire n_15941;
wire n_10426;
wire n_9558;
wire n_11594;
wire n_7453;
wire n_16468;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_15639;
wire n_10684;
wire n_7162;
wire n_16655;
wire n_11436;
wire n_12346;
wire n_18095;
wire n_11729;
wire n_18167;
wire n_15039;
wire n_8371;
wire n_17929;
wire n_8702;
wire n_13916;
wire n_15195;
wire n_17158;
wire n_8116;
wire n_7946;
wire n_8195;
wire n_17027;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_14069;
wire n_17056;
wire n_12244;
wire n_18452;
wire n_17400;
wire n_5877;
wire n_9991;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_11366;
wire n_17438;
wire n_11872;
wire n_7681;
wire n_8845;
wire n_15198;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_13620;
wire n_16434;
wire n_5189;
wire n_17902;
wire n_13930;
wire n_7702;
wire n_6676;
wire n_13981;
wire n_8149;
wire n_16850;
wire n_10823;
wire n_9976;
wire n_8042;
wire n_11516;
wire n_17144;
wire n_14766;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_8392;
wire n_9560;
wire n_14659;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_14592;
wire n_10830;
wire n_15109;
wire n_18362;
wire n_11132;
wire n_16868;
wire n_17625;
wire n_6718;
wire n_18546;
wire n_18034;
wire n_15007;
wire n_17644;
wire n_18181;
wire n_7503;
wire n_17126;
wire n_10824;
wire n_6854;
wire n_17254;
wire n_15400;
wire n_17411;
wire n_15197;
wire n_16866;
wire n_16216;
wire n_15485;
wire n_18499;
wire n_14841;
wire n_16726;
wire n_13624;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_14277;
wire n_5425;
wire n_18603;
wire n_5886;
wire n_8269;
wire n_13493;
wire n_6032;
wire n_9047;
wire n_13805;
wire n_16389;
wire n_12953;
wire n_12842;
wire n_15224;
wire n_18569;
wire n_8968;
wire n_12481;
wire n_16243;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_18168;
wire n_5446;
wire n_11316;
wire n_7855;
wire n_14029;
wire n_11047;
wire n_14963;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_8399;
wire n_16916;
wire n_14648;
wire n_11767;
wire n_9599;
wire n_14056;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_13866;
wire n_9401;
wire n_5678;
wire n_13695;
wire n_12435;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_17463;
wire n_11586;
wire n_6981;
wire n_18106;
wire n_15817;
wire n_15344;
wire n_13288;
wire n_7065;
wire n_12149;
wire n_13669;
wire n_9216;
wire n_12002;
wire n_12836;
wire n_16917;
wire n_17179;
wire n_17245;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_17084;
wire n_13840;
wire n_11229;
wire n_13548;
wire n_15710;
wire n_16601;
wire n_16159;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_14251;
wire n_17570;
wire n_6122;
wire n_11397;
wire n_11225;
wire n_16240;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_17486;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_17504;
wire n_17190;
wire n_12840;
wire n_7330;
wire n_14605;
wire n_17973;
wire n_5437;
wire n_8883;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_11058;
wire n_9058;
wire n_15888;
wire n_7336;
wire n_11471;
wire n_14705;
wire n_7446;
wire n_13543;
wire n_18547;
wire n_17660;
wire n_8401;
wire n_16700;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_10577;
wire n_13772;
wire n_14679;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_15487;
wire n_7357;
wire n_17940;
wire n_8756;
wire n_11324;
wire n_17064;
wire n_8737;
wire n_18045;
wire n_13925;
wire n_10334;
wire n_13406;
wire n_12945;
wire n_16371;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_18334;
wire n_17385;
wire n_10151;
wire n_6439;
wire n_11614;
wire n_14040;
wire n_16704;
wire n_8602;
wire n_14054;
wire n_18223;
wire n_13368;
wire n_8240;
wire n_12850;
wire n_13469;
wire n_14507;
wire n_7714;
wire n_5407;
wire n_10411;
wire n_15242;
wire n_13249;
wire n_9484;
wire n_12984;
wire n_16193;
wire n_10989;
wire n_8422;
wire n_17725;
wire n_10939;
wire n_13587;
wire n_12224;
wire n_5913;
wire n_7088;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_17495;
wire n_8878;
wire n_11144;
wire n_11361;
wire n_10090;
wire n_7440;
wire n_6406;
wire n_14872;
wire n_6945;
wire n_8112;
wire n_14034;
wire n_17681;
wire n_11567;
wire n_10962;
wire n_7029;
wire n_17676;
wire n_14797;
wire n_11128;
wire n_9292;
wire n_9622;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_12197;
wire n_14177;
wire n_17753;
wire n_14093;
wire n_10186;
wire n_14607;
wire n_17236;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_6618;
wire n_13326;
wire n_15901;
wire n_6474;
wire n_13082;
wire n_14453;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_17545;
wire n_6226;
wire n_13094;
wire n_18518;
wire n_7317;
wire n_10856;
wire n_12403;
wire n_17919;
wire n_6000;
wire n_12679;
wire n_13481;
wire n_9584;
wire n_13692;
wire n_8194;
wire n_9461;
wire n_8055;
wire n_11168;
wire n_14921;
wire n_17558;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_8360;
wire n_12018;
wire n_18040;
wire n_6425;
wire n_17393;
wire n_14457;
wire n_5294;
wire n_6493;
wire n_16097;
wire n_16931;
wire n_9845;
wire n_16147;
wire n_7374;
wire n_6250;
wire n_6502;
wire n_6288;
wire n_5974;
wire n_14382;
wire n_14389;
wire n_11937;
wire n_12872;
wire n_18189;
wire n_13396;
wire n_7522;
wire n_17277;
wire n_6492;
wire n_10071;
wire n_14517;
wire n_8755;
wire n_6046;
wire n_11460;
wire n_8251;
wire n_13713;
wire n_5323;
wire n_11565;
wire n_14621;
wire n_12372;
wire n_9618;
wire n_14911;
wire n_6118;
wire n_13608;
wire n_5810;
wire n_15405;
wire n_7046;
wire n_17875;
wire n_11192;
wire n_11808;
wire n_17970;
wire n_15643;
wire n_13257;
wire n_10956;
wire n_6852;
wire n_15420;
wire n_17160;
wire n_8677;
wire n_13052;
wire n_18509;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_5991;
wire n_14934;
wire n_17206;
wire n_17636;
wire n_13914;
wire n_16634;
wire n_12572;
wire n_12453;
wire n_14663;
wire n_16762;
wire n_10035;
wire n_5702;
wire n_16921;
wire n_17559;
wire n_18094;
wire n_17870;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_14962;
wire n_15652;
wire n_13922;
wire n_9699;
wire n_17435;
wire n_13277;
wire n_12340;
wire n_13423;
wire n_8108;
wire n_18149;
wire n_16713;
wire n_14578;
wire n_18143;
wire n_15653;
wire n_5243;
wire n_5914;
wire n_16742;
wire n_12955;
wire n_17065;
wire n_12068;
wire n_10252;
wire n_18464;
wire n_5250;
wire n_16641;
wire n_11555;
wire n_13494;
wire n_6869;
wire n_17285;
wire n_10041;
wire n_9321;
wire n_15499;
wire n_14625;
wire n_5590;
wire n_16856;
wire n_10345;
wire n_14514;
wire n_18555;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_17612;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_5809;
wire n_14256;
wire n_15016;
wire n_16773;
wire n_10543;
wire n_7924;
wire n_17225;
wire n_18493;
wire n_12394;
wire n_13578;
wire n_7659;
wire n_9005;
wire n_9161;
wire n_14204;
wire n_16203;
wire n_8875;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_15855;
wire n_7153;
wire n_11101;
wire n_12954;
wire n_7836;
wire n_10737;
wire n_12662;
wire n_15697;
wire n_17879;
wire n_17910;
wire n_14082;
wire n_17750;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_7280;
wire n_10644;
wire n_12801;
wire n_13448;
wire n_14688;
wire n_15865;
wire n_16928;
wire n_5813;
wire n_18594;
wire n_9293;
wire n_12503;
wire n_13708;
wire n_10365;
wire n_13767;
wire n_5833;
wire n_11781;
wire n_11055;
wire n_18510;
wire n_7886;
wire n_15728;
wire n_16616;
wire n_14832;
wire n_15202;
wire n_18218;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_17599;
wire n_18292;
wire n_7012;
wire n_12965;
wire n_13029;
wire n_17354;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_14571;
wire n_18224;
wire n_16400;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_15707;
wire n_18297;
wire n_16328;
wire n_5816;
wire n_10809;
wire n_15396;
wire n_8927;
wire n_16934;
wire n_10899;
wire n_17985;
wire n_15347;
wire n_15909;
wire n_16396;
wire n_17531;
wire n_9639;
wire n_15155;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_15250;
wire n_17193;
wire n_6228;
wire n_6711;
wire n_11884;
wire n_11997;
wire n_5416;
wire n_8946;
wire n_16517;
wire n_14881;
wire n_18588;
wire n_13090;
wire n_14527;
wire n_12822;
wire n_13541;
wire n_13307;
wire n_13371;
wire n_11863;
wire n_16958;
wire n_17868;
wire n_7279;
wire n_7971;
wire n_13908;
wire n_9646;
wire n_17460;
wire n_8017;
wire n_17396;
wire n_12264;
wire n_13312;
wire n_17033;
wire n_11761;
wire n_17234;
wire n_8474;
wire n_9984;
wire n_16174;
wire n_7275;
wire n_8232;
wire n_18059;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_9649;
wire n_14703;
wire n_8904;
wire n_16977;
wire n_11199;
wire n_13533;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_16283;
wire n_17642;
wire n_10629;
wire n_18329;
wire n_9562;
wire n_7007;
wire n_7070;
wire n_8382;
wire n_13023;
wire n_16088;
wire n_7610;
wire n_6072;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_13856;
wire n_16229;
wire n_15607;
wire n_10006;
wire n_11757;
wire n_7259;
wire n_12320;
wire n_12274;
wire n_14588;
wire n_15879;
wire n_18447;
wire n_15315;
wire n_9759;
wire n_6353;
wire n_12622;
wire n_6992;
wire n_11185;
wire n_12659;
wire n_8128;
wire n_13440;
wire n_15226;
wire n_6818;
wire n_15746;
wire n_13436;
wire n_10206;
wire n_15921;
wire n_17736;
wire n_6322;
wire n_15425;
wire n_5661;
wire n_16878;
wire n_5932;
wire n_5830;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_16982;
wire n_12629;
wire n_7539;
wire n_12586;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_18294;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_11081;
wire n_8481;
wire n_10275;
wire n_7775;
wire n_13011;
wire n_16687;
wire n_11392;
wire n_9981;
wire n_18514;
wire n_14858;
wire n_7930;
wire n_17222;
wire n_5558;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_16513;
wire n_6378;
wire n_13911;
wire n_5383;
wire n_14495;
wire n_16498;
wire n_16879;
wire n_8205;
wire n_14165;
wire n_9907;
wire n_17544;
wire n_13088;
wire n_6976;
wire n_5587;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_12269;
wire n_13538;
wire n_7640;
wire n_14617;
wire n_17309;
wire n_13701;
wire n_9816;
wire n_13787;
wire n_10498;
wire n_11424;
wire n_13486;
wire n_12585;
wire n_14021;
wire n_13674;
wire n_14263;
wire n_11463;
wire n_17132;
wire n_13912;
wire n_18311;
wire n_14303;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_8605;
wire n_11278;
wire n_14445;
wire n_10358;
wire n_7548;
wire n_10635;
wire n_13626;
wire n_17541;
wire n_17593;
wire n_16732;
wire n_9944;
wire n_5954;
wire n_6156;
wire n_12832;
wire n_12913;
wire n_6998;
wire n_8067;
wire n_17394;
wire n_7587;
wire n_7064;
wire n_16158;
wire n_12301;
wire n_16839;
wire n_17496;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_16798;
wire n_17472;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_14427;
wire n_18402;
wire n_7197;
wire n_9676;
wire n_5645;
wire n_15822;
wire n_11881;
wire n_7393;
wire n_18327;
wire n_11332;
wire n_6917;
wire n_13629;
wire n_6937;
wire n_7591;
wire n_13207;
wire n_14980;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_7727;
wire n_18025;
wire n_7358;
wire n_17211;
wire n_16488;
wire n_15994;
wire n_7324;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_18088;
wire n_11935;
wire n_13589;
wire n_15730;
wire n_17568;
wire n_17561;
wire n_15685;
wire n_18089;
wire n_17967;
wire n_6301;
wire n_9788;
wire n_18061;
wire n_16815;
wire n_18022;
wire n_6929;
wire n_15570;
wire n_15562;
wire n_11309;
wire n_16273;
wire n_16706;
wire n_17207;
wire n_8719;
wire n_16140;
wire n_8045;
wire n_10785;
wire n_16032;
wire n_18262;
wire n_7729;
wire n_13872;
wire n_18046;
wire n_15493;
wire n_17646;
wire n_12341;
wire n_12615;
wire n_6436;
wire n_18389;
wire n_5412;
wire n_14475;
wire n_16987;
wire n_18337;
wire n_16959;
wire n_8209;
wire n_13357;
wire n_10802;
wire n_14477;
wire n_10815;
wire n_17148;
wire n_7565;
wire n_6699;
wire n_12926;
wire n_16624;
wire n_14809;
wire n_9213;
wire n_7291;
wire n_14725;
wire n_7631;
wire n_14522;
wire n_16971;
wire n_8784;
wire n_16892;
wire n_7382;
wire n_13869;
wire n_13955;
wire n_16903;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_17708;
wire n_9340;
wire n_16527;
wire n_13561;
wire n_12167;
wire n_14720;
wire n_9473;
wire n_14400;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_16725;
wire n_16904;
wire n_17963;
wire n_15019;
wire n_6677;
wire n_12161;
wire n_16432;
wire n_13499;
wire n_16873;
wire n_12085;
wire n_17107;
wire n_14843;
wire n_11735;
wire n_7618;
wire n_10647;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_16781;
wire n_18190;
wire n_6764;
wire n_8575;
wire n_13554;
wire n_12298;
wire n_10081;
wire n_18421;
wire n_5733;
wire n_10324;
wire n_11189;
wire n_6780;
wire n_12569;
wire n_8815;
wire n_11582;
wire n_14929;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_18497;
wire n_9303;
wire n_11105;
wire n_11705;
wire n_8261;
wire n_7673;
wire n_13698;
wire n_6830;
wire n_17391;
wire n_13894;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_17039;
wire n_17682;
wire n_7282;
wire n_6586;
wire n_9968;
wire n_10808;
wire n_11474;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_16819;
wire n_18504;
wire n_8086;
wire n_16612;
wire n_15466;
wire n_13595;
wire n_8789;
wire n_5946;
wire n_5997;
wire n_13943;
wire n_7953;
wire n_13540;
wire n_17124;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_14642;
wire n_9722;
wire n_13283;
wire n_12042;
wire n_12155;
wire n_14827;
wire n_5657;
wire n_15481;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_13465;
wire n_8695;
wire n_12373;
wire n_15615;
wire n_5975;
wire n_15664;
wire n_16149;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_17430;
wire n_14579;
wire n_17930;
wire n_8363;
wire n_15388;
wire n_17802;
wire n_10652;
wire n_10545;
wire n_9669;
wire n_17775;
wire n_17945;
wire n_8665;
wire n_13098;
wire n_13733;
wire n_16557;
wire n_8282;
wire n_6510;
wire n_15847;
wire n_9388;
wire n_5938;
wire n_15972;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_12654;
wire n_14141;
wire n_17446;
wire n_5602;
wire n_9379;
wire n_11992;
wire n_15790;
wire n_7751;
wire n_17061;
wire n_10869;
wire n_14880;
wire n_18573;
wire n_14718;
wire n_14975;
wire n_13142;
wire n_18298;
wire n_7581;
wire n_13180;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_17960;
wire n_17314;
wire n_15217;
wire n_14589;
wire n_17837;
wire n_5246;
wire n_10453;
wire n_12386;
wire n_14257;
wire n_13308;
wire n_9952;
wire n_16492;
wire n_16811;
wire n_16975;
wire n_16716;
wire n_15323;
wire n_9911;
wire n_12183;
wire n_5579;
wire n_8835;
wire n_16317;
wire n_15187;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_5750;
wire n_10688;
wire n_13785;
wire n_5831;
wire n_7742;
wire n_16771;
wire n_9274;
wire n_12964;
wire n_10473;
wire n_15712;
wire n_16404;
wire n_14007;
wire n_16985;
wire n_15099;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_10957;
wire n_13373;
wire n_7579;
wire n_13517;
wire n_17230;
wire n_12863;
wire n_16874;
wire n_10352;
wire n_11188;
wire n_7428;
wire n_5666;
wire n_12221;
wire n_9195;
wire n_10442;
wire n_16236;
wire n_11687;
wire n_17787;
wire n_16830;
wire n_8870;
wire n_13973;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_11774;
wire n_7283;
wire n_8507;
wire n_6475;
wire n_7015;
wire n_7699;
wire n_17530;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_13206;
wire n_9623;
wire n_6103;
wire n_15951;
wire n_5546;
wire n_7249;
wire n_10713;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_15939;
wire n_14102;
wire n_6680;
wire n_10954;
wire n_7985;
wire n_17196;
wire n_13637;
wire n_12267;
wire n_15803;
wire n_7432;
wire n_8365;
wire n_16036;
wire n_16705;
wire n_18163;
wire n_13978;
wire n_13941;
wire n_15339;
wire n_13439;
wire n_16702;
wire n_13780;
wire n_8893;
wire n_16699;
wire n_16152;
wire n_6372;
wire n_14133;
wire n_14433;
wire n_11329;
wire n_15904;
wire n_7194;
wire n_5994;
wire n_6495;
wire n_17280;
wire n_9516;
wire n_13241;
wire n_16027;
wire n_13187;
wire n_13162;
wire n_12768;
wire n_6752;
wire n_8976;
wire n_6426;
wire n_7505;
wire n_17844;
wire n_5626;
wire n_18136;
wire n_18369;
wire n_16047;
wire n_18521;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_15059;
wire n_8244;
wire n_10130;
wire n_8156;
wire n_7612;
wire n_11661;
wire n_7494;
wire n_16999;
wire n_18380;
wire n_11120;
wire n_14923;
wire n_9222;
wire n_13031;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_16391;
wire n_7736;
wire n_15949;
wire n_17071;
wire n_16040;
wire n_10622;
wire n_5633;
wire n_13661;
wire n_13155;
wire n_9546;
wire n_17912;
wire n_5664;
wire n_7589;
wire n_14259;
wire n_17764;
wire n_5921;
wire n_6797;
wire n_15673;
wire n_13410;
wire n_14012;
wire n_8759;
wire n_16941;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_13066;
wire n_8660;
wire n_13360;
wire n_11296;
wire n_13665;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_13770;
wire n_12993;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_11314;
wire n_8723;
wire n_13511;
wire n_18016;
wire n_11019;
wire n_17784;
wire n_8606;
wire n_9663;
wire n_7843;
wire n_6235;
wire n_15678;
wire n_17306;
wire n_8235;
wire n_13083;
wire n_17996;
wire n_12647;
wire n_7662;
wire n_16164;
wire n_16584;
wire n_6152;
wire n_16444;
wire n_15340;
wire n_16061;
wire n_18340;
wire n_9820;
wire n_14569;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_14071;
wire n_9743;
wire n_6496;
wire n_15744;
wire n_7756;
wire n_12749;
wire n_15557;
wire n_8342;
wire n_8940;
wire n_16776;
wire n_18244;
wire n_13048;
wire n_11584;
wire n_5280;
wire n_8448;
wire n_13563;
wire n_14154;
wire n_8472;
wire n_7700;
wire n_14169;
wire n_17905;
wire n_7555;
wire n_10000;
wire n_10158;
wire n_12812;
wire n_10582;
wire n_12066;
wire n_16151;
wire n_10427;
wire n_12060;
wire n_11816;
wire n_18254;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_14174;
wire n_7500;
wire n_6513;
wire n_10246;
wire n_11910;
wire n_15377;
wire n_16420;
wire n_11693;
wire n_18236;
wire n_15583;
wire n_15429;
wire n_13347;
wire n_15908;
wire n_14269;
wire n_5925;
wire n_9248;
wire n_8866;
wire n_5369;
wire n_8061;
wire n_6138;
wire n_9822;
wire n_10835;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_13991;
wire n_13823;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_17523;
wire n_14821;
wire n_17330;
wire n_13323;
wire n_12164;
wire n_15096;
wire n_16623;
wire n_5272;
wire n_16919;
wire n_11368;
wire n_14992;
wire n_17186;
wire n_10125;
wire n_13111;
wire n_12824;
wire n_13434;
wire n_6330;
wire n_15563;
wire n_16680;
wire n_10117;
wire n_9065;
wire n_12716;
wire n_16938;
wire n_10844;
wire n_17842;
wire n_16341;
wire n_16679;
wire n_16637;
wire n_17793;
wire n_14153;
wire n_8457;
wire n_18605;
wire n_6802;
wire n_13456;
wire n_10654;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_9339;
wire n_10198;
wire n_6909;
wire n_7157;
wire n_11064;
wire n_13237;
wire n_6908;
wire n_14312;
wire n_8237;
wire n_13445;
wire n_15448;
wire n_17177;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_15045;
wire n_11409;
wire n_16851;
wire n_18182;
wire n_15760;
wire n_7266;
wire n_16712;
wire n_17928;
wire n_8046;
wire n_14746;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_13284;
wire n_12437;
wire n_5624;
wire n_10840;
wire n_12052;
wire n_14606;
wire n_6477;
wire n_9746;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_15501;
wire n_5440;
wire n_6490;
wire n_15751;
wire n_16521;
wire n_15298;
wire n_11605;
wire n_11533;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_7198;
wire n_8335;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_17697;
wire n_9440;
wire n_10144;
wire n_17891;
wire n_9684;
wire n_17253;
wire n_15741;
wire n_16195;
wire n_6184;
wire n_14793;
wire n_15820;
wire n_5817;
wire n_18239;
wire n_5214;
wire n_15486;
wire n_10973;
wire n_13472;
wire n_15596;
wire n_17264;
wire n_9493;
wire n_15475;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_11330;
wire n_12720;
wire n_17362;
wire n_7794;
wire n_10267;
wire n_18316;
wire n_6038;
wire n_10551;
wire n_13318;
wire n_15379;
wire n_5861;
wire n_17029;
wire n_10553;
wire n_18589;
wire n_16272;
wire n_15917;
wire n_17924;
wire n_18323;
wire n_13127;
wire n_14884;
wire n_8309;
wire n_18004;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_15121;
wire n_12687;
wire n_18278;
wire n_8964;
wire n_10988;
wire n_14075;
wire n_9032;
wire n_9814;
wire n_16629;
wire n_17510;
wire n_6313;
wire n_16184;
wire n_5619;
wire n_6112;
wire n_16192;
wire n_13208;
wire n_7145;
wire n_18030;
wire n_9041;
wire n_13867;
wire n_15594;
wire n_5859;
wire n_12325;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_5380;
wire n_17841;
wire n_9245;
wire n_13443;
wire n_5776;
wire n_8166;
wire n_5606;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_14626;
wire n_5826;
wire n_15766;
wire n_18339;
wire n_16881;
wire n_10108;
wire n_18121;
wire n_8960;
wire n_13865;
wire n_12789;
wire n_5920;
wire n_10307;
wire n_16759;
wire n_14530;
wire n_17724;
wire n_15402;
wire n_7994;
wire n_14206;
wire n_17328;
wire n_18026;
wire n_8443;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_17497;
wire n_8683;
wire n_6180;
wire n_14481;
wire n_8809;
wire n_17993;
wire n_18558;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_15044;
wire n_12127;
wire n_12504;
wire n_12382;
wire n_5756;
wire n_15306;
wire n_12602;
wire n_17232;
wire n_5527;
wire n_16976;
wire n_8037;
wire n_6476;
wire n_13673;
wire n_12062;
wire n_14119;
wire n_15981;
wire n_15375;
wire n_12573;
wire n_16100;

BUFx10_ASAP7_75t_L g5169 ( 
.A(n_4361),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4343),
.Y(n_5170)
);

CKINVDCx5p33_ASAP7_75t_R g5171 ( 
.A(n_1832),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_3256),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_3605),
.Y(n_5173)
);

CKINVDCx5p33_ASAP7_75t_R g5174 ( 
.A(n_2728),
.Y(n_5174)
);

CKINVDCx5p33_ASAP7_75t_R g5175 ( 
.A(n_1950),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_2547),
.Y(n_5176)
);

CKINVDCx5p33_ASAP7_75t_R g5177 ( 
.A(n_4186),
.Y(n_5177)
);

CKINVDCx5p33_ASAP7_75t_R g5178 ( 
.A(n_2611),
.Y(n_5178)
);

BUFx5_ASAP7_75t_L g5179 ( 
.A(n_5040),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_1726),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_2881),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_2024),
.Y(n_5182)
);

CKINVDCx5p33_ASAP7_75t_R g5183 ( 
.A(n_712),
.Y(n_5183)
);

CKINVDCx5p33_ASAP7_75t_R g5184 ( 
.A(n_4363),
.Y(n_5184)
);

INVxp67_ASAP7_75t_SL g5185 ( 
.A(n_1836),
.Y(n_5185)
);

INVx1_ASAP7_75t_SL g5186 ( 
.A(n_3651),
.Y(n_5186)
);

CKINVDCx20_ASAP7_75t_R g5187 ( 
.A(n_4568),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_2170),
.Y(n_5188)
);

INVx2_ASAP7_75t_L g5189 ( 
.A(n_2245),
.Y(n_5189)
);

CKINVDCx5p33_ASAP7_75t_R g5190 ( 
.A(n_2179),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_4429),
.Y(n_5191)
);

CKINVDCx5p33_ASAP7_75t_R g5192 ( 
.A(n_2617),
.Y(n_5192)
);

CKINVDCx5p33_ASAP7_75t_R g5193 ( 
.A(n_4794),
.Y(n_5193)
);

INVx2_ASAP7_75t_SL g5194 ( 
.A(n_4052),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_1158),
.Y(n_5195)
);

CKINVDCx5p33_ASAP7_75t_R g5196 ( 
.A(n_635),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_882),
.Y(n_5197)
);

CKINVDCx5p33_ASAP7_75t_R g5198 ( 
.A(n_4796),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_4912),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_4459),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_537),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_3028),
.Y(n_5202)
);

BUFx5_ASAP7_75t_L g5203 ( 
.A(n_519),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_3331),
.Y(n_5204)
);

CKINVDCx5p33_ASAP7_75t_R g5205 ( 
.A(n_2360),
.Y(n_5205)
);

CKINVDCx5p33_ASAP7_75t_R g5206 ( 
.A(n_5154),
.Y(n_5206)
);

CKINVDCx5p33_ASAP7_75t_R g5207 ( 
.A(n_4008),
.Y(n_5207)
);

BUFx6f_ASAP7_75t_L g5208 ( 
.A(n_4470),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_2636),
.Y(n_5209)
);

CKINVDCx5p33_ASAP7_75t_R g5210 ( 
.A(n_1478),
.Y(n_5210)
);

BUFx6f_ASAP7_75t_L g5211 ( 
.A(n_677),
.Y(n_5211)
);

CKINVDCx5p33_ASAP7_75t_R g5212 ( 
.A(n_2232),
.Y(n_5212)
);

BUFx10_ASAP7_75t_L g5213 ( 
.A(n_2971),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_403),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_3163),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_1266),
.Y(n_5216)
);

CKINVDCx5p33_ASAP7_75t_R g5217 ( 
.A(n_1524),
.Y(n_5217)
);

CKINVDCx5p33_ASAP7_75t_R g5218 ( 
.A(n_2808),
.Y(n_5218)
);

CKINVDCx5p33_ASAP7_75t_R g5219 ( 
.A(n_2198),
.Y(n_5219)
);

INVx3_ASAP7_75t_L g5220 ( 
.A(n_4159),
.Y(n_5220)
);

CKINVDCx5p33_ASAP7_75t_R g5221 ( 
.A(n_4404),
.Y(n_5221)
);

INVx1_ASAP7_75t_SL g5222 ( 
.A(n_977),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4513),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_4501),
.Y(n_5224)
);

CKINVDCx5p33_ASAP7_75t_R g5225 ( 
.A(n_835),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5090),
.Y(n_5226)
);

CKINVDCx5p33_ASAP7_75t_R g5227 ( 
.A(n_3979),
.Y(n_5227)
);

BUFx2_ASAP7_75t_L g5228 ( 
.A(n_4692),
.Y(n_5228)
);

INVx2_ASAP7_75t_SL g5229 ( 
.A(n_206),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_3438),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4740),
.Y(n_5231)
);

CKINVDCx20_ASAP7_75t_R g5232 ( 
.A(n_4374),
.Y(n_5232)
);

CKINVDCx5p33_ASAP7_75t_R g5233 ( 
.A(n_4078),
.Y(n_5233)
);

BUFx6f_ASAP7_75t_L g5234 ( 
.A(n_2673),
.Y(n_5234)
);

CKINVDCx16_ASAP7_75t_R g5235 ( 
.A(n_1043),
.Y(n_5235)
);

CKINVDCx16_ASAP7_75t_R g5236 ( 
.A(n_1922),
.Y(n_5236)
);

CKINVDCx14_ASAP7_75t_R g5237 ( 
.A(n_4985),
.Y(n_5237)
);

CKINVDCx5p33_ASAP7_75t_R g5238 ( 
.A(n_4492),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_4144),
.Y(n_5239)
);

CKINVDCx5p33_ASAP7_75t_R g5240 ( 
.A(n_4494),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_1429),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4036),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_3164),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_4816),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_2287),
.Y(n_5245)
);

CKINVDCx20_ASAP7_75t_R g5246 ( 
.A(n_4078),
.Y(n_5246)
);

CKINVDCx5p33_ASAP7_75t_R g5247 ( 
.A(n_4438),
.Y(n_5247)
);

CKINVDCx5p33_ASAP7_75t_R g5248 ( 
.A(n_2137),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_2713),
.Y(n_5249)
);

CKINVDCx20_ASAP7_75t_R g5250 ( 
.A(n_902),
.Y(n_5250)
);

CKINVDCx5p33_ASAP7_75t_R g5251 ( 
.A(n_818),
.Y(n_5251)
);

CKINVDCx20_ASAP7_75t_R g5252 ( 
.A(n_3379),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_4727),
.Y(n_5253)
);

CKINVDCx5p33_ASAP7_75t_R g5254 ( 
.A(n_4665),
.Y(n_5254)
);

CKINVDCx5p33_ASAP7_75t_R g5255 ( 
.A(n_3230),
.Y(n_5255)
);

CKINVDCx5p33_ASAP7_75t_R g5256 ( 
.A(n_4141),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_3019),
.Y(n_5257)
);

CKINVDCx5p33_ASAP7_75t_R g5258 ( 
.A(n_2706),
.Y(n_5258)
);

INVx1_ASAP7_75t_SL g5259 ( 
.A(n_4554),
.Y(n_5259)
);

CKINVDCx5p33_ASAP7_75t_R g5260 ( 
.A(n_2499),
.Y(n_5260)
);

CKINVDCx5p33_ASAP7_75t_R g5261 ( 
.A(n_4406),
.Y(n_5261)
);

CKINVDCx20_ASAP7_75t_R g5262 ( 
.A(n_3992),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_2662),
.Y(n_5263)
);

CKINVDCx5p33_ASAP7_75t_R g5264 ( 
.A(n_3322),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_1500),
.Y(n_5265)
);

CKINVDCx5p33_ASAP7_75t_R g5266 ( 
.A(n_560),
.Y(n_5266)
);

INVx2_ASAP7_75t_L g5267 ( 
.A(n_4472),
.Y(n_5267)
);

CKINVDCx5p33_ASAP7_75t_R g5268 ( 
.A(n_4302),
.Y(n_5268)
);

INVx2_ASAP7_75t_SL g5269 ( 
.A(n_4217),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_4013),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_1309),
.Y(n_5271)
);

CKINVDCx5p33_ASAP7_75t_R g5272 ( 
.A(n_1561),
.Y(n_5272)
);

CKINVDCx5p33_ASAP7_75t_R g5273 ( 
.A(n_4548),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_2527),
.Y(n_5274)
);

BUFx2_ASAP7_75t_L g5275 ( 
.A(n_3607),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_4043),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_3650),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_2933),
.Y(n_5278)
);

CKINVDCx5p33_ASAP7_75t_R g5279 ( 
.A(n_4586),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_2556),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_3362),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_3352),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_670),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_4114),
.Y(n_5284)
);

INVx1_ASAP7_75t_SL g5285 ( 
.A(n_1986),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_3140),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_4510),
.Y(n_5287)
);

CKINVDCx20_ASAP7_75t_R g5288 ( 
.A(n_1861),
.Y(n_5288)
);

CKINVDCx5p33_ASAP7_75t_R g5289 ( 
.A(n_876),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_3797),
.Y(n_5290)
);

CKINVDCx5p33_ASAP7_75t_R g5291 ( 
.A(n_359),
.Y(n_5291)
);

CKINVDCx16_ASAP7_75t_R g5292 ( 
.A(n_76),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_1479),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_4255),
.Y(n_5294)
);

CKINVDCx20_ASAP7_75t_R g5295 ( 
.A(n_4553),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_151),
.Y(n_5296)
);

CKINVDCx5p33_ASAP7_75t_R g5297 ( 
.A(n_2000),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4496),
.Y(n_5298)
);

CKINVDCx20_ASAP7_75t_R g5299 ( 
.A(n_897),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_4924),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_1478),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_4152),
.Y(n_5302)
);

CKINVDCx5p33_ASAP7_75t_R g5303 ( 
.A(n_350),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_1257),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4542),
.Y(n_5305)
);

CKINVDCx20_ASAP7_75t_R g5306 ( 
.A(n_3140),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_843),
.Y(n_5307)
);

BUFx10_ASAP7_75t_L g5308 ( 
.A(n_4464),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_2927),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_4787),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4127),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_1180),
.Y(n_5312)
);

CKINVDCx5p33_ASAP7_75t_R g5313 ( 
.A(n_4574),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_1610),
.Y(n_5314)
);

CKINVDCx5p33_ASAP7_75t_R g5315 ( 
.A(n_1451),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_3100),
.Y(n_5316)
);

CKINVDCx5p33_ASAP7_75t_R g5317 ( 
.A(n_3796),
.Y(n_5317)
);

CKINVDCx5p33_ASAP7_75t_R g5318 ( 
.A(n_3566),
.Y(n_5318)
);

CKINVDCx5p33_ASAP7_75t_R g5319 ( 
.A(n_467),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_3510),
.Y(n_5320)
);

INVx2_ASAP7_75t_SL g5321 ( 
.A(n_4384),
.Y(n_5321)
);

CKINVDCx16_ASAP7_75t_R g5322 ( 
.A(n_4534),
.Y(n_5322)
);

CKINVDCx5p33_ASAP7_75t_R g5323 ( 
.A(n_2836),
.Y(n_5323)
);

CKINVDCx20_ASAP7_75t_R g5324 ( 
.A(n_768),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_4491),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_3840),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_3201),
.Y(n_5327)
);

CKINVDCx5p33_ASAP7_75t_R g5328 ( 
.A(n_1989),
.Y(n_5328)
);

CKINVDCx5p33_ASAP7_75t_R g5329 ( 
.A(n_4493),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_2371),
.Y(n_5330)
);

BUFx10_ASAP7_75t_L g5331 ( 
.A(n_2971),
.Y(n_5331)
);

CKINVDCx5p33_ASAP7_75t_R g5332 ( 
.A(n_1048),
.Y(n_5332)
);

CKINVDCx5p33_ASAP7_75t_R g5333 ( 
.A(n_4439),
.Y(n_5333)
);

CKINVDCx5p33_ASAP7_75t_R g5334 ( 
.A(n_3154),
.Y(n_5334)
);

CKINVDCx5p33_ASAP7_75t_R g5335 ( 
.A(n_420),
.Y(n_5335)
);

CKINVDCx5p33_ASAP7_75t_R g5336 ( 
.A(n_3454),
.Y(n_5336)
);

CKINVDCx5p33_ASAP7_75t_R g5337 ( 
.A(n_5032),
.Y(n_5337)
);

CKINVDCx5p33_ASAP7_75t_R g5338 ( 
.A(n_3452),
.Y(n_5338)
);

CKINVDCx5p33_ASAP7_75t_R g5339 ( 
.A(n_3102),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_2477),
.Y(n_5340)
);

CKINVDCx5p33_ASAP7_75t_R g5341 ( 
.A(n_4308),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_5152),
.Y(n_5342)
);

CKINVDCx5p33_ASAP7_75t_R g5343 ( 
.A(n_4477),
.Y(n_5343)
);

BUFx6f_ASAP7_75t_L g5344 ( 
.A(n_2347),
.Y(n_5344)
);

INVx2_ASAP7_75t_SL g5345 ( 
.A(n_4762),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_4382),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_769),
.Y(n_5347)
);

CKINVDCx5p33_ASAP7_75t_R g5348 ( 
.A(n_1874),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_4437),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_4466),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_3913),
.Y(n_5351)
);

CKINVDCx5p33_ASAP7_75t_R g5352 ( 
.A(n_2084),
.Y(n_5352)
);

BUFx10_ASAP7_75t_L g5353 ( 
.A(n_4345),
.Y(n_5353)
);

BUFx10_ASAP7_75t_L g5354 ( 
.A(n_1028),
.Y(n_5354)
);

CKINVDCx5p33_ASAP7_75t_R g5355 ( 
.A(n_3854),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_3142),
.Y(n_5356)
);

CKINVDCx5p33_ASAP7_75t_R g5357 ( 
.A(n_4580),
.Y(n_5357)
);

CKINVDCx5p33_ASAP7_75t_R g5358 ( 
.A(n_88),
.Y(n_5358)
);

CKINVDCx5p33_ASAP7_75t_R g5359 ( 
.A(n_4487),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_956),
.Y(n_5360)
);

CKINVDCx5p33_ASAP7_75t_R g5361 ( 
.A(n_4534),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4526),
.Y(n_5362)
);

CKINVDCx5p33_ASAP7_75t_R g5363 ( 
.A(n_4180),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_3738),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_4774),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_4255),
.Y(n_5366)
);

BUFx6f_ASAP7_75t_L g5367 ( 
.A(n_4520),
.Y(n_5367)
);

BUFx10_ASAP7_75t_L g5368 ( 
.A(n_4441),
.Y(n_5368)
);

CKINVDCx5p33_ASAP7_75t_R g5369 ( 
.A(n_4668),
.Y(n_5369)
);

CKINVDCx20_ASAP7_75t_R g5370 ( 
.A(n_3962),
.Y(n_5370)
);

CKINVDCx5p33_ASAP7_75t_R g5371 ( 
.A(n_5084),
.Y(n_5371)
);

CKINVDCx5p33_ASAP7_75t_R g5372 ( 
.A(n_4380),
.Y(n_5372)
);

CKINVDCx5p33_ASAP7_75t_R g5373 ( 
.A(n_4734),
.Y(n_5373)
);

INVx2_ASAP7_75t_L g5374 ( 
.A(n_4439),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_3690),
.Y(n_5375)
);

HB1xp67_ASAP7_75t_L g5376 ( 
.A(n_4461),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_3721),
.Y(n_5377)
);

CKINVDCx20_ASAP7_75t_R g5378 ( 
.A(n_2912),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_2143),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_209),
.Y(n_5380)
);

CKINVDCx20_ASAP7_75t_R g5381 ( 
.A(n_4914),
.Y(n_5381)
);

HB1xp67_ASAP7_75t_L g5382 ( 
.A(n_2270),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_1938),
.Y(n_5383)
);

CKINVDCx5p33_ASAP7_75t_R g5384 ( 
.A(n_2444),
.Y(n_5384)
);

CKINVDCx5p33_ASAP7_75t_R g5385 ( 
.A(n_4481),
.Y(n_5385)
);

CKINVDCx5p33_ASAP7_75t_R g5386 ( 
.A(n_4386),
.Y(n_5386)
);

CKINVDCx5p33_ASAP7_75t_R g5387 ( 
.A(n_469),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_912),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_1586),
.Y(n_5389)
);

CKINVDCx5p33_ASAP7_75t_R g5390 ( 
.A(n_715),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_2460),
.Y(n_5391)
);

CKINVDCx20_ASAP7_75t_R g5392 ( 
.A(n_311),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_3098),
.Y(n_5393)
);

BUFx8_ASAP7_75t_SL g5394 ( 
.A(n_4489),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_2766),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_289),
.Y(n_5396)
);

BUFx5_ASAP7_75t_L g5397 ( 
.A(n_1571),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_517),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_1157),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_191),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_3973),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_3815),
.Y(n_5402)
);

CKINVDCx16_ASAP7_75t_R g5403 ( 
.A(n_4502),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_2792),
.Y(n_5404)
);

INVx1_ASAP7_75t_SL g5405 ( 
.A(n_4612),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4460),
.Y(n_5406)
);

CKINVDCx5p33_ASAP7_75t_R g5407 ( 
.A(n_2609),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_2088),
.Y(n_5408)
);

INVx2_ASAP7_75t_L g5409 ( 
.A(n_764),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_358),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_4374),
.Y(n_5411)
);

CKINVDCx5p33_ASAP7_75t_R g5412 ( 
.A(n_5063),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_1973),
.Y(n_5413)
);

BUFx2_ASAP7_75t_L g5414 ( 
.A(n_2661),
.Y(n_5414)
);

CKINVDCx5p33_ASAP7_75t_R g5415 ( 
.A(n_627),
.Y(n_5415)
);

CKINVDCx5p33_ASAP7_75t_R g5416 ( 
.A(n_4071),
.Y(n_5416)
);

CKINVDCx5p33_ASAP7_75t_R g5417 ( 
.A(n_97),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_935),
.Y(n_5418)
);

INVx2_ASAP7_75t_SL g5419 ( 
.A(n_4000),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_4365),
.Y(n_5420)
);

CKINVDCx5p33_ASAP7_75t_R g5421 ( 
.A(n_294),
.Y(n_5421)
);

INVx1_ASAP7_75t_SL g5422 ( 
.A(n_358),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_2044),
.Y(n_5423)
);

BUFx3_ASAP7_75t_L g5424 ( 
.A(n_2334),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_4454),
.Y(n_5425)
);

BUFx10_ASAP7_75t_L g5426 ( 
.A(n_480),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_1700),
.Y(n_5427)
);

CKINVDCx5p33_ASAP7_75t_R g5428 ( 
.A(n_3787),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_4584),
.Y(n_5429)
);

CKINVDCx5p33_ASAP7_75t_R g5430 ( 
.A(n_5168),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_4414),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_3790),
.Y(n_5432)
);

CKINVDCx5p33_ASAP7_75t_R g5433 ( 
.A(n_1608),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_2310),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_2123),
.Y(n_5435)
);

CKINVDCx20_ASAP7_75t_R g5436 ( 
.A(n_4469),
.Y(n_5436)
);

CKINVDCx14_ASAP7_75t_R g5437 ( 
.A(n_926),
.Y(n_5437)
);

INVx1_ASAP7_75t_SL g5438 ( 
.A(n_3060),
.Y(n_5438)
);

CKINVDCx5p33_ASAP7_75t_R g5439 ( 
.A(n_3620),
.Y(n_5439)
);

CKINVDCx5p33_ASAP7_75t_R g5440 ( 
.A(n_1132),
.Y(n_5440)
);

CKINVDCx5p33_ASAP7_75t_R g5441 ( 
.A(n_4177),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_4546),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_2555),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_1560),
.Y(n_5444)
);

CKINVDCx5p33_ASAP7_75t_R g5445 ( 
.A(n_3775),
.Y(n_5445)
);

CKINVDCx20_ASAP7_75t_R g5446 ( 
.A(n_2980),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_3145),
.Y(n_5447)
);

CKINVDCx5p33_ASAP7_75t_R g5448 ( 
.A(n_1135),
.Y(n_5448)
);

CKINVDCx5p33_ASAP7_75t_R g5449 ( 
.A(n_2804),
.Y(n_5449)
);

BUFx3_ASAP7_75t_L g5450 ( 
.A(n_242),
.Y(n_5450)
);

CKINVDCx5p33_ASAP7_75t_R g5451 ( 
.A(n_281),
.Y(n_5451)
);

INVx2_ASAP7_75t_L g5452 ( 
.A(n_4376),
.Y(n_5452)
);

CKINVDCx5p33_ASAP7_75t_R g5453 ( 
.A(n_4479),
.Y(n_5453)
);

BUFx8_ASAP7_75t_SL g5454 ( 
.A(n_3831),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_3101),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_2275),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_1806),
.Y(n_5457)
);

CKINVDCx5p33_ASAP7_75t_R g5458 ( 
.A(n_3536),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_3938),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_4388),
.Y(n_5460)
);

CKINVDCx20_ASAP7_75t_R g5461 ( 
.A(n_913),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_1447),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_824),
.Y(n_5463)
);

BUFx6f_ASAP7_75t_L g5464 ( 
.A(n_3817),
.Y(n_5464)
);

CKINVDCx5p33_ASAP7_75t_R g5465 ( 
.A(n_4364),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_2373),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_3966),
.Y(n_5467)
);

INVx2_ASAP7_75t_SL g5468 ( 
.A(n_1500),
.Y(n_5468)
);

CKINVDCx20_ASAP7_75t_R g5469 ( 
.A(n_162),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_4392),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_861),
.Y(n_5471)
);

CKINVDCx5p33_ASAP7_75t_R g5472 ( 
.A(n_262),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_1009),
.Y(n_5473)
);

CKINVDCx5p33_ASAP7_75t_R g5474 ( 
.A(n_1901),
.Y(n_5474)
);

CKINVDCx5p33_ASAP7_75t_R g5475 ( 
.A(n_3171),
.Y(n_5475)
);

CKINVDCx5p33_ASAP7_75t_R g5476 ( 
.A(n_4913),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_276),
.Y(n_5477)
);

CKINVDCx5p33_ASAP7_75t_R g5478 ( 
.A(n_1064),
.Y(n_5478)
);

CKINVDCx20_ASAP7_75t_R g5479 ( 
.A(n_4555),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_4430),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_628),
.Y(n_5481)
);

INVx1_ASAP7_75t_SL g5482 ( 
.A(n_621),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_3347),
.Y(n_5483)
);

CKINVDCx20_ASAP7_75t_R g5484 ( 
.A(n_4262),
.Y(n_5484)
);

BUFx6f_ASAP7_75t_L g5485 ( 
.A(n_4454),
.Y(n_5485)
);

INVxp67_ASAP7_75t_SL g5486 ( 
.A(n_4366),
.Y(n_5486)
);

CKINVDCx5p33_ASAP7_75t_R g5487 ( 
.A(n_2377),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_3228),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_4860),
.Y(n_5489)
);

CKINVDCx20_ASAP7_75t_R g5490 ( 
.A(n_1827),
.Y(n_5490)
);

CKINVDCx5p33_ASAP7_75t_R g5491 ( 
.A(n_1291),
.Y(n_5491)
);

CKINVDCx5p33_ASAP7_75t_R g5492 ( 
.A(n_199),
.Y(n_5492)
);

CKINVDCx5p33_ASAP7_75t_R g5493 ( 
.A(n_4284),
.Y(n_5493)
);

CKINVDCx5p33_ASAP7_75t_R g5494 ( 
.A(n_3649),
.Y(n_5494)
);

BUFx3_ASAP7_75t_L g5495 ( 
.A(n_4605),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_3024),
.Y(n_5496)
);

CKINVDCx5p33_ASAP7_75t_R g5497 ( 
.A(n_4292),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_485),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_1108),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_2368),
.Y(n_5500)
);

BUFx6f_ASAP7_75t_L g5501 ( 
.A(n_4649),
.Y(n_5501)
);

BUFx10_ASAP7_75t_L g5502 ( 
.A(n_4413),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_3496),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_3726),
.Y(n_5504)
);

INVx1_ASAP7_75t_SL g5505 ( 
.A(n_3841),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_4098),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_494),
.Y(n_5507)
);

CKINVDCx5p33_ASAP7_75t_R g5508 ( 
.A(n_4833),
.Y(n_5508)
);

CKINVDCx5p33_ASAP7_75t_R g5509 ( 
.A(n_1525),
.Y(n_5509)
);

INVxp67_ASAP7_75t_L g5510 ( 
.A(n_4372),
.Y(n_5510)
);

CKINVDCx5p33_ASAP7_75t_R g5511 ( 
.A(n_1080),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_4716),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_1182),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_1858),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_1379),
.Y(n_5515)
);

CKINVDCx14_ASAP7_75t_R g5516 ( 
.A(n_1595),
.Y(n_5516)
);

INVx1_ASAP7_75t_SL g5517 ( 
.A(n_5159),
.Y(n_5517)
);

CKINVDCx5p33_ASAP7_75t_R g5518 ( 
.A(n_1587),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_1454),
.Y(n_5519)
);

BUFx10_ASAP7_75t_L g5520 ( 
.A(n_2209),
.Y(n_5520)
);

CKINVDCx5p33_ASAP7_75t_R g5521 ( 
.A(n_1995),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_2961),
.Y(n_5522)
);

BUFx6f_ASAP7_75t_L g5523 ( 
.A(n_2524),
.Y(n_5523)
);

CKINVDCx5p33_ASAP7_75t_R g5524 ( 
.A(n_2400),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_4574),
.Y(n_5525)
);

CKINVDCx5p33_ASAP7_75t_R g5526 ( 
.A(n_1685),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_4143),
.Y(n_5527)
);

CKINVDCx5p33_ASAP7_75t_R g5528 ( 
.A(n_1094),
.Y(n_5528)
);

INVx1_ASAP7_75t_SL g5529 ( 
.A(n_1279),
.Y(n_5529)
);

INVx1_ASAP7_75t_SL g5530 ( 
.A(n_3398),
.Y(n_5530)
);

BUFx10_ASAP7_75t_L g5531 ( 
.A(n_1739),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_2648),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_4494),
.Y(n_5533)
);

BUFx8_ASAP7_75t_SL g5534 ( 
.A(n_4431),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_2395),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_472),
.Y(n_5536)
);

BUFx3_ASAP7_75t_L g5537 ( 
.A(n_1226),
.Y(n_5537)
);

CKINVDCx5p33_ASAP7_75t_R g5538 ( 
.A(n_1851),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_3118),
.Y(n_5539)
);

CKINVDCx5p33_ASAP7_75t_R g5540 ( 
.A(n_2501),
.Y(n_5540)
);

CKINVDCx5p33_ASAP7_75t_R g5541 ( 
.A(n_2098),
.Y(n_5541)
);

CKINVDCx5p33_ASAP7_75t_R g5542 ( 
.A(n_4614),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_3639),
.Y(n_5543)
);

CKINVDCx5p33_ASAP7_75t_R g5544 ( 
.A(n_3524),
.Y(n_5544)
);

CKINVDCx5p33_ASAP7_75t_R g5545 ( 
.A(n_1856),
.Y(n_5545)
);

BUFx3_ASAP7_75t_L g5546 ( 
.A(n_2261),
.Y(n_5546)
);

CKINVDCx5p33_ASAP7_75t_R g5547 ( 
.A(n_3378),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_2653),
.Y(n_5548)
);

INVx2_ASAP7_75t_SL g5549 ( 
.A(n_4975),
.Y(n_5549)
);

CKINVDCx5p33_ASAP7_75t_R g5550 ( 
.A(n_3404),
.Y(n_5550)
);

CKINVDCx20_ASAP7_75t_R g5551 ( 
.A(n_1094),
.Y(n_5551)
);

CKINVDCx5p33_ASAP7_75t_R g5552 ( 
.A(n_4123),
.Y(n_5552)
);

CKINVDCx5p33_ASAP7_75t_R g5553 ( 
.A(n_2180),
.Y(n_5553)
);

CKINVDCx5p33_ASAP7_75t_R g5554 ( 
.A(n_41),
.Y(n_5554)
);

CKINVDCx5p33_ASAP7_75t_R g5555 ( 
.A(n_3160),
.Y(n_5555)
);

CKINVDCx20_ASAP7_75t_R g5556 ( 
.A(n_2009),
.Y(n_5556)
);

CKINVDCx5p33_ASAP7_75t_R g5557 ( 
.A(n_873),
.Y(n_5557)
);

CKINVDCx20_ASAP7_75t_R g5558 ( 
.A(n_1192),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_1099),
.Y(n_5559)
);

CKINVDCx5p33_ASAP7_75t_R g5560 ( 
.A(n_1138),
.Y(n_5560)
);

CKINVDCx16_ASAP7_75t_R g5561 ( 
.A(n_4475),
.Y(n_5561)
);

BUFx8_ASAP7_75t_SL g5562 ( 
.A(n_1097),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_15),
.Y(n_5563)
);

CKINVDCx5p33_ASAP7_75t_R g5564 ( 
.A(n_3663),
.Y(n_5564)
);

CKINVDCx5p33_ASAP7_75t_R g5565 ( 
.A(n_605),
.Y(n_5565)
);

CKINVDCx5p33_ASAP7_75t_R g5566 ( 
.A(n_1166),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_536),
.Y(n_5567)
);

INVxp33_ASAP7_75t_R g5568 ( 
.A(n_2235),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_2833),
.Y(n_5569)
);

BUFx6f_ASAP7_75t_L g5570 ( 
.A(n_4517),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_3917),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_1298),
.Y(n_5572)
);

CKINVDCx5p33_ASAP7_75t_R g5573 ( 
.A(n_4385),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_4105),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_2521),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_1588),
.Y(n_5576)
);

CKINVDCx5p33_ASAP7_75t_R g5577 ( 
.A(n_3384),
.Y(n_5577)
);

CKINVDCx5p33_ASAP7_75t_R g5578 ( 
.A(n_3171),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_4725),
.Y(n_5579)
);

CKINVDCx5p33_ASAP7_75t_R g5580 ( 
.A(n_3106),
.Y(n_5580)
);

INVx2_ASAP7_75t_L g5581 ( 
.A(n_4378),
.Y(n_5581)
);

CKINVDCx5p33_ASAP7_75t_R g5582 ( 
.A(n_487),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_4310),
.Y(n_5583)
);

CKINVDCx5p33_ASAP7_75t_R g5584 ( 
.A(n_5137),
.Y(n_5584)
);

CKINVDCx5p33_ASAP7_75t_R g5585 ( 
.A(n_4095),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_1111),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_3883),
.Y(n_5587)
);

CKINVDCx5p33_ASAP7_75t_R g5588 ( 
.A(n_1400),
.Y(n_5588)
);

CKINVDCx5p33_ASAP7_75t_R g5589 ( 
.A(n_4082),
.Y(n_5589)
);

CKINVDCx5p33_ASAP7_75t_R g5590 ( 
.A(n_1606),
.Y(n_5590)
);

CKINVDCx20_ASAP7_75t_R g5591 ( 
.A(n_1546),
.Y(n_5591)
);

CKINVDCx5p33_ASAP7_75t_R g5592 ( 
.A(n_2140),
.Y(n_5592)
);

CKINVDCx5p33_ASAP7_75t_R g5593 ( 
.A(n_4390),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_4399),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_4237),
.Y(n_5595)
);

CKINVDCx5p33_ASAP7_75t_R g5596 ( 
.A(n_3918),
.Y(n_5596)
);

CKINVDCx5p33_ASAP7_75t_R g5597 ( 
.A(n_432),
.Y(n_5597)
);

CKINVDCx5p33_ASAP7_75t_R g5598 ( 
.A(n_2281),
.Y(n_5598)
);

INVx1_ASAP7_75t_SL g5599 ( 
.A(n_1260),
.Y(n_5599)
);

CKINVDCx5p33_ASAP7_75t_R g5600 ( 
.A(n_3571),
.Y(n_5600)
);

CKINVDCx5p33_ASAP7_75t_R g5601 ( 
.A(n_3409),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_4314),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_2435),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_1421),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_163),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_4756),
.Y(n_5606)
);

CKINVDCx5p33_ASAP7_75t_R g5607 ( 
.A(n_3496),
.Y(n_5607)
);

CKINVDCx5p33_ASAP7_75t_R g5608 ( 
.A(n_4533),
.Y(n_5608)
);

CKINVDCx5p33_ASAP7_75t_R g5609 ( 
.A(n_1964),
.Y(n_5609)
);

CKINVDCx5p33_ASAP7_75t_R g5610 ( 
.A(n_248),
.Y(n_5610)
);

INVxp67_ASAP7_75t_L g5611 ( 
.A(n_3863),
.Y(n_5611)
);

BUFx3_ASAP7_75t_L g5612 ( 
.A(n_3128),
.Y(n_5612)
);

BUFx5_ASAP7_75t_L g5613 ( 
.A(n_4403),
.Y(n_5613)
);

CKINVDCx5p33_ASAP7_75t_R g5614 ( 
.A(n_4278),
.Y(n_5614)
);

BUFx6f_ASAP7_75t_L g5615 ( 
.A(n_795),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_4498),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_1188),
.Y(n_5617)
);

INVx1_ASAP7_75t_SL g5618 ( 
.A(n_2200),
.Y(n_5618)
);

INVxp67_ASAP7_75t_L g5619 ( 
.A(n_288),
.Y(n_5619)
);

BUFx3_ASAP7_75t_L g5620 ( 
.A(n_3052),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_950),
.Y(n_5621)
);

CKINVDCx5p33_ASAP7_75t_R g5622 ( 
.A(n_466),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_4452),
.Y(n_5623)
);

INVxp67_ASAP7_75t_SL g5624 ( 
.A(n_3206),
.Y(n_5624)
);

CKINVDCx5p33_ASAP7_75t_R g5625 ( 
.A(n_4258),
.Y(n_5625)
);

CKINVDCx5p33_ASAP7_75t_R g5626 ( 
.A(n_4395),
.Y(n_5626)
);

CKINVDCx5p33_ASAP7_75t_R g5627 ( 
.A(n_2843),
.Y(n_5627)
);

CKINVDCx5p33_ASAP7_75t_R g5628 ( 
.A(n_803),
.Y(n_5628)
);

INVxp67_ASAP7_75t_L g5629 ( 
.A(n_4696),
.Y(n_5629)
);

CKINVDCx5p33_ASAP7_75t_R g5630 ( 
.A(n_1567),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_2475),
.Y(n_5631)
);

INVx1_ASAP7_75t_SL g5632 ( 
.A(n_3350),
.Y(n_5632)
);

CKINVDCx5p33_ASAP7_75t_R g5633 ( 
.A(n_4434),
.Y(n_5633)
);

INVx1_ASAP7_75t_SL g5634 ( 
.A(n_4042),
.Y(n_5634)
);

CKINVDCx5p33_ASAP7_75t_R g5635 ( 
.A(n_1140),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_2753),
.Y(n_5636)
);

INVx2_ASAP7_75t_SL g5637 ( 
.A(n_1649),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_4171),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_3752),
.Y(n_5639)
);

INVx1_ASAP7_75t_SL g5640 ( 
.A(n_4308),
.Y(n_5640)
);

CKINVDCx5p33_ASAP7_75t_R g5641 ( 
.A(n_2093),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_666),
.Y(n_5642)
);

CKINVDCx5p33_ASAP7_75t_R g5643 ( 
.A(n_1270),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_4398),
.Y(n_5644)
);

BUFx10_ASAP7_75t_L g5645 ( 
.A(n_2),
.Y(n_5645)
);

INVx2_ASAP7_75t_L g5646 ( 
.A(n_4370),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_4440),
.Y(n_5647)
);

CKINVDCx20_ASAP7_75t_R g5648 ( 
.A(n_4405),
.Y(n_5648)
);

CKINVDCx5p33_ASAP7_75t_R g5649 ( 
.A(n_1907),
.Y(n_5649)
);

CKINVDCx20_ASAP7_75t_R g5650 ( 
.A(n_4266),
.Y(n_5650)
);

INVxp33_ASAP7_75t_L g5651 ( 
.A(n_4549),
.Y(n_5651)
);

CKINVDCx5p33_ASAP7_75t_R g5652 ( 
.A(n_3603),
.Y(n_5652)
);

CKINVDCx20_ASAP7_75t_R g5653 ( 
.A(n_4449),
.Y(n_5653)
);

CKINVDCx5p33_ASAP7_75t_R g5654 ( 
.A(n_5085),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_2947),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_3803),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_4693),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_2719),
.Y(n_5658)
);

CKINVDCx20_ASAP7_75t_R g5659 ( 
.A(n_2782),
.Y(n_5659)
);

CKINVDCx5p33_ASAP7_75t_R g5660 ( 
.A(n_1536),
.Y(n_5660)
);

CKINVDCx5p33_ASAP7_75t_R g5661 ( 
.A(n_4478),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_2079),
.Y(n_5662)
);

CKINVDCx20_ASAP7_75t_R g5663 ( 
.A(n_1347),
.Y(n_5663)
);

BUFx3_ASAP7_75t_L g5664 ( 
.A(n_2049),
.Y(n_5664)
);

CKINVDCx20_ASAP7_75t_R g5665 ( 
.A(n_4401),
.Y(n_5665)
);

CKINVDCx5p33_ASAP7_75t_R g5666 ( 
.A(n_2475),
.Y(n_5666)
);

CKINVDCx5p33_ASAP7_75t_R g5667 ( 
.A(n_2408),
.Y(n_5667)
);

INVx1_ASAP7_75t_L g5668 ( 
.A(n_1037),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_2250),
.Y(n_5669)
);

INVx1_ASAP7_75t_SL g5670 ( 
.A(n_4123),
.Y(n_5670)
);

CKINVDCx5p33_ASAP7_75t_R g5671 ( 
.A(n_4381),
.Y(n_5671)
);

CKINVDCx5p33_ASAP7_75t_R g5672 ( 
.A(n_4776),
.Y(n_5672)
);

INVxp33_ASAP7_75t_SL g5673 ( 
.A(n_1641),
.Y(n_5673)
);

CKINVDCx5p33_ASAP7_75t_R g5674 ( 
.A(n_610),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_575),
.Y(n_5675)
);

BUFx3_ASAP7_75t_L g5676 ( 
.A(n_4452),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_514),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_2303),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_1061),
.Y(n_5679)
);

INVx1_ASAP7_75t_SL g5680 ( 
.A(n_3218),
.Y(n_5680)
);

CKINVDCx5p33_ASAP7_75t_R g5681 ( 
.A(n_2613),
.Y(n_5681)
);

BUFx2_ASAP7_75t_L g5682 ( 
.A(n_1870),
.Y(n_5682)
);

BUFx3_ASAP7_75t_L g5683 ( 
.A(n_4267),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_2919),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_2260),
.Y(n_5685)
);

CKINVDCx5p33_ASAP7_75t_R g5686 ( 
.A(n_3007),
.Y(n_5686)
);

BUFx6f_ASAP7_75t_L g5687 ( 
.A(n_4378),
.Y(n_5687)
);

CKINVDCx20_ASAP7_75t_R g5688 ( 
.A(n_4713),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_765),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_4362),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_2678),
.Y(n_5691)
);

CKINVDCx20_ASAP7_75t_R g5692 ( 
.A(n_422),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_790),
.Y(n_5693)
);

CKINVDCx5p33_ASAP7_75t_R g5694 ( 
.A(n_3024),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_4422),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_4847),
.Y(n_5696)
);

CKINVDCx5p33_ASAP7_75t_R g5697 ( 
.A(n_4346),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_620),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_2318),
.Y(n_5699)
);

INVxp67_ASAP7_75t_SL g5700 ( 
.A(n_3078),
.Y(n_5700)
);

CKINVDCx5p33_ASAP7_75t_R g5701 ( 
.A(n_3326),
.Y(n_5701)
);

INVxp67_ASAP7_75t_SL g5702 ( 
.A(n_3058),
.Y(n_5702)
);

INVx3_ASAP7_75t_L g5703 ( 
.A(n_1442),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_4135),
.Y(n_5704)
);

CKINVDCx20_ASAP7_75t_R g5705 ( 
.A(n_4402),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_643),
.Y(n_5706)
);

BUFx10_ASAP7_75t_L g5707 ( 
.A(n_2207),
.Y(n_5707)
);

CKINVDCx5p33_ASAP7_75t_R g5708 ( 
.A(n_4309),
.Y(n_5708)
);

CKINVDCx20_ASAP7_75t_R g5709 ( 
.A(n_3596),
.Y(n_5709)
);

BUFx2_ASAP7_75t_L g5710 ( 
.A(n_2514),
.Y(n_5710)
);

BUFx6f_ASAP7_75t_L g5711 ( 
.A(n_268),
.Y(n_5711)
);

CKINVDCx5p33_ASAP7_75t_R g5712 ( 
.A(n_4606),
.Y(n_5712)
);

CKINVDCx5p33_ASAP7_75t_R g5713 ( 
.A(n_4447),
.Y(n_5713)
);

INVx1_ASAP7_75t_SL g5714 ( 
.A(n_1563),
.Y(n_5714)
);

CKINVDCx5p33_ASAP7_75t_R g5715 ( 
.A(n_3833),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_1745),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_3890),
.Y(n_5717)
);

CKINVDCx5p33_ASAP7_75t_R g5718 ( 
.A(n_1494),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_3966),
.Y(n_5719)
);

CKINVDCx5p33_ASAP7_75t_R g5720 ( 
.A(n_1040),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_3545),
.Y(n_5721)
);

CKINVDCx14_ASAP7_75t_R g5722 ( 
.A(n_3654),
.Y(n_5722)
);

CKINVDCx5p33_ASAP7_75t_R g5723 ( 
.A(n_4528),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_2098),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_4436),
.Y(n_5725)
);

CKINVDCx20_ASAP7_75t_R g5726 ( 
.A(n_4602),
.Y(n_5726)
);

CKINVDCx5p33_ASAP7_75t_R g5727 ( 
.A(n_4680),
.Y(n_5727)
);

CKINVDCx5p33_ASAP7_75t_R g5728 ( 
.A(n_2846),
.Y(n_5728)
);

CKINVDCx5p33_ASAP7_75t_R g5729 ( 
.A(n_2323),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_3621),
.Y(n_5730)
);

CKINVDCx5p33_ASAP7_75t_R g5731 ( 
.A(n_2123),
.Y(n_5731)
);

INVxp67_ASAP7_75t_L g5732 ( 
.A(n_1838),
.Y(n_5732)
);

CKINVDCx5p33_ASAP7_75t_R g5733 ( 
.A(n_4629),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_1092),
.Y(n_5734)
);

BUFx6f_ASAP7_75t_L g5735 ( 
.A(n_2473),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_57),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_4427),
.Y(n_5737)
);

CKINVDCx16_ASAP7_75t_R g5738 ( 
.A(n_64),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_4165),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_3254),
.Y(n_5740)
);

CKINVDCx5p33_ASAP7_75t_R g5741 ( 
.A(n_4709),
.Y(n_5741)
);

BUFx6f_ASAP7_75t_L g5742 ( 
.A(n_4398),
.Y(n_5742)
);

CKINVDCx5p33_ASAP7_75t_R g5743 ( 
.A(n_4479),
.Y(n_5743)
);

INVxp67_ASAP7_75t_L g5744 ( 
.A(n_2877),
.Y(n_5744)
);

CKINVDCx5p33_ASAP7_75t_R g5745 ( 
.A(n_4412),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_3445),
.Y(n_5746)
);

BUFx5_ASAP7_75t_L g5747 ( 
.A(n_1475),
.Y(n_5747)
);

CKINVDCx5p33_ASAP7_75t_R g5748 ( 
.A(n_377),
.Y(n_5748)
);

CKINVDCx5p33_ASAP7_75t_R g5749 ( 
.A(n_3197),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_4120),
.Y(n_5750)
);

BUFx10_ASAP7_75t_L g5751 ( 
.A(n_2361),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_2963),
.Y(n_5752)
);

CKINVDCx5p33_ASAP7_75t_R g5753 ( 
.A(n_2711),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_4465),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_4639),
.Y(n_5755)
);

CKINVDCx5p33_ASAP7_75t_R g5756 ( 
.A(n_4537),
.Y(n_5756)
);

BUFx6f_ASAP7_75t_L g5757 ( 
.A(n_2917),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_1546),
.Y(n_5758)
);

CKINVDCx5p33_ASAP7_75t_R g5759 ( 
.A(n_2530),
.Y(n_5759)
);

CKINVDCx5p33_ASAP7_75t_R g5760 ( 
.A(n_3975),
.Y(n_5760)
);

CKINVDCx5p33_ASAP7_75t_R g5761 ( 
.A(n_4184),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_4932),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_3581),
.Y(n_5763)
);

CKINVDCx5p33_ASAP7_75t_R g5764 ( 
.A(n_2319),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_4264),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_4387),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_3894),
.Y(n_5767)
);

CKINVDCx5p33_ASAP7_75t_R g5768 ( 
.A(n_3056),
.Y(n_5768)
);

CKINVDCx20_ASAP7_75t_R g5769 ( 
.A(n_2790),
.Y(n_5769)
);

INVx1_ASAP7_75t_SL g5770 ( 
.A(n_4761),
.Y(n_5770)
);

CKINVDCx5p33_ASAP7_75t_R g5771 ( 
.A(n_4213),
.Y(n_5771)
);

CKINVDCx5p33_ASAP7_75t_R g5772 ( 
.A(n_3010),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_4946),
.Y(n_5773)
);

BUFx2_ASAP7_75t_L g5774 ( 
.A(n_4456),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_4125),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_3723),
.Y(n_5776)
);

INVx2_ASAP7_75t_SL g5777 ( 
.A(n_4279),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_4664),
.Y(n_5778)
);

CKINVDCx5p33_ASAP7_75t_R g5779 ( 
.A(n_2160),
.Y(n_5779)
);

CKINVDCx5p33_ASAP7_75t_R g5780 ( 
.A(n_4770),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_1092),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_4578),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_54),
.Y(n_5783)
);

BUFx3_ASAP7_75t_L g5784 ( 
.A(n_5056),
.Y(n_5784)
);

CKINVDCx5p33_ASAP7_75t_R g5785 ( 
.A(n_1356),
.Y(n_5785)
);

BUFx10_ASAP7_75t_L g5786 ( 
.A(n_2314),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_1623),
.Y(n_5787)
);

CKINVDCx5p33_ASAP7_75t_R g5788 ( 
.A(n_1016),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_4426),
.Y(n_5789)
);

CKINVDCx20_ASAP7_75t_R g5790 ( 
.A(n_3909),
.Y(n_5790)
);

CKINVDCx5p33_ASAP7_75t_R g5791 ( 
.A(n_2633),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_3567),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_498),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_1758),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_2199),
.Y(n_5795)
);

CKINVDCx5p33_ASAP7_75t_R g5796 ( 
.A(n_1723),
.Y(n_5796)
);

CKINVDCx5p33_ASAP7_75t_R g5797 ( 
.A(n_3829),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_1327),
.Y(n_5798)
);

CKINVDCx5p33_ASAP7_75t_R g5799 ( 
.A(n_4371),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_3313),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_4480),
.Y(n_5801)
);

INVxp67_ASAP7_75t_L g5802 ( 
.A(n_1049),
.Y(n_5802)
);

CKINVDCx5p33_ASAP7_75t_R g5803 ( 
.A(n_156),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_970),
.Y(n_5804)
);

CKINVDCx5p33_ASAP7_75t_R g5805 ( 
.A(n_3293),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_2692),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_3701),
.Y(n_5807)
);

INVx2_ASAP7_75t_L g5808 ( 
.A(n_3042),
.Y(n_5808)
);

INVx1_ASAP7_75t_SL g5809 ( 
.A(n_4710),
.Y(n_5809)
);

CKINVDCx5p33_ASAP7_75t_R g5810 ( 
.A(n_2169),
.Y(n_5810)
);

CKINVDCx5p33_ASAP7_75t_R g5811 ( 
.A(n_4758),
.Y(n_5811)
);

CKINVDCx5p33_ASAP7_75t_R g5812 ( 
.A(n_4726),
.Y(n_5812)
);

CKINVDCx20_ASAP7_75t_R g5813 ( 
.A(n_4580),
.Y(n_5813)
);

BUFx3_ASAP7_75t_L g5814 ( 
.A(n_1221),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_4531),
.Y(n_5815)
);

BUFx3_ASAP7_75t_L g5816 ( 
.A(n_3018),
.Y(n_5816)
);

CKINVDCx5p33_ASAP7_75t_R g5817 ( 
.A(n_1167),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_3919),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_166),
.Y(n_5819)
);

BUFx6f_ASAP7_75t_L g5820 ( 
.A(n_1133),
.Y(n_5820)
);

CKINVDCx5p33_ASAP7_75t_R g5821 ( 
.A(n_456),
.Y(n_5821)
);

CKINVDCx5p33_ASAP7_75t_R g5822 ( 
.A(n_2704),
.Y(n_5822)
);

CKINVDCx5p33_ASAP7_75t_R g5823 ( 
.A(n_5158),
.Y(n_5823)
);

BUFx6f_ASAP7_75t_L g5824 ( 
.A(n_1569),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_1172),
.Y(n_5825)
);

BUFx6f_ASAP7_75t_L g5826 ( 
.A(n_1292),
.Y(n_5826)
);

CKINVDCx16_ASAP7_75t_R g5827 ( 
.A(n_119),
.Y(n_5827)
);

INVx1_ASAP7_75t_SL g5828 ( 
.A(n_2),
.Y(n_5828)
);

CKINVDCx5p33_ASAP7_75t_R g5829 ( 
.A(n_740),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_3972),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_1842),
.Y(n_5831)
);

CKINVDCx5p33_ASAP7_75t_R g5832 ( 
.A(n_4260),
.Y(n_5832)
);

CKINVDCx5p33_ASAP7_75t_R g5833 ( 
.A(n_2095),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_467),
.Y(n_5834)
);

CKINVDCx5p33_ASAP7_75t_R g5835 ( 
.A(n_2224),
.Y(n_5835)
);

BUFx8_ASAP7_75t_SL g5836 ( 
.A(n_2801),
.Y(n_5836)
);

CKINVDCx5p33_ASAP7_75t_R g5837 ( 
.A(n_3392),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_4488),
.Y(n_5838)
);

CKINVDCx5p33_ASAP7_75t_R g5839 ( 
.A(n_4423),
.Y(n_5839)
);

INVxp67_ASAP7_75t_SL g5840 ( 
.A(n_2859),
.Y(n_5840)
);

CKINVDCx5p33_ASAP7_75t_R g5841 ( 
.A(n_1898),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_1715),
.Y(n_5842)
);

CKINVDCx5p33_ASAP7_75t_R g5843 ( 
.A(n_3263),
.Y(n_5843)
);

CKINVDCx5p33_ASAP7_75t_R g5844 ( 
.A(n_3547),
.Y(n_5844)
);

CKINVDCx5p33_ASAP7_75t_R g5845 ( 
.A(n_4457),
.Y(n_5845)
);

CKINVDCx5p33_ASAP7_75t_R g5846 ( 
.A(n_1185),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_3637),
.Y(n_5847)
);

CKINVDCx5p33_ASAP7_75t_R g5848 ( 
.A(n_2785),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_2700),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_4139),
.Y(n_5850)
);

CKINVDCx20_ASAP7_75t_R g5851 ( 
.A(n_4383),
.Y(n_5851)
);

BUFx2_ASAP7_75t_L g5852 ( 
.A(n_4186),
.Y(n_5852)
);

BUFx5_ASAP7_75t_L g5853 ( 
.A(n_597),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_2932),
.Y(n_5854)
);

INVx1_ASAP7_75t_SL g5855 ( 
.A(n_1271),
.Y(n_5855)
);

CKINVDCx16_ASAP7_75t_R g5856 ( 
.A(n_1184),
.Y(n_5856)
);

CKINVDCx5p33_ASAP7_75t_R g5857 ( 
.A(n_4346),
.Y(n_5857)
);

BUFx3_ASAP7_75t_L g5858 ( 
.A(n_4317),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_664),
.Y(n_5859)
);

CKINVDCx5p33_ASAP7_75t_R g5860 ( 
.A(n_4421),
.Y(n_5860)
);

CKINVDCx5p33_ASAP7_75t_R g5861 ( 
.A(n_232),
.Y(n_5861)
);

BUFx2_ASAP7_75t_SL g5862 ( 
.A(n_4337),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5053),
.Y(n_5863)
);

CKINVDCx5p33_ASAP7_75t_R g5864 ( 
.A(n_3103),
.Y(n_5864)
);

CKINVDCx5p33_ASAP7_75t_R g5865 ( 
.A(n_4486),
.Y(n_5865)
);

CKINVDCx5p33_ASAP7_75t_R g5866 ( 
.A(n_5076),
.Y(n_5866)
);

CKINVDCx20_ASAP7_75t_R g5867 ( 
.A(n_2552),
.Y(n_5867)
);

CKINVDCx5p33_ASAP7_75t_R g5868 ( 
.A(n_563),
.Y(n_5868)
);

CKINVDCx5p33_ASAP7_75t_R g5869 ( 
.A(n_4511),
.Y(n_5869)
);

CKINVDCx5p33_ASAP7_75t_R g5870 ( 
.A(n_1623),
.Y(n_5870)
);

CKINVDCx5p33_ASAP7_75t_R g5871 ( 
.A(n_4462),
.Y(n_5871)
);

CKINVDCx5p33_ASAP7_75t_R g5872 ( 
.A(n_3980),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_4407),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_1017),
.Y(n_5874)
);

CKINVDCx20_ASAP7_75t_R g5875 ( 
.A(n_4768),
.Y(n_5875)
);

CKINVDCx5p33_ASAP7_75t_R g5876 ( 
.A(n_4191),
.Y(n_5876)
);

CKINVDCx5p33_ASAP7_75t_R g5877 ( 
.A(n_350),
.Y(n_5877)
);

CKINVDCx5p33_ASAP7_75t_R g5878 ( 
.A(n_2783),
.Y(n_5878)
);

CKINVDCx20_ASAP7_75t_R g5879 ( 
.A(n_175),
.Y(n_5879)
);

CKINVDCx5p33_ASAP7_75t_R g5880 ( 
.A(n_1061),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_4415),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_3731),
.Y(n_5882)
);

CKINVDCx5p33_ASAP7_75t_R g5883 ( 
.A(n_5165),
.Y(n_5883)
);

CKINVDCx5p33_ASAP7_75t_R g5884 ( 
.A(n_4362),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_347),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_2504),
.Y(n_5886)
);

CKINVDCx5p33_ASAP7_75t_R g5887 ( 
.A(n_693),
.Y(n_5887)
);

CKINVDCx5p33_ASAP7_75t_R g5888 ( 
.A(n_4947),
.Y(n_5888)
);

INVx1_ASAP7_75t_SL g5889 ( 
.A(n_3826),
.Y(n_5889)
);

BUFx2_ASAP7_75t_L g5890 ( 
.A(n_2776),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_1320),
.Y(n_5891)
);

CKINVDCx5p33_ASAP7_75t_R g5892 ( 
.A(n_2549),
.Y(n_5892)
);

CKINVDCx5p33_ASAP7_75t_R g5893 ( 
.A(n_4540),
.Y(n_5893)
);

INVx1_ASAP7_75t_SL g5894 ( 
.A(n_1566),
.Y(n_5894)
);

BUFx8_ASAP7_75t_SL g5895 ( 
.A(n_3187),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_21),
.Y(n_5896)
);

HB1xp67_ASAP7_75t_L g5897 ( 
.A(n_1985),
.Y(n_5897)
);

INVx1_ASAP7_75t_SL g5898 ( 
.A(n_1968),
.Y(n_5898)
);

CKINVDCx5p33_ASAP7_75t_R g5899 ( 
.A(n_1112),
.Y(n_5899)
);

CKINVDCx5p33_ASAP7_75t_R g5900 ( 
.A(n_3943),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_101),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_2993),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_4234),
.Y(n_5903)
);

CKINVDCx5p33_ASAP7_75t_R g5904 ( 
.A(n_1880),
.Y(n_5904)
);

CKINVDCx5p33_ASAP7_75t_R g5905 ( 
.A(n_3735),
.Y(n_5905)
);

CKINVDCx5p33_ASAP7_75t_R g5906 ( 
.A(n_1600),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_4207),
.Y(n_5907)
);

CKINVDCx5p33_ASAP7_75t_R g5908 ( 
.A(n_2460),
.Y(n_5908)
);

CKINVDCx5p33_ASAP7_75t_R g5909 ( 
.A(n_4095),
.Y(n_5909)
);

CKINVDCx5p33_ASAP7_75t_R g5910 ( 
.A(n_1020),
.Y(n_5910)
);

INVx1_ASAP7_75t_L g5911 ( 
.A(n_2409),
.Y(n_5911)
);

CKINVDCx5p33_ASAP7_75t_R g5912 ( 
.A(n_2489),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_4524),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_540),
.Y(n_5914)
);

CKINVDCx14_ASAP7_75t_R g5915 ( 
.A(n_636),
.Y(n_5915)
);

CKINVDCx5p33_ASAP7_75t_R g5916 ( 
.A(n_4522),
.Y(n_5916)
);

CKINVDCx5p33_ASAP7_75t_R g5917 ( 
.A(n_2316),
.Y(n_5917)
);

CKINVDCx5p33_ASAP7_75t_R g5918 ( 
.A(n_1824),
.Y(n_5918)
);

CKINVDCx5p33_ASAP7_75t_R g5919 ( 
.A(n_944),
.Y(n_5919)
);

CKINVDCx20_ASAP7_75t_R g5920 ( 
.A(n_4581),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_2178),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_4507),
.Y(n_5922)
);

CKINVDCx5p33_ASAP7_75t_R g5923 ( 
.A(n_4417),
.Y(n_5923)
);

BUFx6f_ASAP7_75t_L g5924 ( 
.A(n_2593),
.Y(n_5924)
);

CKINVDCx5p33_ASAP7_75t_R g5925 ( 
.A(n_2784),
.Y(n_5925)
);

CKINVDCx5p33_ASAP7_75t_R g5926 ( 
.A(n_1585),
.Y(n_5926)
);

CKINVDCx5p33_ASAP7_75t_R g5927 ( 
.A(n_570),
.Y(n_5927)
);

CKINVDCx5p33_ASAP7_75t_R g5928 ( 
.A(n_894),
.Y(n_5928)
);

CKINVDCx5p33_ASAP7_75t_R g5929 ( 
.A(n_2091),
.Y(n_5929)
);

CKINVDCx5p33_ASAP7_75t_R g5930 ( 
.A(n_4657),
.Y(n_5930)
);

BUFx3_ASAP7_75t_L g5931 ( 
.A(n_1181),
.Y(n_5931)
);

INVx1_ASAP7_75t_SL g5932 ( 
.A(n_326),
.Y(n_5932)
);

CKINVDCx5p33_ASAP7_75t_R g5933 ( 
.A(n_1078),
.Y(n_5933)
);

BUFx10_ASAP7_75t_L g5934 ( 
.A(n_3845),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_2979),
.Y(n_5935)
);

BUFx5_ASAP7_75t_L g5936 ( 
.A(n_824),
.Y(n_5936)
);

INVx2_ASAP7_75t_L g5937 ( 
.A(n_1888),
.Y(n_5937)
);

BUFx6f_ASAP7_75t_L g5938 ( 
.A(n_1142),
.Y(n_5938)
);

CKINVDCx5p33_ASAP7_75t_R g5939 ( 
.A(n_4518),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_4406),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_4425),
.Y(n_5941)
);

BUFx3_ASAP7_75t_L g5942 ( 
.A(n_386),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_1526),
.Y(n_5943)
);

CKINVDCx5p33_ASAP7_75t_R g5944 ( 
.A(n_3004),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_4392),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_4004),
.Y(n_5946)
);

CKINVDCx5p33_ASAP7_75t_R g5947 ( 
.A(n_207),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_4489),
.Y(n_5948)
);

BUFx3_ASAP7_75t_L g5949 ( 
.A(n_1667),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_1514),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_4458),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_4551),
.Y(n_5952)
);

BUFx6f_ASAP7_75t_L g5953 ( 
.A(n_2540),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_1752),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_2938),
.Y(n_5955)
);

CKINVDCx5p33_ASAP7_75t_R g5956 ( 
.A(n_1249),
.Y(n_5956)
);

CKINVDCx5p33_ASAP7_75t_R g5957 ( 
.A(n_3135),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_4467),
.Y(n_5958)
);

CKINVDCx5p33_ASAP7_75t_R g5959 ( 
.A(n_34),
.Y(n_5959)
);

CKINVDCx5p33_ASAP7_75t_R g5960 ( 
.A(n_3490),
.Y(n_5960)
);

CKINVDCx5p33_ASAP7_75t_R g5961 ( 
.A(n_4220),
.Y(n_5961)
);

CKINVDCx5p33_ASAP7_75t_R g5962 ( 
.A(n_4459),
.Y(n_5962)
);

BUFx10_ASAP7_75t_L g5963 ( 
.A(n_783),
.Y(n_5963)
);

CKINVDCx5p33_ASAP7_75t_R g5964 ( 
.A(n_2770),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_120),
.Y(n_5965)
);

BUFx6f_ASAP7_75t_L g5966 ( 
.A(n_1460),
.Y(n_5966)
);

CKINVDCx16_ASAP7_75t_R g5967 ( 
.A(n_1679),
.Y(n_5967)
);

CKINVDCx5p33_ASAP7_75t_R g5968 ( 
.A(n_4455),
.Y(n_5968)
);

CKINVDCx5p33_ASAP7_75t_R g5969 ( 
.A(n_4541),
.Y(n_5969)
);

CKINVDCx20_ASAP7_75t_R g5970 ( 
.A(n_2094),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_729),
.Y(n_5971)
);

CKINVDCx5p33_ASAP7_75t_R g5972 ( 
.A(n_1819),
.Y(n_5972)
);

CKINVDCx5p33_ASAP7_75t_R g5973 ( 
.A(n_4379),
.Y(n_5973)
);

CKINVDCx5p33_ASAP7_75t_R g5974 ( 
.A(n_1106),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_973),
.Y(n_5975)
);

CKINVDCx5p33_ASAP7_75t_R g5976 ( 
.A(n_3818),
.Y(n_5976)
);

CKINVDCx5p33_ASAP7_75t_R g5977 ( 
.A(n_3734),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_784),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_1516),
.Y(n_5979)
);

BUFx6f_ASAP7_75t_L g5980 ( 
.A(n_4104),
.Y(n_5980)
);

BUFx10_ASAP7_75t_L g5981 ( 
.A(n_4516),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_4360),
.Y(n_5982)
);

CKINVDCx5p33_ASAP7_75t_R g5983 ( 
.A(n_3302),
.Y(n_5983)
);

CKINVDCx5p33_ASAP7_75t_R g5984 ( 
.A(n_653),
.Y(n_5984)
);

CKINVDCx20_ASAP7_75t_R g5985 ( 
.A(n_2375),
.Y(n_5985)
);

CKINVDCx5p33_ASAP7_75t_R g5986 ( 
.A(n_2628),
.Y(n_5986)
);

CKINVDCx5p33_ASAP7_75t_R g5987 ( 
.A(n_1254),
.Y(n_5987)
);

CKINVDCx5p33_ASAP7_75t_R g5988 ( 
.A(n_1498),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_192),
.Y(n_5989)
);

CKINVDCx5p33_ASAP7_75t_R g5990 ( 
.A(n_2343),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_1004),
.Y(n_5991)
);

INVx2_ASAP7_75t_SL g5992 ( 
.A(n_3492),
.Y(n_5992)
);

CKINVDCx5p33_ASAP7_75t_R g5993 ( 
.A(n_2557),
.Y(n_5993)
);

CKINVDCx5p33_ASAP7_75t_R g5994 ( 
.A(n_4072),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_1512),
.Y(n_5995)
);

CKINVDCx5p33_ASAP7_75t_R g5996 ( 
.A(n_2224),
.Y(n_5996)
);

CKINVDCx20_ASAP7_75t_R g5997 ( 
.A(n_3044),
.Y(n_5997)
);

CKINVDCx20_ASAP7_75t_R g5998 ( 
.A(n_4497),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_2726),
.Y(n_5999)
);

CKINVDCx20_ASAP7_75t_R g6000 ( 
.A(n_4017),
.Y(n_6000)
);

CKINVDCx5p33_ASAP7_75t_R g6001 ( 
.A(n_4081),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_3918),
.Y(n_6002)
);

CKINVDCx5p33_ASAP7_75t_R g6003 ( 
.A(n_3998),
.Y(n_6003)
);

CKINVDCx20_ASAP7_75t_R g6004 ( 
.A(n_4521),
.Y(n_6004)
);

CKINVDCx20_ASAP7_75t_R g6005 ( 
.A(n_2335),
.Y(n_6005)
);

CKINVDCx16_ASAP7_75t_R g6006 ( 
.A(n_4476),
.Y(n_6006)
);

INVx2_ASAP7_75t_L g6007 ( 
.A(n_1054),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_2257),
.Y(n_6008)
);

CKINVDCx5p33_ASAP7_75t_R g6009 ( 
.A(n_462),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_3788),
.Y(n_6010)
);

CKINVDCx5p33_ASAP7_75t_R g6011 ( 
.A(n_4418),
.Y(n_6011)
);

CKINVDCx5p33_ASAP7_75t_R g6012 ( 
.A(n_2990),
.Y(n_6012)
);

CKINVDCx5p33_ASAP7_75t_R g6013 ( 
.A(n_2599),
.Y(n_6013)
);

CKINVDCx5p33_ASAP7_75t_R g6014 ( 
.A(n_662),
.Y(n_6014)
);

CKINVDCx5p33_ASAP7_75t_R g6015 ( 
.A(n_4490),
.Y(n_6015)
);

CKINVDCx5p33_ASAP7_75t_R g6016 ( 
.A(n_928),
.Y(n_6016)
);

BUFx10_ASAP7_75t_L g6017 ( 
.A(n_2787),
.Y(n_6017)
);

BUFx8_ASAP7_75t_SL g6018 ( 
.A(n_1903),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_3663),
.Y(n_6019)
);

CKINVDCx5p33_ASAP7_75t_R g6020 ( 
.A(n_2911),
.Y(n_6020)
);

BUFx5_ASAP7_75t_L g6021 ( 
.A(n_4373),
.Y(n_6021)
);

CKINVDCx5p33_ASAP7_75t_R g6022 ( 
.A(n_546),
.Y(n_6022)
);

CKINVDCx5p33_ASAP7_75t_R g6023 ( 
.A(n_1968),
.Y(n_6023)
);

CKINVDCx5p33_ASAP7_75t_R g6024 ( 
.A(n_2840),
.Y(n_6024)
);

CKINVDCx14_ASAP7_75t_R g6025 ( 
.A(n_273),
.Y(n_6025)
);

INVx1_ASAP7_75t_SL g6026 ( 
.A(n_4530),
.Y(n_6026)
);

CKINVDCx5p33_ASAP7_75t_R g6027 ( 
.A(n_153),
.Y(n_6027)
);

INVx3_ASAP7_75t_L g6028 ( 
.A(n_3783),
.Y(n_6028)
);

CKINVDCx5p33_ASAP7_75t_R g6029 ( 
.A(n_3383),
.Y(n_6029)
);

CKINVDCx5p33_ASAP7_75t_R g6030 ( 
.A(n_1518),
.Y(n_6030)
);

INVx2_ASAP7_75t_L g6031 ( 
.A(n_3790),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_4474),
.Y(n_6032)
);

CKINVDCx5p33_ASAP7_75t_R g6033 ( 
.A(n_3877),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_3524),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_4432),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5127),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_72),
.Y(n_6037)
);

BUFx10_ASAP7_75t_L g6038 ( 
.A(n_1153),
.Y(n_6038)
);

CKINVDCx20_ASAP7_75t_R g6039 ( 
.A(n_2726),
.Y(n_6039)
);

CKINVDCx5p33_ASAP7_75t_R g6040 ( 
.A(n_1387),
.Y(n_6040)
);

INVx2_ASAP7_75t_SL g6041 ( 
.A(n_3170),
.Y(n_6041)
);

CKINVDCx20_ASAP7_75t_R g6042 ( 
.A(n_126),
.Y(n_6042)
);

CKINVDCx5p33_ASAP7_75t_R g6043 ( 
.A(n_2022),
.Y(n_6043)
);

CKINVDCx5p33_ASAP7_75t_R g6044 ( 
.A(n_3552),
.Y(n_6044)
);

BUFx5_ASAP7_75t_L g6045 ( 
.A(n_4342),
.Y(n_6045)
);

CKINVDCx5p33_ASAP7_75t_R g6046 ( 
.A(n_4064),
.Y(n_6046)
);

BUFx6f_ASAP7_75t_L g6047 ( 
.A(n_4514),
.Y(n_6047)
);

CKINVDCx20_ASAP7_75t_R g6048 ( 
.A(n_4784),
.Y(n_6048)
);

INVx2_ASAP7_75t_SL g6049 ( 
.A(n_3984),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_635),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_3034),
.Y(n_6051)
);

CKINVDCx16_ASAP7_75t_R g6052 ( 
.A(n_128),
.Y(n_6052)
);

CKINVDCx20_ASAP7_75t_R g6053 ( 
.A(n_4027),
.Y(n_6053)
);

CKINVDCx5p33_ASAP7_75t_R g6054 ( 
.A(n_4977),
.Y(n_6054)
);

CKINVDCx5p33_ASAP7_75t_R g6055 ( 
.A(n_3889),
.Y(n_6055)
);

CKINVDCx20_ASAP7_75t_R g6056 ( 
.A(n_2062),
.Y(n_6056)
);

CKINVDCx5p33_ASAP7_75t_R g6057 ( 
.A(n_172),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_3685),
.Y(n_6058)
);

CKINVDCx5p33_ASAP7_75t_R g6059 ( 
.A(n_3279),
.Y(n_6059)
);

BUFx6f_ASAP7_75t_L g6060 ( 
.A(n_1497),
.Y(n_6060)
);

CKINVDCx5p33_ASAP7_75t_R g6061 ( 
.A(n_2025),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_4411),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_3759),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_671),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_4524),
.Y(n_6065)
);

CKINVDCx20_ASAP7_75t_R g6066 ( 
.A(n_4506),
.Y(n_6066)
);

CKINVDCx20_ASAP7_75t_R g6067 ( 
.A(n_4270),
.Y(n_6067)
);

CKINVDCx5p33_ASAP7_75t_R g6068 ( 
.A(n_451),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_113),
.Y(n_6069)
);

CKINVDCx5p33_ASAP7_75t_R g6070 ( 
.A(n_44),
.Y(n_6070)
);

CKINVDCx5p33_ASAP7_75t_R g6071 ( 
.A(n_3560),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_3160),
.Y(n_6072)
);

CKINVDCx5p33_ASAP7_75t_R g6073 ( 
.A(n_439),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_3403),
.Y(n_6074)
);

CKINVDCx5p33_ASAP7_75t_R g6075 ( 
.A(n_4525),
.Y(n_6075)
);

BUFx6f_ASAP7_75t_L g6076 ( 
.A(n_1941),
.Y(n_6076)
);

CKINVDCx5p33_ASAP7_75t_R g6077 ( 
.A(n_4311),
.Y(n_6077)
);

CKINVDCx5p33_ASAP7_75t_R g6078 ( 
.A(n_1248),
.Y(n_6078)
);

CKINVDCx5p33_ASAP7_75t_R g6079 ( 
.A(n_3896),
.Y(n_6079)
);

CKINVDCx5p33_ASAP7_75t_R g6080 ( 
.A(n_4608),
.Y(n_6080)
);

INVxp67_ASAP7_75t_L g6081 ( 
.A(n_3258),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_4258),
.Y(n_6082)
);

CKINVDCx5p33_ASAP7_75t_R g6083 ( 
.A(n_4450),
.Y(n_6083)
);

CKINVDCx5p33_ASAP7_75t_R g6084 ( 
.A(n_3940),
.Y(n_6084)
);

CKINVDCx5p33_ASAP7_75t_R g6085 ( 
.A(n_4410),
.Y(n_6085)
);

CKINVDCx5p33_ASAP7_75t_R g6086 ( 
.A(n_4545),
.Y(n_6086)
);

BUFx8_ASAP7_75t_SL g6087 ( 
.A(n_1550),
.Y(n_6087)
);

CKINVDCx5p33_ASAP7_75t_R g6088 ( 
.A(n_2034),
.Y(n_6088)
);

CKINVDCx5p33_ASAP7_75t_R g6089 ( 
.A(n_4471),
.Y(n_6089)
);

CKINVDCx14_ASAP7_75t_R g6090 ( 
.A(n_4327),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_1571),
.Y(n_6091)
);

CKINVDCx5p33_ASAP7_75t_R g6092 ( 
.A(n_5061),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_93),
.Y(n_6093)
);

INVx3_ASAP7_75t_L g6094 ( 
.A(n_2847),
.Y(n_6094)
);

BUFx2_ASAP7_75t_SL g6095 ( 
.A(n_2064),
.Y(n_6095)
);

INVx3_ASAP7_75t_L g6096 ( 
.A(n_2834),
.Y(n_6096)
);

CKINVDCx5p33_ASAP7_75t_R g6097 ( 
.A(n_1396),
.Y(n_6097)
);

BUFx3_ASAP7_75t_L g6098 ( 
.A(n_952),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5092),
.Y(n_6099)
);

INVx1_ASAP7_75t_SL g6100 ( 
.A(n_3871),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_2021),
.Y(n_6101)
);

CKINVDCx5p33_ASAP7_75t_R g6102 ( 
.A(n_645),
.Y(n_6102)
);

BUFx10_ASAP7_75t_L g6103 ( 
.A(n_4700),
.Y(n_6103)
);

CKINVDCx5p33_ASAP7_75t_R g6104 ( 
.A(n_3595),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_2731),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_1592),
.Y(n_6106)
);

CKINVDCx5p33_ASAP7_75t_R g6107 ( 
.A(n_1994),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_2497),
.Y(n_6108)
);

BUFx10_ASAP7_75t_L g6109 ( 
.A(n_4368),
.Y(n_6109)
);

CKINVDCx5p33_ASAP7_75t_R g6110 ( 
.A(n_315),
.Y(n_6110)
);

BUFx3_ASAP7_75t_L g6111 ( 
.A(n_318),
.Y(n_6111)
);

CKINVDCx20_ASAP7_75t_R g6112 ( 
.A(n_36),
.Y(n_6112)
);

CKINVDCx5p33_ASAP7_75t_R g6113 ( 
.A(n_4951),
.Y(n_6113)
);

CKINVDCx5p33_ASAP7_75t_R g6114 ( 
.A(n_1746),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_2199),
.Y(n_6115)
);

CKINVDCx5p33_ASAP7_75t_R g6116 ( 
.A(n_4798),
.Y(n_6116)
);

CKINVDCx5p33_ASAP7_75t_R g6117 ( 
.A(n_2440),
.Y(n_6117)
);

CKINVDCx14_ASAP7_75t_R g6118 ( 
.A(n_2002),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_342),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_4559),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_3310),
.Y(n_6121)
);

INVx1_ASAP7_75t_SL g6122 ( 
.A(n_1716),
.Y(n_6122)
);

CKINVDCx5p33_ASAP7_75t_R g6123 ( 
.A(n_2876),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_715),
.Y(n_6124)
);

CKINVDCx5p33_ASAP7_75t_R g6125 ( 
.A(n_3771),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_1353),
.Y(n_6126)
);

CKINVDCx20_ASAP7_75t_R g6127 ( 
.A(n_4025),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_4423),
.Y(n_6128)
);

CKINVDCx5p33_ASAP7_75t_R g6129 ( 
.A(n_2413),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_1961),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_4927),
.Y(n_6131)
);

CKINVDCx5p33_ASAP7_75t_R g6132 ( 
.A(n_3677),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_3113),
.Y(n_6133)
);

CKINVDCx5p33_ASAP7_75t_R g6134 ( 
.A(n_3649),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_4023),
.Y(n_6135)
);

INVx2_ASAP7_75t_L g6136 ( 
.A(n_2432),
.Y(n_6136)
);

CKINVDCx5p33_ASAP7_75t_R g6137 ( 
.A(n_1757),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_2190),
.Y(n_6138)
);

CKINVDCx5p33_ASAP7_75t_R g6139 ( 
.A(n_1144),
.Y(n_6139)
);

CKINVDCx5p33_ASAP7_75t_R g6140 ( 
.A(n_2426),
.Y(n_6140)
);

BUFx10_ASAP7_75t_L g6141 ( 
.A(n_5078),
.Y(n_6141)
);

BUFx10_ASAP7_75t_L g6142 ( 
.A(n_3602),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_4157),
.Y(n_6143)
);

CKINVDCx5p33_ASAP7_75t_R g6144 ( 
.A(n_2167),
.Y(n_6144)
);

CKINVDCx5p33_ASAP7_75t_R g6145 ( 
.A(n_838),
.Y(n_6145)
);

CKINVDCx5p33_ASAP7_75t_R g6146 ( 
.A(n_3632),
.Y(n_6146)
);

CKINVDCx20_ASAP7_75t_R g6147 ( 
.A(n_4229),
.Y(n_6147)
);

CKINVDCx5p33_ASAP7_75t_R g6148 ( 
.A(n_4477),
.Y(n_6148)
);

CKINVDCx16_ASAP7_75t_R g6149 ( 
.A(n_105),
.Y(n_6149)
);

CKINVDCx14_ASAP7_75t_R g6150 ( 
.A(n_2708),
.Y(n_6150)
);

CKINVDCx5p33_ASAP7_75t_R g6151 ( 
.A(n_1954),
.Y(n_6151)
);

BUFx2_ASAP7_75t_L g6152 ( 
.A(n_4478),
.Y(n_6152)
);

CKINVDCx5p33_ASAP7_75t_R g6153 ( 
.A(n_4003),
.Y(n_6153)
);

CKINVDCx20_ASAP7_75t_R g6154 ( 
.A(n_4433),
.Y(n_6154)
);

CKINVDCx5p33_ASAP7_75t_R g6155 ( 
.A(n_3441),
.Y(n_6155)
);

CKINVDCx5p33_ASAP7_75t_R g6156 ( 
.A(n_4532),
.Y(n_6156)
);

CKINVDCx5p33_ASAP7_75t_R g6157 ( 
.A(n_744),
.Y(n_6157)
);

CKINVDCx5p33_ASAP7_75t_R g6158 ( 
.A(n_86),
.Y(n_6158)
);

CKINVDCx5p33_ASAP7_75t_R g6159 ( 
.A(n_4435),
.Y(n_6159)
);

INVx2_ASAP7_75t_L g6160 ( 
.A(n_3166),
.Y(n_6160)
);

CKINVDCx5p33_ASAP7_75t_R g6161 ( 
.A(n_942),
.Y(n_6161)
);

BUFx3_ASAP7_75t_L g6162 ( 
.A(n_4402),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_3301),
.Y(n_6163)
);

CKINVDCx5p33_ASAP7_75t_R g6164 ( 
.A(n_689),
.Y(n_6164)
);

CKINVDCx5p33_ASAP7_75t_R g6165 ( 
.A(n_4589),
.Y(n_6165)
);

INVx1_ASAP7_75t_SL g6166 ( 
.A(n_5160),
.Y(n_6166)
);

HB1xp67_ASAP7_75t_L g6167 ( 
.A(n_2916),
.Y(n_6167)
);

INVx1_ASAP7_75t_SL g6168 ( 
.A(n_4451),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_3093),
.Y(n_6169)
);

INVx2_ASAP7_75t_SL g6170 ( 
.A(n_36),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_3038),
.Y(n_6171)
);

CKINVDCx5p33_ASAP7_75t_R g6172 ( 
.A(n_3009),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_4400),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_1987),
.Y(n_6174)
);

CKINVDCx20_ASAP7_75t_R g6175 ( 
.A(n_851),
.Y(n_6175)
);

CKINVDCx5p33_ASAP7_75t_R g6176 ( 
.A(n_3779),
.Y(n_6176)
);

CKINVDCx5p33_ASAP7_75t_R g6177 ( 
.A(n_4698),
.Y(n_6177)
);

BUFx3_ASAP7_75t_L g6178 ( 
.A(n_4375),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_3805),
.Y(n_6179)
);

CKINVDCx5p33_ASAP7_75t_R g6180 ( 
.A(n_28),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_3697),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_1910),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_4473),
.Y(n_6183)
);

CKINVDCx5p33_ASAP7_75t_R g6184 ( 
.A(n_404),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_4503),
.Y(n_6185)
);

CKINVDCx5p33_ASAP7_75t_R g6186 ( 
.A(n_4712),
.Y(n_6186)
);

CKINVDCx5p33_ASAP7_75t_R g6187 ( 
.A(n_1168),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_4369),
.Y(n_6188)
);

CKINVDCx5p33_ASAP7_75t_R g6189 ( 
.A(n_1360),
.Y(n_6189)
);

CKINVDCx20_ASAP7_75t_R g6190 ( 
.A(n_4499),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_916),
.Y(n_6191)
);

INVx1_ASAP7_75t_SL g6192 ( 
.A(n_863),
.Y(n_6192)
);

CKINVDCx5p33_ASAP7_75t_R g6193 ( 
.A(n_4791),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_4495),
.Y(n_6194)
);

INVx1_ASAP7_75t_SL g6195 ( 
.A(n_3590),
.Y(n_6195)
);

CKINVDCx5p33_ASAP7_75t_R g6196 ( 
.A(n_3565),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_749),
.Y(n_6197)
);

CKINVDCx5p33_ASAP7_75t_R g6198 ( 
.A(n_4509),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_2546),
.Y(n_6199)
);

CKINVDCx5p33_ASAP7_75t_R g6200 ( 
.A(n_2161),
.Y(n_6200)
);

CKINVDCx5p33_ASAP7_75t_R g6201 ( 
.A(n_813),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_980),
.Y(n_6202)
);

CKINVDCx14_ASAP7_75t_R g6203 ( 
.A(n_4380),
.Y(n_6203)
);

CKINVDCx5p33_ASAP7_75t_R g6204 ( 
.A(n_4285),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_2496),
.Y(n_6205)
);

CKINVDCx5p33_ASAP7_75t_R g6206 ( 
.A(n_2770),
.Y(n_6206)
);

CKINVDCx5p33_ASAP7_75t_R g6207 ( 
.A(n_2637),
.Y(n_6207)
);

CKINVDCx5p33_ASAP7_75t_R g6208 ( 
.A(n_1862),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_4552),
.Y(n_6209)
);

CKINVDCx5p33_ASAP7_75t_R g6210 ( 
.A(n_1133),
.Y(n_6210)
);

BUFx3_ASAP7_75t_L g6211 ( 
.A(n_665),
.Y(n_6211)
);

CKINVDCx5p33_ASAP7_75t_R g6212 ( 
.A(n_2222),
.Y(n_6212)
);

CKINVDCx5p33_ASAP7_75t_R g6213 ( 
.A(n_2150),
.Y(n_6213)
);

CKINVDCx5p33_ASAP7_75t_R g6214 ( 
.A(n_3435),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_4902),
.Y(n_6215)
);

CKINVDCx5p33_ASAP7_75t_R g6216 ( 
.A(n_3368),
.Y(n_6216)
);

INVx2_ASAP7_75t_SL g6217 ( 
.A(n_4539),
.Y(n_6217)
);

CKINVDCx20_ASAP7_75t_R g6218 ( 
.A(n_2724),
.Y(n_6218)
);

BUFx6f_ASAP7_75t_L g6219 ( 
.A(n_2799),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_3462),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_5089),
.Y(n_6221)
);

CKINVDCx5p33_ASAP7_75t_R g6222 ( 
.A(n_3894),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_2410),
.Y(n_6223)
);

INVx1_ASAP7_75t_SL g6224 ( 
.A(n_4321),
.Y(n_6224)
);

CKINVDCx5p33_ASAP7_75t_R g6225 ( 
.A(n_1594),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_1722),
.Y(n_6226)
);

CKINVDCx5p33_ASAP7_75t_R g6227 ( 
.A(n_4595),
.Y(n_6227)
);

CKINVDCx5p33_ASAP7_75t_R g6228 ( 
.A(n_5006),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_2170),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_4389),
.Y(n_6230)
);

CKINVDCx5p33_ASAP7_75t_R g6231 ( 
.A(n_1653),
.Y(n_6231)
);

CKINVDCx5p33_ASAP7_75t_R g6232 ( 
.A(n_2689),
.Y(n_6232)
);

CKINVDCx5p33_ASAP7_75t_R g6233 ( 
.A(n_1481),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_4474),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_3176),
.Y(n_6235)
);

CKINVDCx5p33_ASAP7_75t_R g6236 ( 
.A(n_2410),
.Y(n_6236)
);

CKINVDCx5p33_ASAP7_75t_R g6237 ( 
.A(n_4507),
.Y(n_6237)
);

CKINVDCx5p33_ASAP7_75t_R g6238 ( 
.A(n_2801),
.Y(n_6238)
);

BUFx3_ASAP7_75t_L g6239 ( 
.A(n_2631),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_4320),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_2063),
.Y(n_6241)
);

CKINVDCx5p33_ASAP7_75t_R g6242 ( 
.A(n_1976),
.Y(n_6242)
);

BUFx2_ASAP7_75t_L g6243 ( 
.A(n_3821),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_305),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_3725),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_1472),
.Y(n_6246)
);

CKINVDCx5p33_ASAP7_75t_R g6247 ( 
.A(n_3999),
.Y(n_6247)
);

CKINVDCx5p33_ASAP7_75t_R g6248 ( 
.A(n_3398),
.Y(n_6248)
);

CKINVDCx5p33_ASAP7_75t_R g6249 ( 
.A(n_691),
.Y(n_6249)
);

CKINVDCx5p33_ASAP7_75t_R g6250 ( 
.A(n_3025),
.Y(n_6250)
);

INVx1_ASAP7_75t_SL g6251 ( 
.A(n_4957),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_4408),
.Y(n_6252)
);

CKINVDCx5p33_ASAP7_75t_R g6253 ( 
.A(n_3931),
.Y(n_6253)
);

CKINVDCx5p33_ASAP7_75t_R g6254 ( 
.A(n_4941),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_3881),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_4354),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_4174),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_1448),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_4268),
.Y(n_6259)
);

CKINVDCx5p33_ASAP7_75t_R g6260 ( 
.A(n_542),
.Y(n_6260)
);

HB1xp67_ASAP7_75t_L g6261 ( 
.A(n_1353),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_4445),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_4350),
.Y(n_6263)
);

CKINVDCx5p33_ASAP7_75t_R g6264 ( 
.A(n_4043),
.Y(n_6264)
);

CKINVDCx20_ASAP7_75t_R g6265 ( 
.A(n_4897),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_885),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_2102),
.Y(n_6267)
);

CKINVDCx5p33_ASAP7_75t_R g6268 ( 
.A(n_704),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_3020),
.Y(n_6269)
);

CKINVDCx5p33_ASAP7_75t_R g6270 ( 
.A(n_4500),
.Y(n_6270)
);

CKINVDCx5p33_ASAP7_75t_R g6271 ( 
.A(n_168),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_1787),
.Y(n_6272)
);

CKINVDCx5p33_ASAP7_75t_R g6273 ( 
.A(n_4655),
.Y(n_6273)
);

CKINVDCx5p33_ASAP7_75t_R g6274 ( 
.A(n_617),
.Y(n_6274)
);

CKINVDCx5p33_ASAP7_75t_R g6275 ( 
.A(n_3156),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_2736),
.Y(n_6276)
);

BUFx10_ASAP7_75t_L g6277 ( 
.A(n_4505),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_3395),
.Y(n_6278)
);

CKINVDCx5p33_ASAP7_75t_R g6279 ( 
.A(n_2394),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_4435),
.Y(n_6280)
);

BUFx8_ASAP7_75t_SL g6281 ( 
.A(n_2709),
.Y(n_6281)
);

BUFx3_ASAP7_75t_L g6282 ( 
.A(n_3641),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_4968),
.Y(n_6283)
);

CKINVDCx5p33_ASAP7_75t_R g6284 ( 
.A(n_1476),
.Y(n_6284)
);

CKINVDCx20_ASAP7_75t_R g6285 ( 
.A(n_4367),
.Y(n_6285)
);

CKINVDCx20_ASAP7_75t_R g6286 ( 
.A(n_179),
.Y(n_6286)
);

INVx1_ASAP7_75t_SL g6287 ( 
.A(n_4420),
.Y(n_6287)
);

CKINVDCx5p33_ASAP7_75t_R g6288 ( 
.A(n_2318),
.Y(n_6288)
);

CKINVDCx5p33_ASAP7_75t_R g6289 ( 
.A(n_2271),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_1108),
.Y(n_6290)
);

INVx2_ASAP7_75t_L g6291 ( 
.A(n_589),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_4230),
.Y(n_6292)
);

BUFx10_ASAP7_75t_L g6293 ( 
.A(n_1639),
.Y(n_6293)
);

CKINVDCx16_ASAP7_75t_R g6294 ( 
.A(n_57),
.Y(n_6294)
);

CKINVDCx5p33_ASAP7_75t_R g6295 ( 
.A(n_3372),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_3703),
.Y(n_6296)
);

CKINVDCx5p33_ASAP7_75t_R g6297 ( 
.A(n_973),
.Y(n_6297)
);

CKINVDCx5p33_ASAP7_75t_R g6298 ( 
.A(n_524),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_915),
.Y(n_6299)
);

CKINVDCx5p33_ASAP7_75t_R g6300 ( 
.A(n_4256),
.Y(n_6300)
);

CKINVDCx5p33_ASAP7_75t_R g6301 ( 
.A(n_4830),
.Y(n_6301)
);

CKINVDCx5p33_ASAP7_75t_R g6302 ( 
.A(n_1215),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_4442),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_3056),
.Y(n_6304)
);

CKINVDCx5p33_ASAP7_75t_R g6305 ( 
.A(n_595),
.Y(n_6305)
);

CKINVDCx5p33_ASAP7_75t_R g6306 ( 
.A(n_2697),
.Y(n_6306)
);

BUFx10_ASAP7_75t_L g6307 ( 
.A(n_5141),
.Y(n_6307)
);

CKINVDCx5p33_ASAP7_75t_R g6308 ( 
.A(n_1253),
.Y(n_6308)
);

CKINVDCx5p33_ASAP7_75t_R g6309 ( 
.A(n_708),
.Y(n_6309)
);

CKINVDCx14_ASAP7_75t_R g6310 ( 
.A(n_1301),
.Y(n_6310)
);

BUFx3_ASAP7_75t_L g6311 ( 
.A(n_1930),
.Y(n_6311)
);

CKINVDCx5p33_ASAP7_75t_R g6312 ( 
.A(n_30),
.Y(n_6312)
);

CKINVDCx5p33_ASAP7_75t_R g6313 ( 
.A(n_3384),
.Y(n_6313)
);

CKINVDCx5p33_ASAP7_75t_R g6314 ( 
.A(n_2454),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_3481),
.Y(n_6315)
);

CKINVDCx5p33_ASAP7_75t_R g6316 ( 
.A(n_2062),
.Y(n_6316)
);

CKINVDCx5p33_ASAP7_75t_R g6317 ( 
.A(n_4391),
.Y(n_6317)
);

BUFx3_ASAP7_75t_L g6318 ( 
.A(n_2758),
.Y(n_6318)
);

INVx2_ASAP7_75t_L g6319 ( 
.A(n_3984),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_4971),
.Y(n_6320)
);

BUFx5_ASAP7_75t_L g6321 ( 
.A(n_2222),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_4883),
.Y(n_6322)
);

CKINVDCx5p33_ASAP7_75t_R g6323 ( 
.A(n_4377),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_1299),
.Y(n_6324)
);

INVx2_ASAP7_75t_SL g6325 ( 
.A(n_696),
.Y(n_6325)
);

CKINVDCx5p33_ASAP7_75t_R g6326 ( 
.A(n_7),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_1675),
.Y(n_6327)
);

CKINVDCx5p33_ASAP7_75t_R g6328 ( 
.A(n_1022),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_3491),
.Y(n_6329)
);

BUFx3_ASAP7_75t_L g6330 ( 
.A(n_2710),
.Y(n_6330)
);

CKINVDCx5p33_ASAP7_75t_R g6331 ( 
.A(n_4708),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_2558),
.Y(n_6332)
);

CKINVDCx5p33_ASAP7_75t_R g6333 ( 
.A(n_86),
.Y(n_6333)
);

CKINVDCx5p33_ASAP7_75t_R g6334 ( 
.A(n_779),
.Y(n_6334)
);

CKINVDCx5p33_ASAP7_75t_R g6335 ( 
.A(n_4136),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_595),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_1823),
.Y(n_6337)
);

CKINVDCx16_ASAP7_75t_R g6338 ( 
.A(n_4806),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_4397),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_3372),
.Y(n_6340)
);

CKINVDCx5p33_ASAP7_75t_R g6341 ( 
.A(n_4527),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_3822),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_4535),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_972),
.Y(n_6344)
);

INVx1_ASAP7_75t_SL g6345 ( 
.A(n_128),
.Y(n_6345)
);

CKINVDCx5p33_ASAP7_75t_R g6346 ( 
.A(n_3480),
.Y(n_6346)
);

CKINVDCx5p33_ASAP7_75t_R g6347 ( 
.A(n_3970),
.Y(n_6347)
);

CKINVDCx5p33_ASAP7_75t_R g6348 ( 
.A(n_4214),
.Y(n_6348)
);

CKINVDCx5p33_ASAP7_75t_R g6349 ( 
.A(n_3241),
.Y(n_6349)
);

BUFx6f_ASAP7_75t_L g6350 ( 
.A(n_484),
.Y(n_6350)
);

CKINVDCx5p33_ASAP7_75t_R g6351 ( 
.A(n_3402),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_1964),
.Y(n_6352)
);

CKINVDCx5p33_ASAP7_75t_R g6353 ( 
.A(n_1321),
.Y(n_6353)
);

CKINVDCx5p33_ASAP7_75t_R g6354 ( 
.A(n_1011),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_4416),
.Y(n_6355)
);

CKINVDCx5p33_ASAP7_75t_R g6356 ( 
.A(n_2851),
.Y(n_6356)
);

CKINVDCx5p33_ASAP7_75t_R g6357 ( 
.A(n_5073),
.Y(n_6357)
);

CKINVDCx5p33_ASAP7_75t_R g6358 ( 
.A(n_3678),
.Y(n_6358)
);

BUFx10_ASAP7_75t_L g6359 ( 
.A(n_3896),
.Y(n_6359)
);

BUFx6f_ASAP7_75t_L g6360 ( 
.A(n_5097),
.Y(n_6360)
);

CKINVDCx5p33_ASAP7_75t_R g6361 ( 
.A(n_4953),
.Y(n_6361)
);

INVx1_ASAP7_75t_SL g6362 ( 
.A(n_5003),
.Y(n_6362)
);

CKINVDCx5p33_ASAP7_75t_R g6363 ( 
.A(n_1427),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_4463),
.Y(n_6364)
);

CKINVDCx20_ASAP7_75t_R g6365 ( 
.A(n_4419),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_2238),
.Y(n_6366)
);

CKINVDCx5p33_ASAP7_75t_R g6367 ( 
.A(n_3113),
.Y(n_6367)
);

CKINVDCx5p33_ASAP7_75t_R g6368 ( 
.A(n_4547),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_1213),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_67),
.Y(n_6370)
);

CKINVDCx5p33_ASAP7_75t_R g6371 ( 
.A(n_2092),
.Y(n_6371)
);

CKINVDCx5p33_ASAP7_75t_R g6372 ( 
.A(n_5029),
.Y(n_6372)
);

INVx2_ASAP7_75t_SL g6373 ( 
.A(n_1297),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_2590),
.Y(n_6374)
);

CKINVDCx5p33_ASAP7_75t_R g6375 ( 
.A(n_3882),
.Y(n_6375)
);

CKINVDCx5p33_ASAP7_75t_R g6376 ( 
.A(n_445),
.Y(n_6376)
);

CKINVDCx5p33_ASAP7_75t_R g6377 ( 
.A(n_2764),
.Y(n_6377)
);

CKINVDCx5p33_ASAP7_75t_R g6378 ( 
.A(n_803),
.Y(n_6378)
);

CKINVDCx5p33_ASAP7_75t_R g6379 ( 
.A(n_1225),
.Y(n_6379)
);

CKINVDCx20_ASAP7_75t_R g6380 ( 
.A(n_1470),
.Y(n_6380)
);

BUFx6f_ASAP7_75t_L g6381 ( 
.A(n_4519),
.Y(n_6381)
);

CKINVDCx20_ASAP7_75t_R g6382 ( 
.A(n_3893),
.Y(n_6382)
);

BUFx2_ASAP7_75t_L g6383 ( 
.A(n_875),
.Y(n_6383)
);

CKINVDCx5p33_ASAP7_75t_R g6384 ( 
.A(n_470),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_4453),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_728),
.Y(n_6386)
);

CKINVDCx5p33_ASAP7_75t_R g6387 ( 
.A(n_2081),
.Y(n_6387)
);

CKINVDCx5p33_ASAP7_75t_R g6388 ( 
.A(n_1949),
.Y(n_6388)
);

CKINVDCx5p33_ASAP7_75t_R g6389 ( 
.A(n_3513),
.Y(n_6389)
);

CKINVDCx5p33_ASAP7_75t_R g6390 ( 
.A(n_60),
.Y(n_6390)
);

CKINVDCx5p33_ASAP7_75t_R g6391 ( 
.A(n_2757),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_3590),
.Y(n_6392)
);

CKINVDCx5p33_ASAP7_75t_R g6393 ( 
.A(n_291),
.Y(n_6393)
);

BUFx10_ASAP7_75t_L g6394 ( 
.A(n_4033),
.Y(n_6394)
);

CKINVDCx5p33_ASAP7_75t_R g6395 ( 
.A(n_4485),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_4701),
.Y(n_6396)
);

BUFx10_ASAP7_75t_L g6397 ( 
.A(n_2739),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_294),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_405),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_238),
.Y(n_6400)
);

BUFx2_ASAP7_75t_L g6401 ( 
.A(n_5121),
.Y(n_6401)
);

CKINVDCx5p33_ASAP7_75t_R g6402 ( 
.A(n_3340),
.Y(n_6402)
);

BUFx5_ASAP7_75t_L g6403 ( 
.A(n_4237),
.Y(n_6403)
);

CKINVDCx5p33_ASAP7_75t_R g6404 ( 
.A(n_4807),
.Y(n_6404)
);

CKINVDCx5p33_ASAP7_75t_R g6405 ( 
.A(n_1606),
.Y(n_6405)
);

CKINVDCx5p33_ASAP7_75t_R g6406 ( 
.A(n_4508),
.Y(n_6406)
);

CKINVDCx5p33_ASAP7_75t_R g6407 ( 
.A(n_4982),
.Y(n_6407)
);

CKINVDCx5p33_ASAP7_75t_R g6408 ( 
.A(n_73),
.Y(n_6408)
);

BUFx10_ASAP7_75t_L g6409 ( 
.A(n_4938),
.Y(n_6409)
);

CKINVDCx20_ASAP7_75t_R g6410 ( 
.A(n_2708),
.Y(n_6410)
);

CKINVDCx5p33_ASAP7_75t_R g6411 ( 
.A(n_4418),
.Y(n_6411)
);

CKINVDCx5p33_ASAP7_75t_R g6412 ( 
.A(n_3162),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_1235),
.Y(n_6413)
);

CKINVDCx5p33_ASAP7_75t_R g6414 ( 
.A(n_3983),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_3336),
.Y(n_6415)
);

CKINVDCx5p33_ASAP7_75t_R g6416 ( 
.A(n_2942),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_4172),
.Y(n_6417)
);

BUFx3_ASAP7_75t_L g6418 ( 
.A(n_2787),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_4102),
.Y(n_6419)
);

CKINVDCx5p33_ASAP7_75t_R g6420 ( 
.A(n_1444),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_368),
.Y(n_6421)
);

BUFx10_ASAP7_75t_L g6422 ( 
.A(n_281),
.Y(n_6422)
);

CKINVDCx5p33_ASAP7_75t_R g6423 ( 
.A(n_1518),
.Y(n_6423)
);

CKINVDCx16_ASAP7_75t_R g6424 ( 
.A(n_2844),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_4482),
.Y(n_6425)
);

CKINVDCx5p33_ASAP7_75t_R g6426 ( 
.A(n_572),
.Y(n_6426)
);

CKINVDCx5p33_ASAP7_75t_R g6427 ( 
.A(n_4448),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_3667),
.Y(n_6428)
);

CKINVDCx5p33_ASAP7_75t_R g6429 ( 
.A(n_649),
.Y(n_6429)
);

CKINVDCx5p33_ASAP7_75t_R g6430 ( 
.A(n_226),
.Y(n_6430)
);

CKINVDCx20_ASAP7_75t_R g6431 ( 
.A(n_2331),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_5016),
.Y(n_6432)
);

CKINVDCx5p33_ASAP7_75t_R g6433 ( 
.A(n_2315),
.Y(n_6433)
);

CKINVDCx20_ASAP7_75t_R g6434 ( 
.A(n_2606),
.Y(n_6434)
);

BUFx10_ASAP7_75t_L g6435 ( 
.A(n_2106),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_1514),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_1428),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_3419),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_2763),
.Y(n_6439)
);

CKINVDCx5p33_ASAP7_75t_R g6440 ( 
.A(n_4394),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_2440),
.Y(n_6441)
);

CKINVDCx5p33_ASAP7_75t_R g6442 ( 
.A(n_817),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_1705),
.Y(n_6443)
);

CKINVDCx16_ASAP7_75t_R g6444 ( 
.A(n_4483),
.Y(n_6444)
);

CKINVDCx5p33_ASAP7_75t_R g6445 ( 
.A(n_309),
.Y(n_6445)
);

CKINVDCx5p33_ASAP7_75t_R g6446 ( 
.A(n_501),
.Y(n_6446)
);

CKINVDCx5p33_ASAP7_75t_R g6447 ( 
.A(n_757),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_4253),
.Y(n_6448)
);

CKINVDCx5p33_ASAP7_75t_R g6449 ( 
.A(n_580),
.Y(n_6449)
);

CKINVDCx5p33_ASAP7_75t_R g6450 ( 
.A(n_4793),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_1874),
.Y(n_6451)
);

CKINVDCx5p33_ASAP7_75t_R g6452 ( 
.A(n_597),
.Y(n_6452)
);

CKINVDCx5p33_ASAP7_75t_R g6453 ( 
.A(n_4581),
.Y(n_6453)
);

CKINVDCx5p33_ASAP7_75t_R g6454 ( 
.A(n_2943),
.Y(n_6454)
);

CKINVDCx5p33_ASAP7_75t_R g6455 ( 
.A(n_3200),
.Y(n_6455)
);

CKINVDCx5p33_ASAP7_75t_R g6456 ( 
.A(n_698),
.Y(n_6456)
);

BUFx3_ASAP7_75t_L g6457 ( 
.A(n_1722),
.Y(n_6457)
);

CKINVDCx5p33_ASAP7_75t_R g6458 ( 
.A(n_5035),
.Y(n_6458)
);

CKINVDCx5p33_ASAP7_75t_R g6459 ( 
.A(n_2122),
.Y(n_6459)
);

CKINVDCx5p33_ASAP7_75t_R g6460 ( 
.A(n_5091),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_3871),
.Y(n_6461)
);

INVx1_ASAP7_75t_SL g6462 ( 
.A(n_1543),
.Y(n_6462)
);

CKINVDCx5p33_ASAP7_75t_R g6463 ( 
.A(n_1957),
.Y(n_6463)
);

CKINVDCx5p33_ASAP7_75t_R g6464 ( 
.A(n_516),
.Y(n_6464)
);

CKINVDCx5p33_ASAP7_75t_R g6465 ( 
.A(n_3225),
.Y(n_6465)
);

CKINVDCx16_ASAP7_75t_R g6466 ( 
.A(n_4512),
.Y(n_6466)
);

INVx1_ASAP7_75t_SL g6467 ( 
.A(n_3099),
.Y(n_6467)
);

HB1xp67_ASAP7_75t_L g6468 ( 
.A(n_1547),
.Y(n_6468)
);

CKINVDCx20_ASAP7_75t_R g6469 ( 
.A(n_470),
.Y(n_6469)
);

CKINVDCx5p33_ASAP7_75t_R g6470 ( 
.A(n_4050),
.Y(n_6470)
);

CKINVDCx5p33_ASAP7_75t_R g6471 ( 
.A(n_4739),
.Y(n_6471)
);

CKINVDCx5p33_ASAP7_75t_R g6472 ( 
.A(n_399),
.Y(n_6472)
);

CKINVDCx5p33_ASAP7_75t_R g6473 ( 
.A(n_1188),
.Y(n_6473)
);

CKINVDCx5p33_ASAP7_75t_R g6474 ( 
.A(n_3105),
.Y(n_6474)
);

CKINVDCx5p33_ASAP7_75t_R g6475 ( 
.A(n_2244),
.Y(n_6475)
);

CKINVDCx5p33_ASAP7_75t_R g6476 ( 
.A(n_2530),
.Y(n_6476)
);

CKINVDCx5p33_ASAP7_75t_R g6477 ( 
.A(n_4235),
.Y(n_6477)
);

BUFx6f_ASAP7_75t_L g6478 ( 
.A(n_4419),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_4504),
.Y(n_6479)
);

BUFx3_ASAP7_75t_L g6480 ( 
.A(n_4528),
.Y(n_6480)
);

CKINVDCx5p33_ASAP7_75t_R g6481 ( 
.A(n_1978),
.Y(n_6481)
);

BUFx5_ASAP7_75t_L g6482 ( 
.A(n_3449),
.Y(n_6482)
);

CKINVDCx20_ASAP7_75t_R g6483 ( 
.A(n_2959),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_719),
.Y(n_6484)
);

CKINVDCx5p33_ASAP7_75t_R g6485 ( 
.A(n_1784),
.Y(n_6485)
);

CKINVDCx5p33_ASAP7_75t_R g6486 ( 
.A(n_2213),
.Y(n_6486)
);

CKINVDCx5p33_ASAP7_75t_R g6487 ( 
.A(n_1455),
.Y(n_6487)
);

CKINVDCx5p33_ASAP7_75t_R g6488 ( 
.A(n_4529),
.Y(n_6488)
);

INVx1_ASAP7_75t_SL g6489 ( 
.A(n_2650),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_4165),
.Y(n_6490)
);

BUFx2_ASAP7_75t_L g6491 ( 
.A(n_3702),
.Y(n_6491)
);

CKINVDCx5p33_ASAP7_75t_R g6492 ( 
.A(n_206),
.Y(n_6492)
);

CKINVDCx5p33_ASAP7_75t_R g6493 ( 
.A(n_4659),
.Y(n_6493)
);

BUFx6f_ASAP7_75t_L g6494 ( 
.A(n_4895),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_3558),
.Y(n_6495)
);

CKINVDCx20_ASAP7_75t_R g6496 ( 
.A(n_4536),
.Y(n_6496)
);

INVx1_ASAP7_75t_SL g6497 ( 
.A(n_2384),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_564),
.Y(n_6498)
);

CKINVDCx5p33_ASAP7_75t_R g6499 ( 
.A(n_1005),
.Y(n_6499)
);

CKINVDCx5p33_ASAP7_75t_R g6500 ( 
.A(n_4550),
.Y(n_6500)
);

CKINVDCx5p33_ASAP7_75t_R g6501 ( 
.A(n_977),
.Y(n_6501)
);

CKINVDCx5p33_ASAP7_75t_R g6502 ( 
.A(n_1059),
.Y(n_6502)
);

BUFx6f_ASAP7_75t_L g6503 ( 
.A(n_2271),
.Y(n_6503)
);

CKINVDCx5p33_ASAP7_75t_R g6504 ( 
.A(n_4515),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_2873),
.Y(n_6505)
);

INVxp67_ASAP7_75t_L g6506 ( 
.A(n_3816),
.Y(n_6506)
);

CKINVDCx5p33_ASAP7_75t_R g6507 ( 
.A(n_1048),
.Y(n_6507)
);

CKINVDCx5p33_ASAP7_75t_R g6508 ( 
.A(n_4825),
.Y(n_6508)
);

CKINVDCx5p33_ASAP7_75t_R g6509 ( 
.A(n_4942),
.Y(n_6509)
);

CKINVDCx5p33_ASAP7_75t_R g6510 ( 
.A(n_2040),
.Y(n_6510)
);

CKINVDCx5p33_ASAP7_75t_R g6511 ( 
.A(n_229),
.Y(n_6511)
);

CKINVDCx5p33_ASAP7_75t_R g6512 ( 
.A(n_1367),
.Y(n_6512)
);

INVx1_ASAP7_75t_SL g6513 ( 
.A(n_2216),
.Y(n_6513)
);

CKINVDCx5p33_ASAP7_75t_R g6514 ( 
.A(n_1484),
.Y(n_6514)
);

CKINVDCx5p33_ASAP7_75t_R g6515 ( 
.A(n_4676),
.Y(n_6515)
);

CKINVDCx5p33_ASAP7_75t_R g6516 ( 
.A(n_4468),
.Y(n_6516)
);

CKINVDCx5p33_ASAP7_75t_R g6517 ( 
.A(n_27),
.Y(n_6517)
);

CKINVDCx5p33_ASAP7_75t_R g6518 ( 
.A(n_2509),
.Y(n_6518)
);

CKINVDCx5p33_ASAP7_75t_R g6519 ( 
.A(n_1356),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_2532),
.Y(n_6520)
);

BUFx3_ASAP7_75t_L g6521 ( 
.A(n_1865),
.Y(n_6521)
);

CKINVDCx5p33_ASAP7_75t_R g6522 ( 
.A(n_5060),
.Y(n_6522)
);

CKINVDCx5p33_ASAP7_75t_R g6523 ( 
.A(n_3112),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_1106),
.Y(n_6524)
);

CKINVDCx16_ASAP7_75t_R g6525 ( 
.A(n_304),
.Y(n_6525)
);

BUFx3_ASAP7_75t_L g6526 ( 
.A(n_1552),
.Y(n_6526)
);

BUFx2_ASAP7_75t_L g6527 ( 
.A(n_2282),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_5149),
.Y(n_6528)
);

INVx1_ASAP7_75t_SL g6529 ( 
.A(n_4393),
.Y(n_6529)
);

CKINVDCx5p33_ASAP7_75t_R g6530 ( 
.A(n_4446),
.Y(n_6530)
);

CKINVDCx5p33_ASAP7_75t_R g6531 ( 
.A(n_4409),
.Y(n_6531)
);

BUFx10_ASAP7_75t_L g6532 ( 
.A(n_766),
.Y(n_6532)
);

BUFx5_ASAP7_75t_L g6533 ( 
.A(n_4484),
.Y(n_6533)
);

HB1xp67_ASAP7_75t_L g6534 ( 
.A(n_2467),
.Y(n_6534)
);

BUFx3_ASAP7_75t_L g6535 ( 
.A(n_3431),
.Y(n_6535)
);

INVx2_ASAP7_75t_SL g6536 ( 
.A(n_315),
.Y(n_6536)
);

INVx1_ASAP7_75t_SL g6537 ( 
.A(n_4424),
.Y(n_6537)
);

CKINVDCx5p33_ASAP7_75t_R g6538 ( 
.A(n_1251),
.Y(n_6538)
);

CKINVDCx5p33_ASAP7_75t_R g6539 ( 
.A(n_4599),
.Y(n_6539)
);

CKINVDCx5p33_ASAP7_75t_R g6540 ( 
.A(n_4948),
.Y(n_6540)
);

CKINVDCx5p33_ASAP7_75t_R g6541 ( 
.A(n_4551),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_3044),
.Y(n_6542)
);

CKINVDCx5p33_ASAP7_75t_R g6543 ( 
.A(n_2649),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_3069),
.Y(n_6544)
);

CKINVDCx5p33_ASAP7_75t_R g6545 ( 
.A(n_3999),
.Y(n_6545)
);

CKINVDCx5p33_ASAP7_75t_R g6546 ( 
.A(n_2039),
.Y(n_6546)
);

BUFx3_ASAP7_75t_L g6547 ( 
.A(n_1253),
.Y(n_6547)
);

CKINVDCx5p33_ASAP7_75t_R g6548 ( 
.A(n_4702),
.Y(n_6548)
);

CKINVDCx20_ASAP7_75t_R g6549 ( 
.A(n_4829),
.Y(n_6549)
);

CKINVDCx5p33_ASAP7_75t_R g6550 ( 
.A(n_2692),
.Y(n_6550)
);

CKINVDCx5p33_ASAP7_75t_R g6551 ( 
.A(n_4751),
.Y(n_6551)
);

INVx2_ASAP7_75t_L g6552 ( 
.A(n_1552),
.Y(n_6552)
);

INVx1_ASAP7_75t_SL g6553 ( 
.A(n_3379),
.Y(n_6553)
);

CKINVDCx5p33_ASAP7_75t_R g6554 ( 
.A(n_3424),
.Y(n_6554)
);

INVx2_ASAP7_75t_L g6555 ( 
.A(n_4443),
.Y(n_6555)
);

BUFx3_ASAP7_75t_L g6556 ( 
.A(n_2446),
.Y(n_6556)
);

BUFx6f_ASAP7_75t_L g6557 ( 
.A(n_3228),
.Y(n_6557)
);

CKINVDCx5p33_ASAP7_75t_R g6558 ( 
.A(n_2389),
.Y(n_6558)
);

BUFx2_ASAP7_75t_L g6559 ( 
.A(n_136),
.Y(n_6559)
);

CKINVDCx20_ASAP7_75t_R g6560 ( 
.A(n_2360),
.Y(n_6560)
);

BUFx6f_ASAP7_75t_L g6561 ( 
.A(n_3117),
.Y(n_6561)
);

CKINVDCx5p33_ASAP7_75t_R g6562 ( 
.A(n_2284),
.Y(n_6562)
);

INVx3_ASAP7_75t_L g6563 ( 
.A(n_2197),
.Y(n_6563)
);

CKINVDCx5p33_ASAP7_75t_R g6564 ( 
.A(n_938),
.Y(n_6564)
);

CKINVDCx5p33_ASAP7_75t_R g6565 ( 
.A(n_3813),
.Y(n_6565)
);

CKINVDCx20_ASAP7_75t_R g6566 ( 
.A(n_424),
.Y(n_6566)
);

CKINVDCx5p33_ASAP7_75t_R g6567 ( 
.A(n_1788),
.Y(n_6567)
);

CKINVDCx5p33_ASAP7_75t_R g6568 ( 
.A(n_324),
.Y(n_6568)
);

CKINVDCx5p33_ASAP7_75t_R g6569 ( 
.A(n_4544),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_4387),
.Y(n_6570)
);

CKINVDCx5p33_ASAP7_75t_R g6571 ( 
.A(n_640),
.Y(n_6571)
);

CKINVDCx5p33_ASAP7_75t_R g6572 ( 
.A(n_2820),
.Y(n_6572)
);

INVx2_ASAP7_75t_L g6573 ( 
.A(n_4242),
.Y(n_6573)
);

INVx2_ASAP7_75t_L g6574 ( 
.A(n_4428),
.Y(n_6574)
);

CKINVDCx5p33_ASAP7_75t_R g6575 ( 
.A(n_4028),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_113),
.Y(n_6576)
);

CKINVDCx20_ASAP7_75t_R g6577 ( 
.A(n_1407),
.Y(n_6577)
);

CKINVDCx5p33_ASAP7_75t_R g6578 ( 
.A(n_259),
.Y(n_6578)
);

INVx2_ASAP7_75t_L g6579 ( 
.A(n_3310),
.Y(n_6579)
);

CKINVDCx5p33_ASAP7_75t_R g6580 ( 
.A(n_314),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_2846),
.Y(n_6581)
);

CKINVDCx5p33_ASAP7_75t_R g6582 ( 
.A(n_4848),
.Y(n_6582)
);

CKINVDCx5p33_ASAP7_75t_R g6583 ( 
.A(n_1614),
.Y(n_6583)
);

CKINVDCx5p33_ASAP7_75t_R g6584 ( 
.A(n_4396),
.Y(n_6584)
);

CKINVDCx5p33_ASAP7_75t_R g6585 ( 
.A(n_4538),
.Y(n_6585)
);

CKINVDCx5p33_ASAP7_75t_R g6586 ( 
.A(n_4523),
.Y(n_6586)
);

CKINVDCx5p33_ASAP7_75t_R g6587 ( 
.A(n_2133),
.Y(n_6587)
);

CKINVDCx5p33_ASAP7_75t_R g6588 ( 
.A(n_1268),
.Y(n_6588)
);

CKINVDCx5p33_ASAP7_75t_R g6589 ( 
.A(n_4444),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_4266),
.Y(n_6590)
);

CKINVDCx5p33_ASAP7_75t_R g6591 ( 
.A(n_4119),
.Y(n_6591)
);

INVx1_ASAP7_75t_L g6592 ( 
.A(n_2000),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_2393),
.Y(n_6593)
);

CKINVDCx5p33_ASAP7_75t_R g6594 ( 
.A(n_4543),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_77),
.Y(n_6595)
);

CKINVDCx5p33_ASAP7_75t_R g6596 ( 
.A(n_3916),
.Y(n_6596)
);

CKINVDCx5p33_ASAP7_75t_R g6597 ( 
.A(n_1921),
.Y(n_6597)
);

INVx1_ASAP7_75t_L g6598 ( 
.A(n_484),
.Y(n_6598)
);

CKINVDCx5p33_ASAP7_75t_R g6599 ( 
.A(n_5162),
.Y(n_6599)
);

INVx2_ASAP7_75t_L g6600 ( 
.A(n_2258),
.Y(n_6600)
);

CKINVDCx5p33_ASAP7_75t_R g6601 ( 
.A(n_1575),
.Y(n_6601)
);

CKINVDCx5p33_ASAP7_75t_R g6602 ( 
.A(n_4472),
.Y(n_6602)
);

CKINVDCx5p33_ASAP7_75t_R g6603 ( 
.A(n_4066),
.Y(n_6603)
);

CKINVDCx5p33_ASAP7_75t_R g6604 ( 
.A(n_4158),
.Y(n_6604)
);

INVx2_ASAP7_75t_L g6605 ( 
.A(n_1696),
.Y(n_6605)
);

CKINVDCx5p33_ASAP7_75t_R g6606 ( 
.A(n_1675),
.Y(n_6606)
);

BUFx6f_ASAP7_75t_L g6607 ( 
.A(n_572),
.Y(n_6607)
);

INVx2_ASAP7_75t_SL g6608 ( 
.A(n_4906),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_4081),
.Y(n_6609)
);

CKINVDCx5p33_ASAP7_75t_R g6610 ( 
.A(n_2049),
.Y(n_6610)
);

CKINVDCx5p33_ASAP7_75t_R g6611 ( 
.A(n_426),
.Y(n_6611)
);

CKINVDCx20_ASAP7_75t_R g6612 ( 
.A(n_2588),
.Y(n_6612)
);

CKINVDCx5p33_ASAP7_75t_R g6613 ( 
.A(n_2701),
.Y(n_6613)
);

CKINVDCx5p33_ASAP7_75t_R g6614 ( 
.A(n_2988),
.Y(n_6614)
);

CKINVDCx20_ASAP7_75t_R g6615 ( 
.A(n_3615),
.Y(n_6615)
);

INVx2_ASAP7_75t_SL g6616 ( 
.A(n_4909),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_3243),
.Y(n_6617)
);

CKINVDCx5p33_ASAP7_75t_R g6618 ( 
.A(n_1369),
.Y(n_6618)
);

CKINVDCx5p33_ASAP7_75t_R g6619 ( 
.A(n_2518),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_2090),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_4997),
.Y(n_6621)
);

HB1xp67_ASAP7_75t_L g6622 ( 
.A(n_5235),
.Y(n_6622)
);

CKINVDCx5p33_ASAP7_75t_R g6623 ( 
.A(n_5394),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_5203),
.Y(n_6624)
);

CKINVDCx5p33_ASAP7_75t_R g6625 ( 
.A(n_5454),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_5203),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_5203),
.Y(n_6627)
);

CKINVDCx5p33_ASAP7_75t_R g6628 ( 
.A(n_5534),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_5203),
.Y(n_6629)
);

BUFx10_ASAP7_75t_L g6630 ( 
.A(n_5376),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_5203),
.Y(n_6631)
);

CKINVDCx20_ASAP7_75t_R g6632 ( 
.A(n_5381),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_5397),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_5397),
.Y(n_6634)
);

INVx3_ASAP7_75t_L g6635 ( 
.A(n_5208),
.Y(n_6635)
);

CKINVDCx5p33_ASAP7_75t_R g6636 ( 
.A(n_5562),
.Y(n_6636)
);

CKINVDCx5p33_ASAP7_75t_R g6637 ( 
.A(n_5836),
.Y(n_6637)
);

CKINVDCx5p33_ASAP7_75t_R g6638 ( 
.A(n_5895),
.Y(n_6638)
);

CKINVDCx5p33_ASAP7_75t_R g6639 ( 
.A(n_6018),
.Y(n_6639)
);

NOR2xp67_ASAP7_75t_L g6640 ( 
.A(n_5220),
.B(n_0),
.Y(n_6640)
);

CKINVDCx5p33_ASAP7_75t_R g6641 ( 
.A(n_6087),
.Y(n_6641)
);

CKINVDCx5p33_ASAP7_75t_R g6642 ( 
.A(n_6281),
.Y(n_6642)
);

CKINVDCx5p33_ASAP7_75t_R g6643 ( 
.A(n_5193),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_5397),
.Y(n_6644)
);

CKINVDCx5p33_ASAP7_75t_R g6645 ( 
.A(n_5198),
.Y(n_6645)
);

CKINVDCx6p67_ASAP7_75t_R g6646 ( 
.A(n_5236),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_5397),
.Y(n_6647)
);

CKINVDCx5p33_ASAP7_75t_R g6648 ( 
.A(n_5206),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_5397),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_5613),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_5613),
.Y(n_6651)
);

BUFx6f_ASAP7_75t_L g6652 ( 
.A(n_5501),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_5613),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5613),
.Y(n_6654)
);

BUFx2_ASAP7_75t_SL g6655 ( 
.A(n_5688),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_5613),
.Y(n_6656)
);

INVx1_ASAP7_75t_L g6657 ( 
.A(n_5747),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_5747),
.Y(n_6658)
);

CKINVDCx5p33_ASAP7_75t_R g6659 ( 
.A(n_5254),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_5747),
.Y(n_6660)
);

CKINVDCx5p33_ASAP7_75t_R g6661 ( 
.A(n_5279),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_5747),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_5747),
.Y(n_6663)
);

NOR2xp67_ASAP7_75t_L g6664 ( 
.A(n_5220),
.B(n_0),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_5853),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_5853),
.Y(n_6666)
);

CKINVDCx5p33_ASAP7_75t_R g6667 ( 
.A(n_5300),
.Y(n_6667)
);

CKINVDCx5p33_ASAP7_75t_R g6668 ( 
.A(n_5337),
.Y(n_6668)
);

CKINVDCx5p33_ASAP7_75t_R g6669 ( 
.A(n_5369),
.Y(n_6669)
);

INVx1_ASAP7_75t_SL g6670 ( 
.A(n_5275),
.Y(n_6670)
);

BUFx2_ASAP7_75t_L g6671 ( 
.A(n_5414),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_5853),
.Y(n_6672)
);

CKINVDCx5p33_ASAP7_75t_R g6673 ( 
.A(n_5371),
.Y(n_6673)
);

BUFx3_ASAP7_75t_L g6674 ( 
.A(n_6103),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_5853),
.Y(n_6675)
);

CKINVDCx20_ASAP7_75t_R g6676 ( 
.A(n_5726),
.Y(n_6676)
);

CKINVDCx20_ASAP7_75t_R g6677 ( 
.A(n_5875),
.Y(n_6677)
);

CKINVDCx16_ASAP7_75t_R g6678 ( 
.A(n_5292),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_5853),
.Y(n_6679)
);

CKINVDCx5p33_ASAP7_75t_R g6680 ( 
.A(n_5373),
.Y(n_6680)
);

INVxp67_ASAP7_75t_L g6681 ( 
.A(n_5682),
.Y(n_6681)
);

CKINVDCx5p33_ASAP7_75t_R g6682 ( 
.A(n_5412),
.Y(n_6682)
);

NOR2xp67_ASAP7_75t_L g6683 ( 
.A(n_5703),
.B(n_1),
.Y(n_6683)
);

CKINVDCx14_ASAP7_75t_R g6684 ( 
.A(n_5437),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_5936),
.Y(n_6685)
);

CKINVDCx5p33_ASAP7_75t_R g6686 ( 
.A(n_5430),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_5936),
.Y(n_6687)
);

INVx2_ASAP7_75t_L g6688 ( 
.A(n_5936),
.Y(n_6688)
);

CKINVDCx5p33_ASAP7_75t_R g6689 ( 
.A(n_5476),
.Y(n_6689)
);

CKINVDCx5p33_ASAP7_75t_R g6690 ( 
.A(n_5489),
.Y(n_6690)
);

CKINVDCx5p33_ASAP7_75t_R g6691 ( 
.A(n_5508),
.Y(n_6691)
);

BUFx3_ASAP7_75t_L g6692 ( 
.A(n_6103),
.Y(n_6692)
);

CKINVDCx5p33_ASAP7_75t_R g6693 ( 
.A(n_5542),
.Y(n_6693)
);

CKINVDCx5p33_ASAP7_75t_R g6694 ( 
.A(n_5579),
.Y(n_6694)
);

BUFx2_ASAP7_75t_L g6695 ( 
.A(n_5710),
.Y(n_6695)
);

BUFx6f_ASAP7_75t_L g6696 ( 
.A(n_5501),
.Y(n_6696)
);

CKINVDCx5p33_ASAP7_75t_R g6697 ( 
.A(n_5584),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_5936),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_5936),
.Y(n_6699)
);

INVx1_ASAP7_75t_SL g6700 ( 
.A(n_5774),
.Y(n_6700)
);

CKINVDCx5p33_ASAP7_75t_R g6701 ( 
.A(n_5654),
.Y(n_6701)
);

INVx2_ASAP7_75t_L g6702 ( 
.A(n_6021),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6021),
.Y(n_6703)
);

CKINVDCx5p33_ASAP7_75t_R g6704 ( 
.A(n_5672),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6021),
.Y(n_6705)
);

CKINVDCx5p33_ASAP7_75t_R g6706 ( 
.A(n_5712),
.Y(n_6706)
);

CKINVDCx5p33_ASAP7_75t_R g6707 ( 
.A(n_5727),
.Y(n_6707)
);

BUFx3_ASAP7_75t_L g6708 ( 
.A(n_6141),
.Y(n_6708)
);

CKINVDCx5p33_ASAP7_75t_R g6709 ( 
.A(n_5733),
.Y(n_6709)
);

CKINVDCx16_ASAP7_75t_R g6710 ( 
.A(n_5322),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_6021),
.Y(n_6711)
);

INVx1_ASAP7_75t_SL g6712 ( 
.A(n_5852),
.Y(n_6712)
);

CKINVDCx5p33_ASAP7_75t_R g6713 ( 
.A(n_5741),
.Y(n_6713)
);

BUFx2_ASAP7_75t_SL g6714 ( 
.A(n_6048),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6021),
.Y(n_6715)
);

CKINVDCx5p33_ASAP7_75t_R g6716 ( 
.A(n_5780),
.Y(n_6716)
);

BUFx6f_ASAP7_75t_L g6717 ( 
.A(n_5501),
.Y(n_6717)
);

CKINVDCx5p33_ASAP7_75t_R g6718 ( 
.A(n_5811),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6045),
.Y(n_6719)
);

CKINVDCx5p33_ASAP7_75t_R g6720 ( 
.A(n_5812),
.Y(n_6720)
);

CKINVDCx5p33_ASAP7_75t_R g6721 ( 
.A(n_5823),
.Y(n_6721)
);

INVx1_ASAP7_75t_L g6722 ( 
.A(n_6045),
.Y(n_6722)
);

CKINVDCx5p33_ASAP7_75t_R g6723 ( 
.A(n_5866),
.Y(n_6723)
);

INVx2_ASAP7_75t_L g6724 ( 
.A(n_6045),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_6045),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6045),
.Y(n_6726)
);

CKINVDCx5p33_ASAP7_75t_R g6727 ( 
.A(n_5883),
.Y(n_6727)
);

CKINVDCx16_ASAP7_75t_R g6728 ( 
.A(n_5403),
.Y(n_6728)
);

INVx2_ASAP7_75t_L g6729 ( 
.A(n_6321),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6321),
.Y(n_6730)
);

BUFx2_ASAP7_75t_L g6731 ( 
.A(n_5890),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6321),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6321),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6321),
.Y(n_6734)
);

CKINVDCx5p33_ASAP7_75t_R g6735 ( 
.A(n_5888),
.Y(n_6735)
);

INVx3_ASAP7_75t_L g6736 ( 
.A(n_5208),
.Y(n_6736)
);

CKINVDCx5p33_ASAP7_75t_R g6737 ( 
.A(n_5930),
.Y(n_6737)
);

BUFx5_ASAP7_75t_L g6738 ( 
.A(n_5199),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6403),
.Y(n_6739)
);

CKINVDCx5p33_ASAP7_75t_R g6740 ( 
.A(n_6054),
.Y(n_6740)
);

CKINVDCx20_ASAP7_75t_R g6741 ( 
.A(n_6265),
.Y(n_6741)
);

CKINVDCx5p33_ASAP7_75t_R g6742 ( 
.A(n_6080),
.Y(n_6742)
);

OR2x2_ASAP7_75t_L g6743 ( 
.A(n_6152),
.B(n_1),
.Y(n_6743)
);

CKINVDCx5p33_ASAP7_75t_R g6744 ( 
.A(n_6092),
.Y(n_6744)
);

INVx2_ASAP7_75t_L g6745 ( 
.A(n_6403),
.Y(n_6745)
);

BUFx10_ASAP7_75t_L g6746 ( 
.A(n_5382),
.Y(n_6746)
);

INVx2_ASAP7_75t_L g6747 ( 
.A(n_6403),
.Y(n_6747)
);

BUFx6f_ASAP7_75t_L g6748 ( 
.A(n_6360),
.Y(n_6748)
);

CKINVDCx5p33_ASAP7_75t_R g6749 ( 
.A(n_6113),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6403),
.Y(n_6750)
);

CKINVDCx5p33_ASAP7_75t_R g6751 ( 
.A(n_6116),
.Y(n_6751)
);

CKINVDCx5p33_ASAP7_75t_R g6752 ( 
.A(n_6131),
.Y(n_6752)
);

BUFx2_ASAP7_75t_SL g6753 ( 
.A(n_6549),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6403),
.Y(n_6754)
);

CKINVDCx5p33_ASAP7_75t_R g6755 ( 
.A(n_6165),
.Y(n_6755)
);

INVx1_ASAP7_75t_L g6756 ( 
.A(n_6482),
.Y(n_6756)
);

INVx1_ASAP7_75t_L g6757 ( 
.A(n_6482),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6482),
.Y(n_6758)
);

BUFx5_ASAP7_75t_L g6759 ( 
.A(n_5226),
.Y(n_6759)
);

INVx1_ASAP7_75t_L g6760 ( 
.A(n_6482),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6482),
.Y(n_6761)
);

INVx1_ASAP7_75t_SL g6762 ( 
.A(n_6243),
.Y(n_6762)
);

BUFx6f_ASAP7_75t_L g6763 ( 
.A(n_6360),
.Y(n_6763)
);

CKINVDCx5p33_ASAP7_75t_R g6764 ( 
.A(n_6177),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6533),
.Y(n_6765)
);

NAND2xp5_ASAP7_75t_L g6766 ( 
.A(n_5516),
.B(n_3),
.Y(n_6766)
);

BUFx3_ASAP7_75t_L g6767 ( 
.A(n_6141),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6533),
.Y(n_6768)
);

INVx2_ASAP7_75t_SL g6769 ( 
.A(n_5169),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6533),
.Y(n_6770)
);

INVx1_ASAP7_75t_L g6771 ( 
.A(n_6533),
.Y(n_6771)
);

CKINVDCx5p33_ASAP7_75t_R g6772 ( 
.A(n_6186),
.Y(n_6772)
);

CKINVDCx5p33_ASAP7_75t_R g6773 ( 
.A(n_6193),
.Y(n_6773)
);

CKINVDCx5p33_ASAP7_75t_R g6774 ( 
.A(n_6221),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_5722),
.B(n_3),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6533),
.Y(n_6776)
);

CKINVDCx20_ASAP7_75t_R g6777 ( 
.A(n_6338),
.Y(n_6777)
);

CKINVDCx5p33_ASAP7_75t_R g6778 ( 
.A(n_6227),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_5703),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6028),
.Y(n_6780)
);

CKINVDCx5p33_ASAP7_75t_R g6781 ( 
.A(n_6228),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6028),
.Y(n_6782)
);

CKINVDCx20_ASAP7_75t_R g6783 ( 
.A(n_5237),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6094),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6094),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6096),
.Y(n_6786)
);

CKINVDCx5p33_ASAP7_75t_R g6787 ( 
.A(n_6254),
.Y(n_6787)
);

CKINVDCx20_ASAP7_75t_R g6788 ( 
.A(n_5915),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6096),
.Y(n_6789)
);

CKINVDCx5p33_ASAP7_75t_R g6790 ( 
.A(n_6273),
.Y(n_6790)
);

CKINVDCx5p33_ASAP7_75t_R g6791 ( 
.A(n_6301),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_6563),
.Y(n_6792)
);

OR2x2_ASAP7_75t_L g6793 ( 
.A(n_6383),
.B(n_4),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6563),
.Y(n_6794)
);

CKINVDCx5p33_ASAP7_75t_R g6795 ( 
.A(n_6331),
.Y(n_6795)
);

CKINVDCx5p33_ASAP7_75t_R g6796 ( 
.A(n_6357),
.Y(n_6796)
);

CKINVDCx20_ASAP7_75t_R g6797 ( 
.A(n_6025),
.Y(n_6797)
);

BUFx2_ASAP7_75t_L g6798 ( 
.A(n_6491),
.Y(n_6798)
);

HB1xp67_ASAP7_75t_L g6799 ( 
.A(n_5561),
.Y(n_6799)
);

CKINVDCx5p33_ASAP7_75t_R g6800 ( 
.A(n_6361),
.Y(n_6800)
);

CKINVDCx5p33_ASAP7_75t_R g6801 ( 
.A(n_6372),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_5208),
.Y(n_6802)
);

INVx2_ASAP7_75t_L g6803 ( 
.A(n_5211),
.Y(n_6803)
);

BUFx3_ASAP7_75t_L g6804 ( 
.A(n_6307),
.Y(n_6804)
);

CKINVDCx5p33_ASAP7_75t_R g6805 ( 
.A(n_6404),
.Y(n_6805)
);

CKINVDCx5p33_ASAP7_75t_R g6806 ( 
.A(n_6407),
.Y(n_6806)
);

CKINVDCx5p33_ASAP7_75t_R g6807 ( 
.A(n_6450),
.Y(n_6807)
);

CKINVDCx20_ASAP7_75t_R g6808 ( 
.A(n_6090),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_5211),
.Y(n_6809)
);

BUFx6f_ASAP7_75t_L g6810 ( 
.A(n_6360),
.Y(n_6810)
);

CKINVDCx5p33_ASAP7_75t_R g6811 ( 
.A(n_6458),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_5211),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_5234),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_5234),
.Y(n_6814)
);

CKINVDCx20_ASAP7_75t_R g6815 ( 
.A(n_6118),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_5234),
.Y(n_6816)
);

CKINVDCx5p33_ASAP7_75t_R g6817 ( 
.A(n_6460),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_5344),
.Y(n_6818)
);

CKINVDCx5p33_ASAP7_75t_R g6819 ( 
.A(n_6471),
.Y(n_6819)
);

CKINVDCx16_ASAP7_75t_R g6820 ( 
.A(n_5738),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_5344),
.Y(n_6821)
);

INVx1_ASAP7_75t_L g6822 ( 
.A(n_5344),
.Y(n_6822)
);

CKINVDCx5p33_ASAP7_75t_R g6823 ( 
.A(n_6493),
.Y(n_6823)
);

CKINVDCx5p33_ASAP7_75t_R g6824 ( 
.A(n_6508),
.Y(n_6824)
);

CKINVDCx5p33_ASAP7_75t_R g6825 ( 
.A(n_6509),
.Y(n_6825)
);

HB1xp67_ASAP7_75t_L g6826 ( 
.A(n_5827),
.Y(n_6826)
);

BUFx10_ASAP7_75t_L g6827 ( 
.A(n_6261),
.Y(n_6827)
);

CKINVDCx5p33_ASAP7_75t_R g6828 ( 
.A(n_6515),
.Y(n_6828)
);

INVx2_ASAP7_75t_L g6829 ( 
.A(n_5367),
.Y(n_6829)
);

CKINVDCx5p33_ASAP7_75t_R g6830 ( 
.A(n_6522),
.Y(n_6830)
);

INVx1_ASAP7_75t_SL g6831 ( 
.A(n_6527),
.Y(n_6831)
);

CKINVDCx5p33_ASAP7_75t_R g6832 ( 
.A(n_6539),
.Y(n_6832)
);

CKINVDCx5p33_ASAP7_75t_R g6833 ( 
.A(n_6540),
.Y(n_6833)
);

CKINVDCx5p33_ASAP7_75t_R g6834 ( 
.A(n_6548),
.Y(n_6834)
);

CKINVDCx5p33_ASAP7_75t_R g6835 ( 
.A(n_6551),
.Y(n_6835)
);

CKINVDCx5p33_ASAP7_75t_R g6836 ( 
.A(n_6582),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_5367),
.Y(n_6837)
);

CKINVDCx5p33_ASAP7_75t_R g6838 ( 
.A(n_6599),
.Y(n_6838)
);

CKINVDCx5p33_ASAP7_75t_R g6839 ( 
.A(n_6150),
.Y(n_6839)
);

CKINVDCx5p33_ASAP7_75t_R g6840 ( 
.A(n_6203),
.Y(n_6840)
);

BUFx2_ASAP7_75t_L g6841 ( 
.A(n_6559),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_5367),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_5464),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_5464),
.Y(n_6844)
);

CKINVDCx5p33_ASAP7_75t_R g6845 ( 
.A(n_6310),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_5464),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_5485),
.Y(n_6847)
);

HB1xp67_ASAP7_75t_L g6848 ( 
.A(n_5856),
.Y(n_6848)
);

INVx1_ASAP7_75t_L g6849 ( 
.A(n_5485),
.Y(n_6849)
);

INVx2_ASAP7_75t_L g6850 ( 
.A(n_5485),
.Y(n_6850)
);

BUFx3_ASAP7_75t_L g6851 ( 
.A(n_6307),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_5523),
.Y(n_6852)
);

CKINVDCx5p33_ASAP7_75t_R g6853 ( 
.A(n_5967),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_5523),
.Y(n_6854)
);

CKINVDCx5p33_ASAP7_75t_R g6855 ( 
.A(n_6006),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_5523),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_5570),
.Y(n_6857)
);

INVx1_ASAP7_75t_L g6858 ( 
.A(n_5570),
.Y(n_6858)
);

CKINVDCx5p33_ASAP7_75t_R g6859 ( 
.A(n_6052),
.Y(n_6859)
);

HB1xp67_ASAP7_75t_L g6860 ( 
.A(n_6149),
.Y(n_6860)
);

CKINVDCx20_ASAP7_75t_R g6861 ( 
.A(n_5228),
.Y(n_6861)
);

CKINVDCx20_ASAP7_75t_R g6862 ( 
.A(n_6401),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_5570),
.Y(n_6863)
);

CKINVDCx5p33_ASAP7_75t_R g6864 ( 
.A(n_6294),
.Y(n_6864)
);

INVxp67_ASAP7_75t_SL g6865 ( 
.A(n_5495),
.Y(n_6865)
);

CKINVDCx5p33_ASAP7_75t_R g6866 ( 
.A(n_6424),
.Y(n_6866)
);

CKINVDCx5p33_ASAP7_75t_R g6867 ( 
.A(n_6444),
.Y(n_6867)
);

CKINVDCx5p33_ASAP7_75t_R g6868 ( 
.A(n_6466),
.Y(n_6868)
);

CKINVDCx5p33_ASAP7_75t_R g6869 ( 
.A(n_6525),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_5615),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_5615),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_5615),
.Y(n_6872)
);

NAND2xp5_ASAP7_75t_L g6873 ( 
.A(n_5345),
.B(n_4),
.Y(n_6873)
);

INVx1_ASAP7_75t_SL g6874 ( 
.A(n_5299),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_5687),
.Y(n_6875)
);

INVx2_ASAP7_75t_L g6876 ( 
.A(n_5687),
.Y(n_6876)
);

HB1xp67_ASAP7_75t_L g6877 ( 
.A(n_5897),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_5687),
.Y(n_6878)
);

CKINVDCx16_ASAP7_75t_R g6879 ( 
.A(n_5169),
.Y(n_6879)
);

BUFx8_ASAP7_75t_SL g6880 ( 
.A(n_5187),
.Y(n_6880)
);

CKINVDCx5p33_ASAP7_75t_R g6881 ( 
.A(n_6610),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_5711),
.Y(n_6882)
);

CKINVDCx20_ASAP7_75t_R g6883 ( 
.A(n_5784),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_5711),
.Y(n_6884)
);

INVxp67_ASAP7_75t_L g6885 ( 
.A(n_6167),
.Y(n_6885)
);

INVx2_ASAP7_75t_L g6886 ( 
.A(n_5711),
.Y(n_6886)
);

INVx2_ASAP7_75t_L g6887 ( 
.A(n_5735),
.Y(n_6887)
);

CKINVDCx5p33_ASAP7_75t_R g6888 ( 
.A(n_6613),
.Y(n_6888)
);

CKINVDCx5p33_ASAP7_75t_R g6889 ( 
.A(n_6614),
.Y(n_6889)
);

CKINVDCx5p33_ASAP7_75t_R g6890 ( 
.A(n_6618),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_5735),
.Y(n_6891)
);

HB1xp67_ASAP7_75t_L g6892 ( 
.A(n_6468),
.Y(n_6892)
);

CKINVDCx5p33_ASAP7_75t_R g6893 ( 
.A(n_6619),
.Y(n_6893)
);

CKINVDCx5p33_ASAP7_75t_R g6894 ( 
.A(n_5171),
.Y(n_6894)
);

CKINVDCx5p33_ASAP7_75t_R g6895 ( 
.A(n_5173),
.Y(n_6895)
);

BUFx6f_ASAP7_75t_L g6896 ( 
.A(n_6494),
.Y(n_6896)
);

CKINVDCx5p33_ASAP7_75t_R g6897 ( 
.A(n_5174),
.Y(n_6897)
);

BUFx3_ASAP7_75t_L g6898 ( 
.A(n_6409),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_5735),
.Y(n_6899)
);

CKINVDCx5p33_ASAP7_75t_R g6900 ( 
.A(n_5175),
.Y(n_6900)
);

BUFx6f_ASAP7_75t_L g6901 ( 
.A(n_6494),
.Y(n_6901)
);

NOR2xp67_ASAP7_75t_L g6902 ( 
.A(n_5510),
.B(n_5),
.Y(n_6902)
);

CKINVDCx16_ASAP7_75t_R g6903 ( 
.A(n_5213),
.Y(n_6903)
);

HB1xp67_ASAP7_75t_L g6904 ( 
.A(n_6534),
.Y(n_6904)
);

INVx2_ASAP7_75t_L g6905 ( 
.A(n_6607),
.Y(n_6905)
);

INVxp67_ASAP7_75t_L g6906 ( 
.A(n_5213),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6607),
.Y(n_6907)
);

CKINVDCx5p33_ASAP7_75t_R g6908 ( 
.A(n_6604),
.Y(n_6908)
);

BUFx10_ASAP7_75t_L g6909 ( 
.A(n_5742),
.Y(n_6909)
);

CKINVDCx5p33_ASAP7_75t_R g6910 ( 
.A(n_6606),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_5742),
.Y(n_6911)
);

CKINVDCx5p33_ASAP7_75t_R g6912 ( 
.A(n_6611),
.Y(n_6912)
);

CKINVDCx5p33_ASAP7_75t_R g6913 ( 
.A(n_5177),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_5742),
.Y(n_6914)
);

CKINVDCx5p33_ASAP7_75t_R g6915 ( 
.A(n_5178),
.Y(n_6915)
);

CKINVDCx5p33_ASAP7_75t_R g6916 ( 
.A(n_5181),
.Y(n_6916)
);

CKINVDCx5p33_ASAP7_75t_R g6917 ( 
.A(n_5183),
.Y(n_6917)
);

CKINVDCx5p33_ASAP7_75t_R g6918 ( 
.A(n_5184),
.Y(n_6918)
);

INVxp33_ASAP7_75t_L g6919 ( 
.A(n_5651),
.Y(n_6919)
);

INVx1_ASAP7_75t_L g6920 ( 
.A(n_5757),
.Y(n_6920)
);

CKINVDCx5p33_ASAP7_75t_R g6921 ( 
.A(n_5190),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_5757),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_5757),
.Y(n_6923)
);

CKINVDCx5p33_ASAP7_75t_R g6924 ( 
.A(n_5191),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_5820),
.Y(n_6925)
);

INVx1_ASAP7_75t_L g6926 ( 
.A(n_5820),
.Y(n_6926)
);

CKINVDCx5p33_ASAP7_75t_R g6927 ( 
.A(n_5192),
.Y(n_6927)
);

CKINVDCx20_ASAP7_75t_R g6928 ( 
.A(n_5232),
.Y(n_6928)
);

INVxp67_ASAP7_75t_SL g6929 ( 
.A(n_5629),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_5820),
.Y(n_6930)
);

BUFx3_ASAP7_75t_L g6931 ( 
.A(n_6409),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_5824),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_5824),
.Y(n_6933)
);

CKINVDCx5p33_ASAP7_75t_R g6934 ( 
.A(n_6603),
.Y(n_6934)
);

CKINVDCx5p33_ASAP7_75t_R g6935 ( 
.A(n_5196),
.Y(n_6935)
);

INVx3_ASAP7_75t_L g6936 ( 
.A(n_5824),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_5826),
.Y(n_6937)
);

CKINVDCx5p33_ASAP7_75t_R g6938 ( 
.A(n_5197),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_5826),
.Y(n_6939)
);

CKINVDCx5p33_ASAP7_75t_R g6940 ( 
.A(n_5200),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_5826),
.Y(n_6941)
);

CKINVDCx5p33_ASAP7_75t_R g6942 ( 
.A(n_5201),
.Y(n_6942)
);

CKINVDCx5p33_ASAP7_75t_R g6943 ( 
.A(n_5204),
.Y(n_6943)
);

BUFx3_ASAP7_75t_L g6944 ( 
.A(n_5424),
.Y(n_6944)
);

INVx1_ASAP7_75t_SL g6945 ( 
.A(n_5252),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_5924),
.Y(n_6946)
);

CKINVDCx5p33_ASAP7_75t_R g6947 ( 
.A(n_5205),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_5924),
.Y(n_6948)
);

INVx2_ASAP7_75t_L g6949 ( 
.A(n_5924),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_5938),
.Y(n_6950)
);

INVx2_ASAP7_75t_L g6951 ( 
.A(n_6607),
.Y(n_6951)
);

HB1xp67_ASAP7_75t_L g6952 ( 
.A(n_5450),
.Y(n_6952)
);

CKINVDCx20_ASAP7_75t_R g6953 ( 
.A(n_5246),
.Y(n_6953)
);

CKINVDCx20_ASAP7_75t_R g6954 ( 
.A(n_5250),
.Y(n_6954)
);

CKINVDCx5p33_ASAP7_75t_R g6955 ( 
.A(n_6601),
.Y(n_6955)
);

CKINVDCx5p33_ASAP7_75t_R g6956 ( 
.A(n_6602),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_5938),
.Y(n_6957)
);

CKINVDCx5p33_ASAP7_75t_R g6958 ( 
.A(n_5207),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_5938),
.Y(n_6959)
);

CKINVDCx5p33_ASAP7_75t_R g6960 ( 
.A(n_5210),
.Y(n_6960)
);

CKINVDCx5p33_ASAP7_75t_R g6961 ( 
.A(n_5212),
.Y(n_6961)
);

CKINVDCx5p33_ASAP7_75t_R g6962 ( 
.A(n_5217),
.Y(n_6962)
);

CKINVDCx20_ASAP7_75t_R g6963 ( 
.A(n_5262),
.Y(n_6963)
);

INVxp33_ASAP7_75t_L g6964 ( 
.A(n_5170),
.Y(n_6964)
);

CKINVDCx20_ASAP7_75t_R g6965 ( 
.A(n_5288),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_5953),
.Y(n_6966)
);

INVx2_ASAP7_75t_L g6967 ( 
.A(n_5953),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_5953),
.Y(n_6968)
);

CKINVDCx20_ASAP7_75t_R g6969 ( 
.A(n_5295),
.Y(n_6969)
);

CKINVDCx5p33_ASAP7_75t_R g6970 ( 
.A(n_6594),
.Y(n_6970)
);

INVx2_ASAP7_75t_L g6971 ( 
.A(n_5966),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_5966),
.Y(n_6972)
);

CKINVDCx5p33_ASAP7_75t_R g6973 ( 
.A(n_6596),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_5966),
.Y(n_6974)
);

BUFx3_ASAP7_75t_L g6975 ( 
.A(n_5537),
.Y(n_6975)
);

INVxp33_ASAP7_75t_SL g6976 ( 
.A(n_5218),
.Y(n_6976)
);

CKINVDCx5p33_ASAP7_75t_R g6977 ( 
.A(n_5219),
.Y(n_6977)
);

CKINVDCx5p33_ASAP7_75t_R g6978 ( 
.A(n_5221),
.Y(n_6978)
);

CKINVDCx5p33_ASAP7_75t_R g6979 ( 
.A(n_5225),
.Y(n_6979)
);

CKINVDCx5p33_ASAP7_75t_R g6980 ( 
.A(n_5227),
.Y(n_6980)
);

INVx1_ASAP7_75t_L g6981 ( 
.A(n_5980),
.Y(n_6981)
);

CKINVDCx5p33_ASAP7_75t_R g6982 ( 
.A(n_5230),
.Y(n_6982)
);

CKINVDCx5p33_ASAP7_75t_R g6983 ( 
.A(n_5233),
.Y(n_6983)
);

CKINVDCx20_ASAP7_75t_R g6984 ( 
.A(n_5306),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_5980),
.Y(n_6985)
);

CKINVDCx5p33_ASAP7_75t_R g6986 ( 
.A(n_5238),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_5980),
.Y(n_6987)
);

CKINVDCx5p33_ASAP7_75t_R g6988 ( 
.A(n_5240),
.Y(n_6988)
);

CKINVDCx5p33_ASAP7_75t_R g6989 ( 
.A(n_5241),
.Y(n_6989)
);

CKINVDCx5p33_ASAP7_75t_R g6990 ( 
.A(n_6597),
.Y(n_6990)
);

INVx2_ASAP7_75t_L g6991 ( 
.A(n_6047),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_6608),
.B(n_5),
.Y(n_6992)
);

CKINVDCx5p33_ASAP7_75t_R g6993 ( 
.A(n_5247),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_6047),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6047),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6060),
.Y(n_6996)
);

CKINVDCx5p33_ASAP7_75t_R g6997 ( 
.A(n_5248),
.Y(n_6997)
);

CKINVDCx5p33_ASAP7_75t_R g6998 ( 
.A(n_5251),
.Y(n_6998)
);

NOR2xp67_ASAP7_75t_L g6999 ( 
.A(n_5611),
.B(n_6),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6060),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6060),
.Y(n_7001)
);

CKINVDCx5p33_ASAP7_75t_R g7002 ( 
.A(n_5255),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6076),
.Y(n_7003)
);

CKINVDCx5p33_ASAP7_75t_R g7004 ( 
.A(n_5256),
.Y(n_7004)
);

CKINVDCx5p33_ASAP7_75t_R g7005 ( 
.A(n_5257),
.Y(n_7005)
);

INVx1_ASAP7_75t_L g7006 ( 
.A(n_6076),
.Y(n_7006)
);

CKINVDCx5p33_ASAP7_75t_R g7007 ( 
.A(n_5258),
.Y(n_7007)
);

BUFx3_ASAP7_75t_L g7008 ( 
.A(n_5546),
.Y(n_7008)
);

CKINVDCx20_ASAP7_75t_R g7009 ( 
.A(n_5324),
.Y(n_7009)
);

BUFx6f_ASAP7_75t_L g7010 ( 
.A(n_6494),
.Y(n_7010)
);

CKINVDCx5p33_ASAP7_75t_R g7011 ( 
.A(n_5260),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6076),
.Y(n_7012)
);

BUFx5_ASAP7_75t_L g7013 ( 
.A(n_5231),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6219),
.Y(n_7014)
);

BUFx10_ASAP7_75t_L g7015 ( 
.A(n_6219),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_6219),
.Y(n_7016)
);

INVxp33_ASAP7_75t_L g7017 ( 
.A(n_5172),
.Y(n_7017)
);

CKINVDCx5p33_ASAP7_75t_R g7018 ( 
.A(n_5261),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6350),
.Y(n_7019)
);

CKINVDCx5p33_ASAP7_75t_R g7020 ( 
.A(n_5264),
.Y(n_7020)
);

CKINVDCx16_ASAP7_75t_R g7021 ( 
.A(n_5308),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6350),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6350),
.Y(n_7023)
);

CKINVDCx5p33_ASAP7_75t_R g7024 ( 
.A(n_5265),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6381),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6381),
.Y(n_7026)
);

CKINVDCx5p33_ASAP7_75t_R g7027 ( 
.A(n_5266),
.Y(n_7027)
);

CKINVDCx5p33_ASAP7_75t_R g7028 ( 
.A(n_5268),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6381),
.Y(n_7029)
);

CKINVDCx5p33_ASAP7_75t_R g7030 ( 
.A(n_5272),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6478),
.Y(n_7031)
);

CKINVDCx5p33_ASAP7_75t_R g7032 ( 
.A(n_5273),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6478),
.Y(n_7033)
);

CKINVDCx5p33_ASAP7_75t_R g7034 ( 
.A(n_5277),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6478),
.Y(n_7035)
);

CKINVDCx20_ASAP7_75t_R g7036 ( 
.A(n_5370),
.Y(n_7036)
);

INVx1_ASAP7_75t_L g7037 ( 
.A(n_6503),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6503),
.Y(n_7038)
);

CKINVDCx5p33_ASAP7_75t_R g7039 ( 
.A(n_6591),
.Y(n_7039)
);

INVx1_ASAP7_75t_L g7040 ( 
.A(n_6503),
.Y(n_7040)
);

BUFx10_ASAP7_75t_L g7041 ( 
.A(n_6557),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6557),
.Y(n_7042)
);

CKINVDCx5p33_ASAP7_75t_R g7043 ( 
.A(n_5284),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6557),
.Y(n_7044)
);

CKINVDCx5p33_ASAP7_75t_R g7045 ( 
.A(n_5289),
.Y(n_7045)
);

CKINVDCx5p33_ASAP7_75t_R g7046 ( 
.A(n_5291),
.Y(n_7046)
);

CKINVDCx5p33_ASAP7_75t_R g7047 ( 
.A(n_5294),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6561),
.Y(n_7048)
);

CKINVDCx5p33_ASAP7_75t_R g7049 ( 
.A(n_5297),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6561),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6561),
.Y(n_7051)
);

CKINVDCx5p33_ASAP7_75t_R g7052 ( 
.A(n_5303),
.Y(n_7052)
);

CKINVDCx12_ASAP7_75t_R g7053 ( 
.A(n_5189),
.Y(n_7053)
);

INVx1_ASAP7_75t_SL g7054 ( 
.A(n_5551),
.Y(n_7054)
);

CKINVDCx5p33_ASAP7_75t_R g7055 ( 
.A(n_5304),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_5612),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_5620),
.Y(n_7057)
);

INVx2_ASAP7_75t_SL g7058 ( 
.A(n_5308),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_5664),
.Y(n_7059)
);

CKINVDCx5p33_ASAP7_75t_R g7060 ( 
.A(n_5313),
.Y(n_7060)
);

CKINVDCx5p33_ASAP7_75t_R g7061 ( 
.A(n_5315),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_5676),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_5683),
.Y(n_7063)
);

CKINVDCx5p33_ASAP7_75t_R g7064 ( 
.A(n_5317),
.Y(n_7064)
);

CKINVDCx5p33_ASAP7_75t_R g7065 ( 
.A(n_5318),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_5758),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_5814),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_5816),
.Y(n_7068)
);

CKINVDCx5p33_ASAP7_75t_R g7069 ( 
.A(n_5319),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_5858),
.Y(n_7070)
);

CKINVDCx5p33_ASAP7_75t_R g7071 ( 
.A(n_5323),
.Y(n_7071)
);

CKINVDCx5p33_ASAP7_75t_R g7072 ( 
.A(n_5326),
.Y(n_7072)
);

CKINVDCx5p33_ASAP7_75t_R g7073 ( 
.A(n_5328),
.Y(n_7073)
);

CKINVDCx5p33_ASAP7_75t_R g7074 ( 
.A(n_5329),
.Y(n_7074)
);

CKINVDCx20_ASAP7_75t_R g7075 ( 
.A(n_5378),
.Y(n_7075)
);

NOR2xp67_ASAP7_75t_L g7076 ( 
.A(n_5619),
.B(n_6),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_5931),
.Y(n_7077)
);

INVxp67_ASAP7_75t_L g7078 ( 
.A(n_5331),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_5942),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_5949),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_5179),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_6098),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6111),
.Y(n_7083)
);

CKINVDCx20_ASAP7_75t_R g7084 ( 
.A(n_6632),
.Y(n_7084)
);

INVx3_ASAP7_75t_L g7085 ( 
.A(n_6652),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6803),
.Y(n_7086)
);

INVxp67_ASAP7_75t_L g7087 ( 
.A(n_6622),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_6829),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6850),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6876),
.Y(n_7090)
);

INVx1_ASAP7_75t_L g7091 ( 
.A(n_6886),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6887),
.Y(n_7092)
);

INVx2_ASAP7_75t_L g7093 ( 
.A(n_6905),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6907),
.Y(n_7094)
);

CKINVDCx5p33_ASAP7_75t_R g7095 ( 
.A(n_6643),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_6949),
.Y(n_7096)
);

CKINVDCx20_ASAP7_75t_R g7097 ( 
.A(n_6676),
.Y(n_7097)
);

HB1xp67_ASAP7_75t_L g7098 ( 
.A(n_6853),
.Y(n_7098)
);

INVxp67_ASAP7_75t_L g7099 ( 
.A(n_6799),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_6951),
.Y(n_7100)
);

INVx1_ASAP7_75t_L g7101 ( 
.A(n_6967),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6971),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6991),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_6802),
.Y(n_7104)
);

INVx1_ASAP7_75t_SL g7105 ( 
.A(n_6874),
.Y(n_7105)
);

INVxp67_ASAP7_75t_SL g7106 ( 
.A(n_6865),
.Y(n_7106)
);

CKINVDCx5p33_ASAP7_75t_R g7107 ( 
.A(n_6645),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6809),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6812),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_6813),
.Y(n_7110)
);

CKINVDCx5p33_ASAP7_75t_R g7111 ( 
.A(n_6648),
.Y(n_7111)
);

CKINVDCx20_ASAP7_75t_R g7112 ( 
.A(n_6677),
.Y(n_7112)
);

CKINVDCx20_ASAP7_75t_R g7113 ( 
.A(n_6741),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6814),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6816),
.Y(n_7115)
);

CKINVDCx16_ASAP7_75t_R g7116 ( 
.A(n_6788),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6818),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6821),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6822),
.Y(n_7119)
);

BUFx2_ASAP7_75t_L g7120 ( 
.A(n_6797),
.Y(n_7120)
);

INVx2_ASAP7_75t_L g7121 ( 
.A(n_6652),
.Y(n_7121)
);

INVxp67_ASAP7_75t_L g7122 ( 
.A(n_6826),
.Y(n_7122)
);

CKINVDCx5p33_ASAP7_75t_R g7123 ( 
.A(n_6659),
.Y(n_7123)
);

CKINVDCx20_ASAP7_75t_R g7124 ( 
.A(n_6783),
.Y(n_7124)
);

CKINVDCx16_ASAP7_75t_R g7125 ( 
.A(n_6808),
.Y(n_7125)
);

INVxp67_ASAP7_75t_L g7126 ( 
.A(n_6848),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6837),
.Y(n_7127)
);

XOR2x2_ASAP7_75t_L g7128 ( 
.A(n_6945),
.B(n_5673),
.Y(n_7128)
);

CKINVDCx16_ASAP7_75t_R g7129 ( 
.A(n_6815),
.Y(n_7129)
);

CKINVDCx5p33_ASAP7_75t_R g7130 ( 
.A(n_6661),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6842),
.Y(n_7131)
);

HB1xp67_ASAP7_75t_L g7132 ( 
.A(n_6855),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6843),
.Y(n_7133)
);

INVx2_ASAP7_75t_L g7134 ( 
.A(n_6652),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6844),
.Y(n_7135)
);

CKINVDCx5p33_ASAP7_75t_R g7136 ( 
.A(n_6667),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6846),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6847),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_6849),
.Y(n_7139)
);

INVx1_ASAP7_75t_L g7140 ( 
.A(n_6852),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6854),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6696),
.Y(n_7142)
);

CKINVDCx16_ASAP7_75t_R g7143 ( 
.A(n_6678),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_6856),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6696),
.Y(n_7145)
);

CKINVDCx20_ASAP7_75t_R g7146 ( 
.A(n_6928),
.Y(n_7146)
);

INVxp67_ASAP7_75t_SL g7147 ( 
.A(n_6952),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6857),
.Y(n_7148)
);

CKINVDCx5p33_ASAP7_75t_R g7149 ( 
.A(n_6668),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_6858),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6863),
.Y(n_7151)
);

HB1xp67_ASAP7_75t_L g7152 ( 
.A(n_6859),
.Y(n_7152)
);

CKINVDCx20_ASAP7_75t_R g7153 ( 
.A(n_6953),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_6870),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6871),
.Y(n_7155)
);

CKINVDCx20_ASAP7_75t_R g7156 ( 
.A(n_6954),
.Y(n_7156)
);

INVx2_ASAP7_75t_L g7157 ( 
.A(n_6696),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6872),
.Y(n_7158)
);

CKINVDCx5p33_ASAP7_75t_R g7159 ( 
.A(n_6669),
.Y(n_7159)
);

INVxp67_ASAP7_75t_L g7160 ( 
.A(n_6860),
.Y(n_7160)
);

CKINVDCx5p33_ASAP7_75t_R g7161 ( 
.A(n_6673),
.Y(n_7161)
);

INVx2_ASAP7_75t_SL g7162 ( 
.A(n_6630),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_6875),
.Y(n_7163)
);

CKINVDCx5p33_ASAP7_75t_R g7164 ( 
.A(n_6680),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6878),
.Y(n_7165)
);

CKINVDCx5p33_ASAP7_75t_R g7166 ( 
.A(n_6682),
.Y(n_7166)
);

INVx2_ASAP7_75t_L g7167 ( 
.A(n_6717),
.Y(n_7167)
);

CKINVDCx20_ASAP7_75t_R g7168 ( 
.A(n_6963),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6882),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_6884),
.Y(n_7170)
);

INVx2_ASAP7_75t_L g7171 ( 
.A(n_6717),
.Y(n_7171)
);

CKINVDCx5p33_ASAP7_75t_R g7172 ( 
.A(n_6686),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_6891),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_6899),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6911),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_6914),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6920),
.Y(n_7177)
);

CKINVDCx16_ASAP7_75t_R g7178 ( 
.A(n_6710),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_6922),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6923),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6925),
.Y(n_7181)
);

INVxp67_ASAP7_75t_L g7182 ( 
.A(n_6674),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6926),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6930),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_6932),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_6933),
.Y(n_7186)
);

INVxp67_ASAP7_75t_SL g7187 ( 
.A(n_6766),
.Y(n_7187)
);

CKINVDCx5p33_ASAP7_75t_R g7188 ( 
.A(n_6689),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_6937),
.Y(n_7189)
);

CKINVDCx5p33_ASAP7_75t_R g7190 ( 
.A(n_6690),
.Y(n_7190)
);

INVxp67_ASAP7_75t_SL g7191 ( 
.A(n_6775),
.Y(n_7191)
);

CKINVDCx5p33_ASAP7_75t_R g7192 ( 
.A(n_6691),
.Y(n_7192)
);

CKINVDCx16_ASAP7_75t_R g7193 ( 
.A(n_6728),
.Y(n_7193)
);

BUFx6f_ASAP7_75t_L g7194 ( 
.A(n_6717),
.Y(n_7194)
);

CKINVDCx5p33_ASAP7_75t_R g7195 ( 
.A(n_6693),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_6939),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_6941),
.Y(n_7197)
);

BUFx3_ASAP7_75t_L g7198 ( 
.A(n_6944),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6946),
.Y(n_7199)
);

CKINVDCx5p33_ASAP7_75t_R g7200 ( 
.A(n_6694),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6948),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6950),
.Y(n_7202)
);

CKINVDCx5p33_ASAP7_75t_R g7203 ( 
.A(n_6697),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_6957),
.Y(n_7204)
);

INVxp67_ASAP7_75t_SL g7205 ( 
.A(n_6975),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_6959),
.Y(n_7206)
);

CKINVDCx20_ASAP7_75t_R g7207 ( 
.A(n_6965),
.Y(n_7207)
);

HB1xp67_ASAP7_75t_L g7208 ( 
.A(n_6864),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_6966),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_6968),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_6972),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6974),
.Y(n_7212)
);

INVxp67_ASAP7_75t_L g7213 ( 
.A(n_6692),
.Y(n_7213)
);

CKINVDCx16_ASAP7_75t_R g7214 ( 
.A(n_6820),
.Y(n_7214)
);

CKINVDCx5p33_ASAP7_75t_R g7215 ( 
.A(n_6701),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_6748),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_6981),
.Y(n_7217)
);

INVx1_ASAP7_75t_L g7218 ( 
.A(n_6985),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_6987),
.Y(n_7219)
);

INVx1_ASAP7_75t_L g7220 ( 
.A(n_6994),
.Y(n_7220)
);

INVxp67_ASAP7_75t_SL g7221 ( 
.A(n_7008),
.Y(n_7221)
);

INVxp67_ASAP7_75t_L g7222 ( 
.A(n_6708),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6995),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_6996),
.Y(n_7224)
);

CKINVDCx20_ASAP7_75t_R g7225 ( 
.A(n_6969),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7000),
.Y(n_7226)
);

INVxp67_ASAP7_75t_SL g7227 ( 
.A(n_6748),
.Y(n_7227)
);

CKINVDCx5p33_ASAP7_75t_R g7228 ( 
.A(n_6704),
.Y(n_7228)
);

CKINVDCx20_ASAP7_75t_R g7229 ( 
.A(n_6984),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_7001),
.Y(n_7230)
);

INVxp67_ASAP7_75t_L g7231 ( 
.A(n_6767),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_7003),
.Y(n_7232)
);

CKINVDCx20_ASAP7_75t_R g7233 ( 
.A(n_7009),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_7006),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_7012),
.Y(n_7235)
);

INVxp67_ASAP7_75t_L g7236 ( 
.A(n_6804),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_7014),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_7016),
.Y(n_7238)
);

CKINVDCx16_ASAP7_75t_R g7239 ( 
.A(n_6777),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7019),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_7022),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_7023),
.Y(n_7242)
);

INVxp67_ASAP7_75t_SL g7243 ( 
.A(n_6748),
.Y(n_7243)
);

CKINVDCx20_ASAP7_75t_R g7244 ( 
.A(n_7036),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_7025),
.Y(n_7245)
);

HB1xp67_ASAP7_75t_L g7246 ( 
.A(n_6866),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7026),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_7029),
.Y(n_7248)
);

CKINVDCx5p33_ASAP7_75t_R g7249 ( 
.A(n_6706),
.Y(n_7249)
);

CKINVDCx5p33_ASAP7_75t_R g7250 ( 
.A(n_6707),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_7031),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_7033),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_7035),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_7037),
.Y(n_7254)
);

CKINVDCx5p33_ASAP7_75t_R g7255 ( 
.A(n_6709),
.Y(n_7255)
);

INVxp67_ASAP7_75t_SL g7256 ( 
.A(n_6763),
.Y(n_7256)
);

CKINVDCx5p33_ASAP7_75t_R g7257 ( 
.A(n_6713),
.Y(n_7257)
);

CKINVDCx20_ASAP7_75t_R g7258 ( 
.A(n_7075),
.Y(n_7258)
);

INVx1_ASAP7_75t_L g7259 ( 
.A(n_7038),
.Y(n_7259)
);

CKINVDCx20_ASAP7_75t_R g7260 ( 
.A(n_6883),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7040),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7042),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7044),
.Y(n_7263)
);

CKINVDCx20_ASAP7_75t_R g7264 ( 
.A(n_6880),
.Y(n_7264)
);

INVxp33_ASAP7_75t_SL g7265 ( 
.A(n_6623),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7048),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_7050),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_7051),
.Y(n_7268)
);

INVxp67_ASAP7_75t_L g7269 ( 
.A(n_6851),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_6763),
.Y(n_7270)
);

CKINVDCx16_ASAP7_75t_R g7271 ( 
.A(n_6684),
.Y(n_7271)
);

CKINVDCx5p33_ASAP7_75t_R g7272 ( 
.A(n_6716),
.Y(n_7272)
);

CKINVDCx5p33_ASAP7_75t_R g7273 ( 
.A(n_6718),
.Y(n_7273)
);

CKINVDCx5p33_ASAP7_75t_R g7274 ( 
.A(n_6720),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_6763),
.Y(n_7275)
);

INVxp67_ASAP7_75t_SL g7276 ( 
.A(n_6810),
.Y(n_7276)
);

INVxp67_ASAP7_75t_SL g7277 ( 
.A(n_6810),
.Y(n_7277)
);

CKINVDCx5p33_ASAP7_75t_R g7278 ( 
.A(n_6721),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_6810),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_6896),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_6896),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_6896),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_6901),
.Y(n_7283)
);

CKINVDCx5p33_ASAP7_75t_R g7284 ( 
.A(n_6723),
.Y(n_7284)
);

INVxp33_ASAP7_75t_L g7285 ( 
.A(n_6919),
.Y(n_7285)
);

INVxp33_ASAP7_75t_L g7286 ( 
.A(n_6877),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6901),
.Y(n_7287)
);

INVx1_ASAP7_75t_L g7288 ( 
.A(n_6901),
.Y(n_7288)
);

CKINVDCx14_ASAP7_75t_R g7289 ( 
.A(n_6646),
.Y(n_7289)
);

CKINVDCx5p33_ASAP7_75t_R g7290 ( 
.A(n_6727),
.Y(n_7290)
);

INVx2_ASAP7_75t_L g7291 ( 
.A(n_7010),
.Y(n_7291)
);

HB1xp67_ASAP7_75t_L g7292 ( 
.A(n_6867),
.Y(n_7292)
);

INVx1_ASAP7_75t_L g7293 ( 
.A(n_7010),
.Y(n_7293)
);

CKINVDCx20_ASAP7_75t_R g7294 ( 
.A(n_6735),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7010),
.Y(n_7295)
);

INVx1_ASAP7_75t_L g7296 ( 
.A(n_6635),
.Y(n_7296)
);

INVxp67_ASAP7_75t_SL g7297 ( 
.A(n_6929),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6635),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6736),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_6736),
.Y(n_7300)
);

CKINVDCx5p33_ASAP7_75t_R g7301 ( 
.A(n_6737),
.Y(n_7301)
);

CKINVDCx5p33_ASAP7_75t_R g7302 ( 
.A(n_6740),
.Y(n_7302)
);

CKINVDCx16_ASAP7_75t_R g7303 ( 
.A(n_6879),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6936),
.Y(n_7304)
);

CKINVDCx5p33_ASAP7_75t_R g7305 ( 
.A(n_6742),
.Y(n_7305)
);

CKINVDCx5p33_ASAP7_75t_R g7306 ( 
.A(n_6744),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_6936),
.Y(n_7307)
);

CKINVDCx5p33_ASAP7_75t_R g7308 ( 
.A(n_6749),
.Y(n_7308)
);

CKINVDCx5p33_ASAP7_75t_R g7309 ( 
.A(n_6751),
.Y(n_7309)
);

CKINVDCx20_ASAP7_75t_R g7310 ( 
.A(n_6752),
.Y(n_7310)
);

CKINVDCx14_ASAP7_75t_R g7311 ( 
.A(n_6839),
.Y(n_7311)
);

INVxp33_ASAP7_75t_SL g7312 ( 
.A(n_6625),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6624),
.Y(n_7313)
);

INVx1_ASAP7_75t_L g7314 ( 
.A(n_6626),
.Y(n_7314)
);

CKINVDCx16_ASAP7_75t_R g7315 ( 
.A(n_6903),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_6627),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_6629),
.Y(n_7317)
);

INVx1_ASAP7_75t_L g7318 ( 
.A(n_6631),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_6633),
.Y(n_7319)
);

INVxp67_ASAP7_75t_SL g7320 ( 
.A(n_6873),
.Y(n_7320)
);

CKINVDCx5p33_ASAP7_75t_R g7321 ( 
.A(n_6755),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_6634),
.Y(n_7322)
);

BUFx3_ASAP7_75t_L g7323 ( 
.A(n_6909),
.Y(n_7323)
);

CKINVDCx20_ASAP7_75t_R g7324 ( 
.A(n_6764),
.Y(n_7324)
);

CKINVDCx5p33_ASAP7_75t_R g7325 ( 
.A(n_6772),
.Y(n_7325)
);

CKINVDCx5p33_ASAP7_75t_R g7326 ( 
.A(n_6773),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_6644),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_6649),
.Y(n_7328)
);

CKINVDCx20_ASAP7_75t_R g7329 ( 
.A(n_6774),
.Y(n_7329)
);

CKINVDCx5p33_ASAP7_75t_R g7330 ( 
.A(n_6778),
.Y(n_7330)
);

CKINVDCx20_ASAP7_75t_R g7331 ( 
.A(n_6781),
.Y(n_7331)
);

CKINVDCx20_ASAP7_75t_R g7332 ( 
.A(n_6787),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6650),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_6651),
.Y(n_7334)
);

CKINVDCx5p33_ASAP7_75t_R g7335 ( 
.A(n_6790),
.Y(n_7335)
);

CKINVDCx20_ASAP7_75t_R g7336 ( 
.A(n_6791),
.Y(n_7336)
);

INVx2_ASAP7_75t_L g7337 ( 
.A(n_6647),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_6653),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6663),
.Y(n_7339)
);

CKINVDCx5p33_ASAP7_75t_R g7340 ( 
.A(n_6795),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6654),
.Y(n_7341)
);

INVxp67_ASAP7_75t_SL g7342 ( 
.A(n_6992),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6656),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_6657),
.Y(n_7344)
);

INVxp67_ASAP7_75t_SL g7345 ( 
.A(n_7056),
.Y(n_7345)
);

HB1xp67_ASAP7_75t_L g7346 ( 
.A(n_6868),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_6658),
.Y(n_7347)
);

CKINVDCx5p33_ASAP7_75t_R g7348 ( 
.A(n_6796),
.Y(n_7348)
);

INVxp67_ASAP7_75t_SL g7349 ( 
.A(n_7057),
.Y(n_7349)
);

CKINVDCx5p33_ASAP7_75t_R g7350 ( 
.A(n_6800),
.Y(n_7350)
);

BUFx2_ASAP7_75t_L g7351 ( 
.A(n_6869),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6660),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_6662),
.Y(n_7353)
);

CKINVDCx5p33_ASAP7_75t_R g7354 ( 
.A(n_6801),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_6665),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_6672),
.Y(n_7356)
);

INVxp33_ASAP7_75t_L g7357 ( 
.A(n_6892),
.Y(n_7357)
);

CKINVDCx20_ASAP7_75t_R g7358 ( 
.A(n_6805),
.Y(n_7358)
);

INVxp67_ASAP7_75t_SL g7359 ( 
.A(n_7059),
.Y(n_7359)
);

CKINVDCx5p33_ASAP7_75t_R g7360 ( 
.A(n_6806),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6675),
.Y(n_7361)
);

INVxp67_ASAP7_75t_SL g7362 ( 
.A(n_7062),
.Y(n_7362)
);

CKINVDCx14_ASAP7_75t_R g7363 ( 
.A(n_6840),
.Y(n_7363)
);

CKINVDCx5p33_ASAP7_75t_R g7364 ( 
.A(n_6807),
.Y(n_7364)
);

CKINVDCx5p33_ASAP7_75t_R g7365 ( 
.A(n_6811),
.Y(n_7365)
);

CKINVDCx5p33_ASAP7_75t_R g7366 ( 
.A(n_6817),
.Y(n_7366)
);

INVx2_ASAP7_75t_L g7367 ( 
.A(n_6666),
.Y(n_7367)
);

BUFx3_ASAP7_75t_L g7368 ( 
.A(n_6909),
.Y(n_7368)
);

INVxp33_ASAP7_75t_L g7369 ( 
.A(n_6904),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_6679),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_6685),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_6687),
.Y(n_7372)
);

INVx1_ASAP7_75t_L g7373 ( 
.A(n_6698),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_6699),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6703),
.Y(n_7375)
);

INVxp67_ASAP7_75t_SL g7376 ( 
.A(n_7063),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_6705),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_6711),
.Y(n_7378)
);

CKINVDCx5p33_ASAP7_75t_R g7379 ( 
.A(n_6819),
.Y(n_7379)
);

CKINVDCx20_ASAP7_75t_R g7380 ( 
.A(n_6823),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_6715),
.Y(n_7381)
);

CKINVDCx5p33_ASAP7_75t_R g7382 ( 
.A(n_6824),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6719),
.Y(n_7383)
);

CKINVDCx20_ASAP7_75t_R g7384 ( 
.A(n_6825),
.Y(n_7384)
);

CKINVDCx5p33_ASAP7_75t_R g7385 ( 
.A(n_6828),
.Y(n_7385)
);

BUFx2_ASAP7_75t_L g7386 ( 
.A(n_6881),
.Y(n_7386)
);

CKINVDCx5p33_ASAP7_75t_R g7387 ( 
.A(n_6830),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_6722),
.Y(n_7388)
);

CKINVDCx20_ASAP7_75t_R g7389 ( 
.A(n_6832),
.Y(n_7389)
);

CKINVDCx20_ASAP7_75t_R g7390 ( 
.A(n_6833),
.Y(n_7390)
);

INVx2_ASAP7_75t_L g7391 ( 
.A(n_6688),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_6725),
.Y(n_7392)
);

CKINVDCx5p33_ASAP7_75t_R g7393 ( 
.A(n_6834),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_6726),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_6835),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_6730),
.Y(n_7396)
);

INVx1_ASAP7_75t_L g7397 ( 
.A(n_6732),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6733),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_6734),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6739),
.Y(n_7400)
);

INVx2_ASAP7_75t_L g7401 ( 
.A(n_6702),
.Y(n_7401)
);

CKINVDCx16_ASAP7_75t_R g7402 ( 
.A(n_7021),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_6750),
.Y(n_7403)
);

CKINVDCx16_ASAP7_75t_R g7404 ( 
.A(n_6655),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_6754),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_6756),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_6757),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_6758),
.Y(n_7408)
);

CKINVDCx20_ASAP7_75t_R g7409 ( 
.A(n_6836),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_6760),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6761),
.Y(n_7411)
);

INVxp67_ASAP7_75t_L g7412 ( 
.A(n_6898),
.Y(n_7412)
);

INVxp67_ASAP7_75t_SL g7413 ( 
.A(n_7066),
.Y(n_7413)
);

CKINVDCx16_ASAP7_75t_R g7414 ( 
.A(n_6714),
.Y(n_7414)
);

CKINVDCx16_ASAP7_75t_R g7415 ( 
.A(n_6753),
.Y(n_7415)
);

CKINVDCx5p33_ASAP7_75t_R g7416 ( 
.A(n_6838),
.Y(n_7416)
);

CKINVDCx5p33_ASAP7_75t_R g7417 ( 
.A(n_6888),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6765),
.Y(n_7418)
);

CKINVDCx5p33_ASAP7_75t_R g7419 ( 
.A(n_6889),
.Y(n_7419)
);

INVx1_ASAP7_75t_L g7420 ( 
.A(n_6770),
.Y(n_7420)
);

CKINVDCx5p33_ASAP7_75t_R g7421 ( 
.A(n_6890),
.Y(n_7421)
);

INVxp33_ASAP7_75t_SL g7422 ( 
.A(n_6628),
.Y(n_7422)
);

INVx2_ASAP7_75t_L g7423 ( 
.A(n_6724),
.Y(n_7423)
);

INVxp67_ASAP7_75t_L g7424 ( 
.A(n_6931),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_6771),
.Y(n_7425)
);

INVxp67_ASAP7_75t_SL g7426 ( 
.A(n_7067),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_6776),
.Y(n_7427)
);

BUFx3_ASAP7_75t_L g7428 ( 
.A(n_7015),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_6779),
.Y(n_7429)
);

INVx1_ASAP7_75t_L g7430 ( 
.A(n_6780),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_6782),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6784),
.Y(n_7432)
);

CKINVDCx20_ASAP7_75t_R g7433 ( 
.A(n_6861),
.Y(n_7433)
);

CKINVDCx20_ASAP7_75t_R g7434 ( 
.A(n_6862),
.Y(n_7434)
);

INVx1_ASAP7_75t_SL g7435 ( 
.A(n_7054),
.Y(n_7435)
);

INVxp33_ASAP7_75t_SL g7436 ( 
.A(n_6636),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_6785),
.Y(n_7437)
);

CKINVDCx5p33_ASAP7_75t_R g7438 ( 
.A(n_6893),
.Y(n_7438)
);

CKINVDCx20_ASAP7_75t_R g7439 ( 
.A(n_6894),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6786),
.Y(n_7440)
);

INVx2_ASAP7_75t_L g7441 ( 
.A(n_6729),
.Y(n_7441)
);

INVxp67_ASAP7_75t_SL g7442 ( 
.A(n_7068),
.Y(n_7442)
);

INVxp33_ASAP7_75t_SL g7443 ( 
.A(n_6637),
.Y(n_7443)
);

CKINVDCx20_ASAP7_75t_R g7444 ( 
.A(n_6895),
.Y(n_7444)
);

HB1xp67_ASAP7_75t_L g7445 ( 
.A(n_6897),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6789),
.Y(n_7446)
);

CKINVDCx5p33_ASAP7_75t_R g7447 ( 
.A(n_6900),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6792),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_6794),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6745),
.Y(n_7450)
);

INVxp67_ASAP7_75t_L g7451 ( 
.A(n_6769),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_6747),
.Y(n_7452)
);

CKINVDCx5p33_ASAP7_75t_R g7453 ( 
.A(n_6908),
.Y(n_7453)
);

INVxp67_ASAP7_75t_L g7454 ( 
.A(n_7058),
.Y(n_7454)
);

BUFx2_ASAP7_75t_L g7455 ( 
.A(n_6910),
.Y(n_7455)
);

CKINVDCx5p33_ASAP7_75t_R g7456 ( 
.A(n_6912),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_6768),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7015),
.Y(n_7458)
);

CKINVDCx5p33_ASAP7_75t_R g7459 ( 
.A(n_6913),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7041),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_7041),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_7070),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_7077),
.Y(n_7463)
);

CKINVDCx16_ASAP7_75t_R g7464 ( 
.A(n_6670),
.Y(n_7464)
);

CKINVDCx16_ASAP7_75t_R g7465 ( 
.A(n_6700),
.Y(n_7465)
);

CKINVDCx5p33_ASAP7_75t_R g7466 ( 
.A(n_6915),
.Y(n_7466)
);

BUFx3_ASAP7_75t_L g7467 ( 
.A(n_7079),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_7080),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7082),
.Y(n_7469)
);

CKINVDCx5p33_ASAP7_75t_R g7470 ( 
.A(n_6916),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_7083),
.Y(n_7471)
);

INVxp67_ASAP7_75t_L g7472 ( 
.A(n_6671),
.Y(n_7472)
);

CKINVDCx20_ASAP7_75t_R g7473 ( 
.A(n_6917),
.Y(n_7473)
);

CKINVDCx5p33_ASAP7_75t_R g7474 ( 
.A(n_6918),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7081),
.Y(n_7475)
);

INVxp67_ASAP7_75t_SL g7476 ( 
.A(n_6640),
.Y(n_7476)
);

CKINVDCx20_ASAP7_75t_R g7477 ( 
.A(n_6921),
.Y(n_7477)
);

CKINVDCx20_ASAP7_75t_R g7478 ( 
.A(n_6924),
.Y(n_7478)
);

CKINVDCx20_ASAP7_75t_R g7479 ( 
.A(n_6927),
.Y(n_7479)
);

BUFx2_ASAP7_75t_L g7480 ( 
.A(n_6934),
.Y(n_7480)
);

INVx1_ASAP7_75t_L g7481 ( 
.A(n_7053),
.Y(n_7481)
);

BUFx3_ASAP7_75t_L g7482 ( 
.A(n_6935),
.Y(n_7482)
);

INVx1_ASAP7_75t_L g7483 ( 
.A(n_6738),
.Y(n_7483)
);

CKINVDCx5p33_ASAP7_75t_R g7484 ( 
.A(n_6938),
.Y(n_7484)
);

CKINVDCx20_ASAP7_75t_R g7485 ( 
.A(n_6940),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_6738),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_6738),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_6738),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_6738),
.Y(n_7489)
);

HB1xp67_ASAP7_75t_L g7490 ( 
.A(n_6942),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_6759),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_6759),
.Y(n_7492)
);

CKINVDCx20_ASAP7_75t_R g7493 ( 
.A(n_6943),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6759),
.Y(n_7494)
);

INVxp67_ASAP7_75t_L g7495 ( 
.A(n_6695),
.Y(n_7495)
);

INVx1_ASAP7_75t_L g7496 ( 
.A(n_6759),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_6759),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7013),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_7013),
.Y(n_7499)
);

CKINVDCx5p33_ASAP7_75t_R g7500 ( 
.A(n_6947),
.Y(n_7500)
);

CKINVDCx5p33_ASAP7_75t_R g7501 ( 
.A(n_6955),
.Y(n_7501)
);

INVxp67_ASAP7_75t_L g7502 ( 
.A(n_6731),
.Y(n_7502)
);

INVx2_ASAP7_75t_L g7503 ( 
.A(n_7013),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_7013),
.Y(n_7504)
);

CKINVDCx5p33_ASAP7_75t_R g7505 ( 
.A(n_6956),
.Y(n_7505)
);

HB1xp67_ASAP7_75t_L g7506 ( 
.A(n_6958),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_7013),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_6664),
.Y(n_7508)
);

CKINVDCx16_ASAP7_75t_R g7509 ( 
.A(n_6712),
.Y(n_7509)
);

CKINVDCx5p33_ASAP7_75t_R g7510 ( 
.A(n_6960),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_6683),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_6961),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_6962),
.Y(n_7513)
);

CKINVDCx5p33_ASAP7_75t_R g7514 ( 
.A(n_6970),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_6973),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_6743),
.Y(n_7516)
);

CKINVDCx5p33_ASAP7_75t_R g7517 ( 
.A(n_6977),
.Y(n_7517)
);

CKINVDCx5p33_ASAP7_75t_R g7518 ( 
.A(n_6978),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_6979),
.Y(n_7519)
);

INVxp67_ASAP7_75t_SL g7520 ( 
.A(n_6885),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_6980),
.Y(n_7521)
);

INVx1_ASAP7_75t_L g7522 ( 
.A(n_6982),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_6983),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6986),
.Y(n_7524)
);

CKINVDCx20_ASAP7_75t_R g7525 ( 
.A(n_6988),
.Y(n_7525)
);

BUFx2_ASAP7_75t_L g7526 ( 
.A(n_6989),
.Y(n_7526)
);

CKINVDCx16_ASAP7_75t_R g7527 ( 
.A(n_6762),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_6990),
.Y(n_7528)
);

INVx1_ASAP7_75t_L g7529 ( 
.A(n_6993),
.Y(n_7529)
);

CKINVDCx20_ASAP7_75t_R g7530 ( 
.A(n_6997),
.Y(n_7530)
);

INVx2_ASAP7_75t_L g7531 ( 
.A(n_6793),
.Y(n_7531)
);

CKINVDCx5p33_ASAP7_75t_R g7532 ( 
.A(n_6998),
.Y(n_7532)
);

INVx2_ASAP7_75t_L g7533 ( 
.A(n_7002),
.Y(n_7533)
);

INVx1_ASAP7_75t_L g7534 ( 
.A(n_7004),
.Y(n_7534)
);

CKINVDCx5p33_ASAP7_75t_R g7535 ( 
.A(n_7005),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7007),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7011),
.Y(n_7537)
);

BUFx6f_ASAP7_75t_L g7538 ( 
.A(n_7018),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_7020),
.Y(n_7539)
);

CKINVDCx5p33_ASAP7_75t_R g7540 ( 
.A(n_7024),
.Y(n_7540)
);

CKINVDCx5p33_ASAP7_75t_R g7541 ( 
.A(n_7027),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7028),
.Y(n_7542)
);

HB1xp67_ASAP7_75t_L g7543 ( 
.A(n_7030),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7032),
.Y(n_7544)
);

CKINVDCx5p33_ASAP7_75t_R g7545 ( 
.A(n_7034),
.Y(n_7545)
);

INVx1_ASAP7_75t_L g7546 ( 
.A(n_7039),
.Y(n_7546)
);

CKINVDCx5p33_ASAP7_75t_R g7547 ( 
.A(n_7043),
.Y(n_7547)
);

CKINVDCx5p33_ASAP7_75t_R g7548 ( 
.A(n_7045),
.Y(n_7548)
);

CKINVDCx5p33_ASAP7_75t_R g7549 ( 
.A(n_7046),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7047),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7049),
.Y(n_7551)
);

INVxp67_ASAP7_75t_SL g7552 ( 
.A(n_6906),
.Y(n_7552)
);

INVx1_ASAP7_75t_L g7553 ( 
.A(n_7052),
.Y(n_7553)
);

INVx1_ASAP7_75t_L g7554 ( 
.A(n_7055),
.Y(n_7554)
);

INVxp67_ASAP7_75t_SL g7555 ( 
.A(n_7078),
.Y(n_7555)
);

CKINVDCx5p33_ASAP7_75t_R g7556 ( 
.A(n_7060),
.Y(n_7556)
);

CKINVDCx5p33_ASAP7_75t_R g7557 ( 
.A(n_7061),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7064),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_7065),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7069),
.Y(n_7560)
);

INVxp67_ASAP7_75t_SL g7561 ( 
.A(n_6681),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_7071),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_7072),
.Y(n_7563)
);

INVx1_ASAP7_75t_L g7564 ( 
.A(n_7073),
.Y(n_7564)
);

INVx1_ASAP7_75t_L g7565 ( 
.A(n_7074),
.Y(n_7565)
);

INVx1_ASAP7_75t_L g7566 ( 
.A(n_6902),
.Y(n_7566)
);

CKINVDCx20_ASAP7_75t_R g7567 ( 
.A(n_6845),
.Y(n_7567)
);

BUFx3_ASAP7_75t_L g7568 ( 
.A(n_6976),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_6999),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_7076),
.Y(n_7570)
);

CKINVDCx5p33_ASAP7_75t_R g7571 ( 
.A(n_6638),
.Y(n_7571)
);

INVxp67_ASAP7_75t_SL g7572 ( 
.A(n_6964),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7017),
.Y(n_7573)
);

CKINVDCx20_ASAP7_75t_R g7574 ( 
.A(n_6639),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_6630),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_6746),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_6746),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6827),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_6827),
.Y(n_7579)
);

CKINVDCx5p33_ASAP7_75t_R g7580 ( 
.A(n_6641),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_6798),
.Y(n_7581)
);

CKINVDCx5p33_ASAP7_75t_R g7582 ( 
.A(n_6642),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_6841),
.Y(n_7583)
);

INVxp33_ASAP7_75t_L g7584 ( 
.A(n_6831),
.Y(n_7584)
);

CKINVDCx5p33_ASAP7_75t_R g7585 ( 
.A(n_6643),
.Y(n_7585)
);

INVx1_ASAP7_75t_L g7586 ( 
.A(n_6803),
.Y(n_7586)
);

INVxp67_ASAP7_75t_SL g7587 ( 
.A(n_6865),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_6803),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_6803),
.Y(n_7589)
);

CKINVDCx16_ASAP7_75t_R g7590 ( 
.A(n_6788),
.Y(n_7590)
);

CKINVDCx20_ASAP7_75t_R g7591 ( 
.A(n_6632),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_6803),
.Y(n_7592)
);

CKINVDCx20_ASAP7_75t_R g7593 ( 
.A(n_6632),
.Y(n_7593)
);

CKINVDCx5p33_ASAP7_75t_R g7594 ( 
.A(n_6643),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_6803),
.Y(n_7595)
);

CKINVDCx16_ASAP7_75t_R g7596 ( 
.A(n_6788),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_6803),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_6803),
.Y(n_7598)
);

CKINVDCx5p33_ASAP7_75t_R g7599 ( 
.A(n_6643),
.Y(n_7599)
);

CKINVDCx5p33_ASAP7_75t_R g7600 ( 
.A(n_6643),
.Y(n_7600)
);

INVxp67_ASAP7_75t_SL g7601 ( 
.A(n_6865),
.Y(n_7601)
);

CKINVDCx5p33_ASAP7_75t_R g7602 ( 
.A(n_6643),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_6803),
.Y(n_7603)
);

HB1xp67_ASAP7_75t_L g7604 ( 
.A(n_6853),
.Y(n_7604)
);

CKINVDCx20_ASAP7_75t_R g7605 ( 
.A(n_6632),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_6803),
.Y(n_7606)
);

CKINVDCx5p33_ASAP7_75t_R g7607 ( 
.A(n_6643),
.Y(n_7607)
);

CKINVDCx20_ASAP7_75t_R g7608 ( 
.A(n_6632),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_6803),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_6803),
.Y(n_7610)
);

CKINVDCx5p33_ASAP7_75t_R g7611 ( 
.A(n_6643),
.Y(n_7611)
);

INVx3_ASAP7_75t_L g7612 ( 
.A(n_7194),
.Y(n_7612)
);

OAI21xp33_ASAP7_75t_L g7613 ( 
.A1(n_7516),
.A2(n_5222),
.B(n_5186),
.Y(n_7613)
);

AOI22xp5_ASAP7_75t_L g7614 ( 
.A1(n_7187),
.A2(n_5486),
.B1(n_5624),
.B2(n_5185),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_SL g7615 ( 
.A(n_7572),
.B(n_5405),
.Y(n_7615)
);

BUFx6f_ASAP7_75t_L g7616 ( 
.A(n_7194),
.Y(n_7616)
);

AND2x6_ASAP7_75t_L g7617 ( 
.A(n_7538),
.B(n_6162),
.Y(n_7617)
);

INVx5_ASAP7_75t_L g7618 ( 
.A(n_7143),
.Y(n_7618)
);

BUFx6f_ASAP7_75t_L g7619 ( 
.A(n_7194),
.Y(n_7619)
);

CKINVDCx5p33_ASAP7_75t_R g7620 ( 
.A(n_7095),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7313),
.Y(n_7621)
);

AND2x2_ASAP7_75t_L g7622 ( 
.A(n_7285),
.B(n_5331),
.Y(n_7622)
);

NOR2xp33_ASAP7_75t_L g7623 ( 
.A(n_7191),
.B(n_5517),
.Y(n_7623)
);

OAI22xp5_ASAP7_75t_L g7624 ( 
.A1(n_7320),
.A2(n_5744),
.B1(n_5802),
.B2(n_5732),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7314),
.Y(n_7625)
);

OAI22x1_ASAP7_75t_SL g7626 ( 
.A1(n_7433),
.A2(n_5436),
.B1(n_5446),
.B2(n_5392),
.Y(n_7626)
);

INVx2_ASAP7_75t_SL g7627 ( 
.A(n_7573),
.Y(n_7627)
);

AOI22xp5_ASAP7_75t_L g7628 ( 
.A1(n_7561),
.A2(n_5702),
.B1(n_5840),
.B2(n_5700),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7316),
.Y(n_7629)
);

BUFx6f_ASAP7_75t_L g7630 ( 
.A(n_7198),
.Y(n_7630)
);

BUFx2_ASAP7_75t_L g7631 ( 
.A(n_7464),
.Y(n_7631)
);

NAND2xp5_ASAP7_75t_L g7632 ( 
.A(n_7342),
.B(n_5549),
.Y(n_7632)
);

INVx1_ASAP7_75t_L g7633 ( 
.A(n_7317),
.Y(n_7633)
);

INVx2_ASAP7_75t_L g7634 ( 
.A(n_7121),
.Y(n_7634)
);

INVx2_ASAP7_75t_SL g7635 ( 
.A(n_7105),
.Y(n_7635)
);

BUFx6f_ASAP7_75t_L g7636 ( 
.A(n_7085),
.Y(n_7636)
);

AND2x4_ASAP7_75t_L g7637 ( 
.A(n_7205),
.B(n_6178),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7318),
.Y(n_7638)
);

AOI22xp5_ASAP7_75t_L g7639 ( 
.A1(n_7297),
.A2(n_5809),
.B1(n_6166),
.B2(n_5770),
.Y(n_7639)
);

OAI22xp5_ASAP7_75t_L g7640 ( 
.A1(n_7531),
.A2(n_6506),
.B1(n_6081),
.B2(n_5333),
.Y(n_7640)
);

BUFx6f_ASAP7_75t_L g7641 ( 
.A(n_7085),
.Y(n_7641)
);

OAI21x1_ASAP7_75t_L g7642 ( 
.A1(n_7483),
.A2(n_5512),
.B(n_5365),
.Y(n_7642)
);

BUFx12f_ASAP7_75t_L g7643 ( 
.A(n_7417),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_7134),
.Y(n_7644)
);

INVx2_ASAP7_75t_L g7645 ( 
.A(n_7142),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7319),
.Y(n_7646)
);

AOI22x1_ASAP7_75t_SL g7647 ( 
.A1(n_7264),
.A2(n_5469),
.B1(n_5479),
.B2(n_5461),
.Y(n_7647)
);

BUFx12f_ASAP7_75t_L g7648 ( 
.A(n_7419),
.Y(n_7648)
);

INVx5_ASAP7_75t_L g7649 ( 
.A(n_7178),
.Y(n_7649)
);

INVx4_ASAP7_75t_L g7650 ( 
.A(n_7538),
.Y(n_7650)
);

AND2x4_ASAP7_75t_L g7651 ( 
.A(n_7221),
.B(n_6211),
.Y(n_7651)
);

INVx1_ASAP7_75t_L g7652 ( 
.A(n_7322),
.Y(n_7652)
);

AND2x4_ASAP7_75t_L g7653 ( 
.A(n_7481),
.B(n_6239),
.Y(n_7653)
);

BUFx2_ASAP7_75t_L g7654 ( 
.A(n_7465),
.Y(n_7654)
);

OAI21x1_ASAP7_75t_L g7655 ( 
.A1(n_7486),
.A2(n_5657),
.B(n_5253),
.Y(n_7655)
);

INVx1_ASAP7_75t_L g7656 ( 
.A(n_7327),
.Y(n_7656)
);

NOR2xp33_ASAP7_75t_L g7657 ( 
.A(n_7106),
.B(n_6251),
.Y(n_7657)
);

INVx2_ASAP7_75t_L g7658 ( 
.A(n_7145),
.Y(n_7658)
);

BUFx6f_ASAP7_75t_L g7659 ( 
.A(n_7157),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7328),
.Y(n_7660)
);

AOI22xp5_ASAP7_75t_L g7661 ( 
.A1(n_7512),
.A2(n_6362),
.B1(n_5285),
.B2(n_5422),
.Y(n_7661)
);

AND2x4_ASAP7_75t_L g7662 ( 
.A(n_7587),
.B(n_6282),
.Y(n_7662)
);

BUFx3_ASAP7_75t_L g7663 ( 
.A(n_7467),
.Y(n_7663)
);

OAI22xp5_ASAP7_75t_L g7664 ( 
.A1(n_7513),
.A2(n_5334),
.B1(n_5335),
.B2(n_5332),
.Y(n_7664)
);

AND2x6_ASAP7_75t_L g7665 ( 
.A(n_7538),
.B(n_6311),
.Y(n_7665)
);

AND2x2_ASAP7_75t_L g7666 ( 
.A(n_7584),
.B(n_5353),
.Y(n_7666)
);

OA21x2_ASAP7_75t_L g7667 ( 
.A1(n_7487),
.A2(n_5310),
.B(n_5244),
.Y(n_7667)
);

OAI22xp5_ASAP7_75t_L g7668 ( 
.A1(n_7515),
.A2(n_5338),
.B1(n_5339),
.B2(n_5336),
.Y(n_7668)
);

CKINVDCx11_ASAP7_75t_R g7669 ( 
.A(n_7146),
.Y(n_7669)
);

NAND2xp5_ASAP7_75t_L g7670 ( 
.A(n_7601),
.B(n_6616),
.Y(n_7670)
);

BUFx6f_ASAP7_75t_L g7671 ( 
.A(n_7167),
.Y(n_7671)
);

INVx2_ASAP7_75t_L g7672 ( 
.A(n_7171),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7333),
.Y(n_7673)
);

OAI21x1_ASAP7_75t_L g7674 ( 
.A1(n_7489),
.A2(n_5429),
.B(n_5342),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7216),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7334),
.Y(n_7676)
);

AND2x2_ASAP7_75t_L g7677 ( 
.A(n_7520),
.B(n_5353),
.Y(n_7677)
);

BUFx8_ASAP7_75t_L g7678 ( 
.A(n_7120),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7476),
.B(n_5606),
.Y(n_7679)
);

INVx2_ASAP7_75t_L g7680 ( 
.A(n_7280),
.Y(n_7680)
);

AND2x4_ASAP7_75t_L g7681 ( 
.A(n_7323),
.B(n_6318),
.Y(n_7681)
);

OAI22xp5_ASAP7_75t_L g7682 ( 
.A1(n_7519),
.A2(n_5341),
.B1(n_5343),
.B2(n_5340),
.Y(n_7682)
);

BUFx2_ASAP7_75t_L g7683 ( 
.A(n_7509),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_7338),
.Y(n_7684)
);

BUFx6f_ASAP7_75t_L g7685 ( 
.A(n_7291),
.Y(n_7685)
);

AND2x4_ASAP7_75t_L g7686 ( 
.A(n_7368),
.B(n_6330),
.Y(n_7686)
);

INVx5_ASAP7_75t_L g7687 ( 
.A(n_7193),
.Y(n_7687)
);

AND2x4_ASAP7_75t_L g7688 ( 
.A(n_7428),
.B(n_6418),
.Y(n_7688)
);

BUFx6f_ASAP7_75t_L g7689 ( 
.A(n_7270),
.Y(n_7689)
);

BUFx8_ASAP7_75t_SL g7690 ( 
.A(n_7260),
.Y(n_7690)
);

AND2x2_ASAP7_75t_L g7691 ( 
.A(n_7435),
.B(n_5354),
.Y(n_7691)
);

BUFx12f_ASAP7_75t_L g7692 ( 
.A(n_7421),
.Y(n_7692)
);

INVx3_ASAP7_75t_L g7693 ( 
.A(n_7337),
.Y(n_7693)
);

BUFx6f_ASAP7_75t_L g7694 ( 
.A(n_7275),
.Y(n_7694)
);

BUFx3_ASAP7_75t_L g7695 ( 
.A(n_7294),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7341),
.Y(n_7696)
);

BUFx6f_ASAP7_75t_L g7697 ( 
.A(n_7279),
.Y(n_7697)
);

AND2x2_ASAP7_75t_L g7698 ( 
.A(n_7286),
.B(n_5354),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7343),
.Y(n_7699)
);

INVxp67_ASAP7_75t_L g7700 ( 
.A(n_7552),
.Y(n_7700)
);

AND2x4_ASAP7_75t_L g7701 ( 
.A(n_7533),
.B(n_7560),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7093),
.Y(n_7702)
);

BUFx2_ASAP7_75t_L g7703 ( 
.A(n_7527),
.Y(n_7703)
);

NAND2xp5_ASAP7_75t_SL g7704 ( 
.A(n_7271),
.B(n_5348),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7344),
.Y(n_7705)
);

INVx3_ASAP7_75t_L g7706 ( 
.A(n_7339),
.Y(n_7706)
);

BUFx3_ASAP7_75t_L g7707 ( 
.A(n_7310),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_7347),
.Y(n_7708)
);

AND2x4_ASAP7_75t_L g7709 ( 
.A(n_7508),
.B(n_6457),
.Y(n_7709)
);

AND2x2_ASAP7_75t_L g7710 ( 
.A(n_7357),
.B(n_5368),
.Y(n_7710)
);

INVx1_ASAP7_75t_L g7711 ( 
.A(n_7352),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7353),
.Y(n_7712)
);

AND2x2_ASAP7_75t_L g7713 ( 
.A(n_7369),
.B(n_5368),
.Y(n_7713)
);

AND2x4_ASAP7_75t_L g7714 ( 
.A(n_7511),
.B(n_6480),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_7355),
.Y(n_7715)
);

OA21x2_ASAP7_75t_L g7716 ( 
.A1(n_7491),
.A2(n_5755),
.B(n_5696),
.Y(n_7716)
);

AND2x2_ASAP7_75t_L g7717 ( 
.A(n_7147),
.B(n_5426),
.Y(n_7717)
);

INVx3_ASAP7_75t_L g7718 ( 
.A(n_7367),
.Y(n_7718)
);

BUFx6f_ASAP7_75t_L g7719 ( 
.A(n_7281),
.Y(n_7719)
);

INVx1_ASAP7_75t_L g7720 ( 
.A(n_7356),
.Y(n_7720)
);

INVx2_ASAP7_75t_L g7721 ( 
.A(n_7391),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_7361),
.Y(n_7722)
);

BUFx12f_ASAP7_75t_L g7723 ( 
.A(n_7438),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7370),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_7371),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_7401),
.Y(n_7726)
);

BUFx6f_ASAP7_75t_L g7727 ( 
.A(n_7282),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7372),
.Y(n_7728)
);

BUFx8_ASAP7_75t_L g7729 ( 
.A(n_7351),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7227),
.B(n_5762),
.Y(n_7730)
);

BUFx6f_ASAP7_75t_L g7731 ( 
.A(n_7283),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7373),
.Y(n_7732)
);

NAND2xp5_ASAP7_75t_L g7733 ( 
.A(n_7243),
.B(n_5773),
.Y(n_7733)
);

BUFx2_ASAP7_75t_L g7734 ( 
.A(n_7434),
.Y(n_7734)
);

BUFx3_ASAP7_75t_L g7735 ( 
.A(n_7324),
.Y(n_7735)
);

BUFx6f_ASAP7_75t_L g7736 ( 
.A(n_7287),
.Y(n_7736)
);

NAND2xp5_ASAP7_75t_L g7737 ( 
.A(n_7256),
.B(n_5778),
.Y(n_7737)
);

INVx2_ASAP7_75t_L g7738 ( 
.A(n_7423),
.Y(n_7738)
);

BUFx3_ASAP7_75t_L g7739 ( 
.A(n_7329),
.Y(n_7739)
);

OAI22xp5_ASAP7_75t_L g7740 ( 
.A1(n_7521),
.A2(n_5350),
.B1(n_5352),
.B2(n_5349),
.Y(n_7740)
);

BUFx12f_ASAP7_75t_L g7741 ( 
.A(n_7447),
.Y(n_7741)
);

CKINVDCx5p33_ASAP7_75t_R g7742 ( 
.A(n_7107),
.Y(n_7742)
);

INVx2_ASAP7_75t_L g7743 ( 
.A(n_7441),
.Y(n_7743)
);

BUFx6f_ASAP7_75t_L g7744 ( 
.A(n_7288),
.Y(n_7744)
);

INVx2_ASAP7_75t_L g7745 ( 
.A(n_7293),
.Y(n_7745)
);

INVx5_ASAP7_75t_L g7746 ( 
.A(n_7214),
.Y(n_7746)
);

AOI22xp5_ASAP7_75t_L g7747 ( 
.A1(n_7522),
.A2(n_5438),
.B1(n_5482),
.B2(n_5259),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7374),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7375),
.Y(n_7749)
);

INVx2_ASAP7_75t_L g7750 ( 
.A(n_7295),
.Y(n_7750)
);

BUFx2_ASAP7_75t_L g7751 ( 
.A(n_7472),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7377),
.Y(n_7752)
);

AND2x2_ASAP7_75t_SL g7753 ( 
.A(n_7239),
.B(n_5195),
.Y(n_7753)
);

NOR2xp33_ASAP7_75t_L g7754 ( 
.A(n_7523),
.B(n_5194),
.Y(n_7754)
);

BUFx3_ASAP7_75t_L g7755 ( 
.A(n_7331),
.Y(n_7755)
);

OAI22x1_ASAP7_75t_SL g7756 ( 
.A1(n_7153),
.A2(n_5490),
.B1(n_5556),
.B2(n_5484),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7378),
.Y(n_7757)
);

AND2x6_ASAP7_75t_L g7758 ( 
.A(n_7524),
.B(n_7528),
.Y(n_7758)
);

INVx4_ASAP7_75t_L g7759 ( 
.A(n_7111),
.Y(n_7759)
);

BUFx6f_ASAP7_75t_L g7760 ( 
.A(n_7450),
.Y(n_7760)
);

CKINVDCx20_ASAP7_75t_R g7761 ( 
.A(n_7084),
.Y(n_7761)
);

BUFx2_ASAP7_75t_L g7762 ( 
.A(n_7495),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_7381),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7383),
.Y(n_7764)
);

AND2x2_ASAP7_75t_L g7765 ( 
.A(n_7555),
.B(n_5426),
.Y(n_7765)
);

OAI22x1_ASAP7_75t_L g7766 ( 
.A1(n_7502),
.A2(n_5568),
.B1(n_5529),
.B2(n_5530),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_L g7767 ( 
.A(n_7276),
.B(n_5863),
.Y(n_7767)
);

AND2x4_ASAP7_75t_L g7768 ( 
.A(n_7458),
.B(n_7460),
.Y(n_7768)
);

AND2x4_ASAP7_75t_L g7769 ( 
.A(n_7461),
.B(n_6521),
.Y(n_7769)
);

AND2x2_ASAP7_75t_L g7770 ( 
.A(n_7386),
.B(n_5502),
.Y(n_7770)
);

OA21x2_ASAP7_75t_L g7771 ( 
.A1(n_7492),
.A2(n_6099),
.B(n_6036),
.Y(n_7771)
);

BUFx3_ASAP7_75t_L g7772 ( 
.A(n_7332),
.Y(n_7772)
);

BUFx2_ASAP7_75t_L g7773 ( 
.A(n_7439),
.Y(n_7773)
);

OAI21x1_ASAP7_75t_L g7774 ( 
.A1(n_7494),
.A2(n_6283),
.B(n_6215),
.Y(n_7774)
);

CKINVDCx20_ASAP7_75t_R g7775 ( 
.A(n_7097),
.Y(n_7775)
);

BUFx8_ASAP7_75t_L g7776 ( 
.A(n_7455),
.Y(n_7776)
);

BUFx6f_ASAP7_75t_L g7777 ( 
.A(n_7452),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7388),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7392),
.Y(n_7779)
);

INVx2_ASAP7_75t_L g7780 ( 
.A(n_7457),
.Y(n_7780)
);

INVx2_ASAP7_75t_L g7781 ( 
.A(n_7104),
.Y(n_7781)
);

AOI22xp33_ASAP7_75t_L g7782 ( 
.A1(n_7394),
.A2(n_5267),
.B1(n_5287),
.B2(n_5214),
.Y(n_7782)
);

OA21x2_ASAP7_75t_L g7783 ( 
.A1(n_7496),
.A2(n_6322),
.B(n_6320),
.Y(n_7783)
);

NOR2xp33_ASAP7_75t_L g7784 ( 
.A(n_7529),
.B(n_5229),
.Y(n_7784)
);

NAND2xp5_ASAP7_75t_L g7785 ( 
.A(n_7277),
.B(n_6396),
.Y(n_7785)
);

AND2x4_ASAP7_75t_L g7786 ( 
.A(n_7534),
.B(n_6526),
.Y(n_7786)
);

CKINVDCx5p33_ASAP7_75t_R g7787 ( 
.A(n_7123),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7396),
.Y(n_7788)
);

INVx6_ASAP7_75t_L g7789 ( 
.A(n_7303),
.Y(n_7789)
);

NAND2xp5_ASAP7_75t_L g7790 ( 
.A(n_7397),
.B(n_6432),
.Y(n_7790)
);

BUFx6f_ASAP7_75t_L g7791 ( 
.A(n_7296),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7398),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_7399),
.Y(n_7793)
);

INVxp67_ASAP7_75t_L g7794 ( 
.A(n_7581),
.Y(n_7794)
);

BUFx12f_ASAP7_75t_L g7795 ( 
.A(n_7453),
.Y(n_7795)
);

NAND2xp5_ASAP7_75t_L g7796 ( 
.A(n_7400),
.B(n_6528),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_L g7797 ( 
.A(n_7403),
.B(n_6621),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7405),
.Y(n_7798)
);

INVx2_ASAP7_75t_L g7799 ( 
.A(n_7108),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_7406),
.Y(n_7800)
);

AND2x2_ASAP7_75t_L g7801 ( 
.A(n_7480),
.B(n_7526),
.Y(n_7801)
);

OA21x2_ASAP7_75t_L g7802 ( 
.A1(n_7497),
.A2(n_5180),
.B(n_5176),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_7109),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7407),
.Y(n_7804)
);

AND2x4_ASAP7_75t_L g7805 ( 
.A(n_7536),
.B(n_6535),
.Y(n_7805)
);

OAI21x1_ASAP7_75t_L g7806 ( 
.A1(n_7498),
.A2(n_5351),
.B(n_5307),
.Y(n_7806)
);

OAI21x1_ASAP7_75t_L g7807 ( 
.A1(n_7499),
.A2(n_5398),
.B(n_5374),
.Y(n_7807)
);

AND2x2_ASAP7_75t_SL g7808 ( 
.A(n_7404),
.B(n_7414),
.Y(n_7808)
);

OAI22x1_ASAP7_75t_L g7809 ( 
.A1(n_7087),
.A2(n_5599),
.B1(n_5618),
.B2(n_5505),
.Y(n_7809)
);

NAND2xp5_ASAP7_75t_L g7810 ( 
.A(n_7408),
.B(n_5179),
.Y(n_7810)
);

INVx2_ASAP7_75t_L g7811 ( 
.A(n_7110),
.Y(n_7811)
);

INVx2_ASAP7_75t_L g7812 ( 
.A(n_7114),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7410),
.Y(n_7813)
);

INVx5_ASAP7_75t_L g7814 ( 
.A(n_7162),
.Y(n_7814)
);

INVx2_ASAP7_75t_L g7815 ( 
.A(n_7115),
.Y(n_7815)
);

INVx2_ASAP7_75t_L g7816 ( 
.A(n_7117),
.Y(n_7816)
);

INVx4_ASAP7_75t_L g7817 ( 
.A(n_7130),
.Y(n_7817)
);

INVx2_ASAP7_75t_L g7818 ( 
.A(n_7118),
.Y(n_7818)
);

NAND2xp5_ASAP7_75t_L g7819 ( 
.A(n_7411),
.B(n_5179),
.Y(n_7819)
);

INVx6_ASAP7_75t_L g7820 ( 
.A(n_7315),
.Y(n_7820)
);

HB1xp67_ASAP7_75t_L g7821 ( 
.A(n_7099),
.Y(n_7821)
);

BUFx6f_ASAP7_75t_L g7822 ( 
.A(n_7298),
.Y(n_7822)
);

BUFx6f_ASAP7_75t_L g7823 ( 
.A(n_7299),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_7418),
.Y(n_7824)
);

NAND2xp5_ASAP7_75t_L g7825 ( 
.A(n_7420),
.B(n_5179),
.Y(n_7825)
);

BUFx8_ASAP7_75t_L g7826 ( 
.A(n_7575),
.Y(n_7826)
);

AND2x2_ASAP7_75t_L g7827 ( 
.A(n_7182),
.B(n_5502),
.Y(n_7827)
);

HB1xp67_ASAP7_75t_L g7828 ( 
.A(n_7122),
.Y(n_7828)
);

BUFx12f_ASAP7_75t_L g7829 ( 
.A(n_7456),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7425),
.Y(n_7830)
);

INVx2_ASAP7_75t_L g7831 ( 
.A(n_7119),
.Y(n_7831)
);

BUFx6f_ASAP7_75t_L g7832 ( 
.A(n_7300),
.Y(n_7832)
);

BUFx6f_ASAP7_75t_L g7833 ( 
.A(n_7304),
.Y(n_7833)
);

INVx2_ASAP7_75t_L g7834 ( 
.A(n_7127),
.Y(n_7834)
);

NAND2xp5_ASAP7_75t_L g7835 ( 
.A(n_7427),
.B(n_5179),
.Y(n_7835)
);

INVx2_ASAP7_75t_L g7836 ( 
.A(n_7131),
.Y(n_7836)
);

INVx4_ASAP7_75t_L g7837 ( 
.A(n_7136),
.Y(n_7837)
);

AND2x2_ASAP7_75t_L g7838 ( 
.A(n_7213),
.B(n_5520),
.Y(n_7838)
);

INVx2_ASAP7_75t_L g7839 ( 
.A(n_7133),
.Y(n_7839)
);

HB1xp67_ASAP7_75t_L g7840 ( 
.A(n_7126),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_7462),
.Y(n_7841)
);

CKINVDCx5p33_ASAP7_75t_R g7842 ( 
.A(n_7149),
.Y(n_7842)
);

BUFx6f_ASAP7_75t_L g7843 ( 
.A(n_7307),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_7463),
.Y(n_7844)
);

CKINVDCx20_ASAP7_75t_R g7845 ( 
.A(n_7112),
.Y(n_7845)
);

AND2x4_ASAP7_75t_L g7846 ( 
.A(n_7537),
.B(n_6547),
.Y(n_7846)
);

CKINVDCx5p33_ASAP7_75t_R g7847 ( 
.A(n_7159),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7135),
.Y(n_7848)
);

BUFx6f_ASAP7_75t_L g7849 ( 
.A(n_7137),
.Y(n_7849)
);

INVx2_ASAP7_75t_L g7850 ( 
.A(n_7138),
.Y(n_7850)
);

CKINVDCx5p33_ASAP7_75t_R g7851 ( 
.A(n_7161),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_L g7852 ( 
.A(n_7475),
.B(n_5269),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7468),
.Y(n_7853)
);

OAI22x1_ASAP7_75t_R g7854 ( 
.A1(n_7574),
.A2(n_5591),
.B1(n_5648),
.B2(n_5558),
.Y(n_7854)
);

INVx1_ASAP7_75t_L g7855 ( 
.A(n_7469),
.Y(n_7855)
);

INVx2_ASAP7_75t_L g7856 ( 
.A(n_7139),
.Y(n_7856)
);

BUFx3_ASAP7_75t_L g7857 ( 
.A(n_7336),
.Y(n_7857)
);

OAI22xp5_ASAP7_75t_L g7858 ( 
.A1(n_7539),
.A2(n_5355),
.B1(n_5358),
.B2(n_5357),
.Y(n_7858)
);

NAND2xp5_ASAP7_75t_L g7859 ( 
.A(n_7504),
.B(n_7507),
.Y(n_7859)
);

INVx2_ASAP7_75t_L g7860 ( 
.A(n_7140),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7471),
.Y(n_7861)
);

BUFx6f_ASAP7_75t_L g7862 ( 
.A(n_7141),
.Y(n_7862)
);

INVx2_ASAP7_75t_L g7863 ( 
.A(n_7144),
.Y(n_7863)
);

BUFx6f_ASAP7_75t_L g7864 ( 
.A(n_7148),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7429),
.Y(n_7865)
);

AND2x6_ASAP7_75t_L g7866 ( 
.A(n_7542),
.B(n_6556),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7430),
.Y(n_7867)
);

BUFx2_ASAP7_75t_L g7868 ( 
.A(n_7444),
.Y(n_7868)
);

AND2x4_ASAP7_75t_L g7869 ( 
.A(n_7544),
.B(n_5321),
.Y(n_7869)
);

OA21x2_ASAP7_75t_L g7870 ( 
.A1(n_7488),
.A2(n_5188),
.B(n_5182),
.Y(n_7870)
);

BUFx6f_ASAP7_75t_L g7871 ( 
.A(n_7150),
.Y(n_7871)
);

AND2x4_ASAP7_75t_L g7872 ( 
.A(n_7546),
.B(n_5419),
.Y(n_7872)
);

INVx2_ASAP7_75t_L g7873 ( 
.A(n_7151),
.Y(n_7873)
);

INVx6_ASAP7_75t_L g7874 ( 
.A(n_7402),
.Y(n_7874)
);

AND2x6_ASAP7_75t_L g7875 ( 
.A(n_7550),
.B(n_5632),
.Y(n_7875)
);

INVx3_ASAP7_75t_L g7876 ( 
.A(n_7431),
.Y(n_7876)
);

OA21x2_ASAP7_75t_L g7877 ( 
.A1(n_7503),
.A2(n_5209),
.B(n_5202),
.Y(n_7877)
);

BUFx8_ASAP7_75t_SL g7878 ( 
.A(n_7156),
.Y(n_7878)
);

HB1xp67_ASAP7_75t_L g7879 ( 
.A(n_7160),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_7432),
.Y(n_7880)
);

BUFx3_ASAP7_75t_L g7881 ( 
.A(n_7358),
.Y(n_7881)
);

BUFx6f_ASAP7_75t_L g7882 ( 
.A(n_7154),
.Y(n_7882)
);

BUFx6f_ASAP7_75t_L g7883 ( 
.A(n_7155),
.Y(n_7883)
);

INVx2_ASAP7_75t_L g7884 ( 
.A(n_7158),
.Y(n_7884)
);

INVx4_ASAP7_75t_L g7885 ( 
.A(n_7164),
.Y(n_7885)
);

INVx1_ASAP7_75t_L g7886 ( 
.A(n_7437),
.Y(n_7886)
);

AND2x2_ASAP7_75t_L g7887 ( 
.A(n_7222),
.B(n_5520),
.Y(n_7887)
);

NAND2xp5_ASAP7_75t_L g7888 ( 
.A(n_7345),
.B(n_5468),
.Y(n_7888)
);

INVx1_ASAP7_75t_L g7889 ( 
.A(n_7440),
.Y(n_7889)
);

INVx1_ASAP7_75t_L g7890 ( 
.A(n_7446),
.Y(n_7890)
);

AND2x6_ASAP7_75t_L g7891 ( 
.A(n_7551),
.B(n_5634),
.Y(n_7891)
);

NAND2xp5_ASAP7_75t_L g7892 ( 
.A(n_7349),
.B(n_5637),
.Y(n_7892)
);

BUFx12f_ASAP7_75t_L g7893 ( 
.A(n_7459),
.Y(n_7893)
);

NOR2xp33_ASAP7_75t_L g7894 ( 
.A(n_7553),
.B(n_5678),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7359),
.B(n_5777),
.Y(n_7895)
);

NOR2xp33_ASAP7_75t_L g7896 ( 
.A(n_7554),
.B(n_5992),
.Y(n_7896)
);

OA21x2_ASAP7_75t_L g7897 ( 
.A1(n_7566),
.A2(n_5216),
.B(n_5215),
.Y(n_7897)
);

INVx2_ASAP7_75t_L g7898 ( 
.A(n_7163),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_7448),
.Y(n_7899)
);

HB1xp67_ASAP7_75t_L g7900 ( 
.A(n_7451),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7449),
.Y(n_7901)
);

INVxp67_ASAP7_75t_L g7902 ( 
.A(n_7583),
.Y(n_7902)
);

NAND2xp5_ASAP7_75t_L g7903 ( 
.A(n_7362),
.B(n_6041),
.Y(n_7903)
);

BUFx8_ASAP7_75t_L g7904 ( 
.A(n_7576),
.Y(n_7904)
);

AND2x2_ASAP7_75t_L g7905 ( 
.A(n_7231),
.B(n_5531),
.Y(n_7905)
);

INVx2_ASAP7_75t_SL g7906 ( 
.A(n_7098),
.Y(n_7906)
);

CKINVDCx5p33_ASAP7_75t_R g7907 ( 
.A(n_7166),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7165),
.Y(n_7908)
);

INVx4_ASAP7_75t_L g7909 ( 
.A(n_7172),
.Y(n_7909)
);

INVx2_ASAP7_75t_L g7910 ( 
.A(n_7169),
.Y(n_7910)
);

INVx3_ASAP7_75t_L g7911 ( 
.A(n_7170),
.Y(n_7911)
);

AOI22xp5_ASAP7_75t_L g7912 ( 
.A1(n_7558),
.A2(n_5670),
.B1(n_5680),
.B2(n_5640),
.Y(n_7912)
);

CKINVDCx16_ASAP7_75t_R g7913 ( 
.A(n_7116),
.Y(n_7913)
);

BUFx3_ASAP7_75t_L g7914 ( 
.A(n_7380),
.Y(n_7914)
);

BUFx6f_ASAP7_75t_L g7915 ( 
.A(n_7173),
.Y(n_7915)
);

NOR2xp33_ASAP7_75t_L g7916 ( 
.A(n_7559),
.B(n_6049),
.Y(n_7916)
);

BUFx2_ASAP7_75t_L g7917 ( 
.A(n_7473),
.Y(n_7917)
);

AND2x4_ASAP7_75t_L g7918 ( 
.A(n_7562),
.B(n_6170),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7174),
.Y(n_7919)
);

CKINVDCx5p33_ASAP7_75t_R g7920 ( 
.A(n_7188),
.Y(n_7920)
);

INVx1_ASAP7_75t_L g7921 ( 
.A(n_7175),
.Y(n_7921)
);

OAI22x1_ASAP7_75t_SL g7922 ( 
.A1(n_7168),
.A2(n_5653),
.B1(n_5659),
.B2(n_5650),
.Y(n_7922)
);

NAND2xp5_ASAP7_75t_L g7923 ( 
.A(n_7376),
.B(n_6217),
.Y(n_7923)
);

AOI22x1_ASAP7_75t_SL g7924 ( 
.A1(n_7124),
.A2(n_5665),
.B1(n_5692),
.B2(n_5663),
.Y(n_7924)
);

BUFx6f_ASAP7_75t_L g7925 ( 
.A(n_7176),
.Y(n_7925)
);

OAI21x1_ASAP7_75t_L g7926 ( 
.A1(n_7569),
.A2(n_5409),
.B(n_5402),
.Y(n_7926)
);

BUFx6f_ASAP7_75t_L g7927 ( 
.A(n_7177),
.Y(n_7927)
);

INVx2_ASAP7_75t_L g7928 ( 
.A(n_7179),
.Y(n_7928)
);

BUFx8_ASAP7_75t_L g7929 ( 
.A(n_7577),
.Y(n_7929)
);

HB1xp67_ASAP7_75t_L g7930 ( 
.A(n_7454),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7180),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7181),
.Y(n_7932)
);

NAND2xp5_ASAP7_75t_L g7933 ( 
.A(n_7413),
.B(n_6325),
.Y(n_7933)
);

AOI22xp5_ASAP7_75t_L g7934 ( 
.A1(n_7563),
.A2(n_5828),
.B1(n_5855),
.B2(n_5714),
.Y(n_7934)
);

OAI22x1_ASAP7_75t_L g7935 ( 
.A1(n_7578),
.A2(n_5894),
.B1(n_5898),
.B2(n_5889),
.Y(n_7935)
);

OA21x2_ASAP7_75t_L g7936 ( 
.A1(n_7570),
.A2(n_5224),
.B(n_5223),
.Y(n_7936)
);

INVx2_ASAP7_75t_L g7937 ( 
.A(n_7183),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7184),
.Y(n_7938)
);

BUFx6f_ASAP7_75t_L g7939 ( 
.A(n_7185),
.Y(n_7939)
);

INVx1_ASAP7_75t_L g7940 ( 
.A(n_7186),
.Y(n_7940)
);

INVx2_ASAP7_75t_L g7941 ( 
.A(n_7189),
.Y(n_7941)
);

BUFx6f_ASAP7_75t_L g7942 ( 
.A(n_7196),
.Y(n_7942)
);

INVx5_ASAP7_75t_L g7943 ( 
.A(n_7128),
.Y(n_7943)
);

INVx2_ASAP7_75t_L g7944 ( 
.A(n_7197),
.Y(n_7944)
);

AND2x2_ASAP7_75t_L g7945 ( 
.A(n_7236),
.B(n_5531),
.Y(n_7945)
);

CKINVDCx5p33_ASAP7_75t_R g7946 ( 
.A(n_7190),
.Y(n_7946)
);

INVx5_ASAP7_75t_L g7947 ( 
.A(n_7568),
.Y(n_7947)
);

INVx3_ASAP7_75t_L g7948 ( 
.A(n_7199),
.Y(n_7948)
);

INVx2_ASAP7_75t_L g7949 ( 
.A(n_7201),
.Y(n_7949)
);

INVx2_ASAP7_75t_L g7950 ( 
.A(n_7202),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7204),
.Y(n_7951)
);

BUFx6f_ASAP7_75t_L g7952 ( 
.A(n_7206),
.Y(n_7952)
);

OA21x2_ASAP7_75t_L g7953 ( 
.A1(n_7426),
.A2(n_5242),
.B(n_5239),
.Y(n_7953)
);

AND2x4_ASAP7_75t_L g7954 ( 
.A(n_7564),
.B(n_6373),
.Y(n_7954)
);

HB1xp67_ASAP7_75t_L g7955 ( 
.A(n_7269),
.Y(n_7955)
);

OAI22xp5_ASAP7_75t_L g7956 ( 
.A1(n_7565),
.A2(n_5360),
.B1(n_5361),
.B2(n_5359),
.Y(n_7956)
);

CKINVDCx6p67_ASAP7_75t_R g7957 ( 
.A(n_7125),
.Y(n_7957)
);

INVx2_ASAP7_75t_L g7958 ( 
.A(n_7209),
.Y(n_7958)
);

INVxp67_ASAP7_75t_L g7959 ( 
.A(n_7579),
.Y(n_7959)
);

INVx2_ASAP7_75t_L g7960 ( 
.A(n_7210),
.Y(n_7960)
);

CKINVDCx16_ASAP7_75t_R g7961 ( 
.A(n_7129),
.Y(n_7961)
);

INVx3_ASAP7_75t_L g7962 ( 
.A(n_7211),
.Y(n_7962)
);

BUFx2_ASAP7_75t_L g7963 ( 
.A(n_7477),
.Y(n_7963)
);

INVx2_ASAP7_75t_L g7964 ( 
.A(n_7212),
.Y(n_7964)
);

BUFx6f_ASAP7_75t_L g7965 ( 
.A(n_7217),
.Y(n_7965)
);

BUFx3_ASAP7_75t_L g7966 ( 
.A(n_7384),
.Y(n_7966)
);

INVx1_ASAP7_75t_L g7967 ( 
.A(n_7218),
.Y(n_7967)
);

NAND2xp5_ASAP7_75t_L g7968 ( 
.A(n_7442),
.B(n_6536),
.Y(n_7968)
);

BUFx6f_ASAP7_75t_L g7969 ( 
.A(n_7219),
.Y(n_7969)
);

INVx3_ASAP7_75t_L g7970 ( 
.A(n_7220),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_7223),
.Y(n_7971)
);

AND2x2_ASAP7_75t_SL g7972 ( 
.A(n_7415),
.B(n_5410),
.Y(n_7972)
);

INVx3_ASAP7_75t_L g7973 ( 
.A(n_7224),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_7226),
.Y(n_7974)
);

BUFx6f_ASAP7_75t_L g7975 ( 
.A(n_7230),
.Y(n_7975)
);

INVx2_ASAP7_75t_L g7976 ( 
.A(n_7232),
.Y(n_7976)
);

INVx2_ASAP7_75t_L g7977 ( 
.A(n_7234),
.Y(n_7977)
);

OA21x2_ASAP7_75t_L g7978 ( 
.A1(n_7235),
.A2(n_5245),
.B(n_5243),
.Y(n_7978)
);

INVx6_ASAP7_75t_L g7979 ( 
.A(n_7590),
.Y(n_7979)
);

INVx3_ASAP7_75t_L g7980 ( 
.A(n_7237),
.Y(n_7980)
);

INVx6_ASAP7_75t_L g7981 ( 
.A(n_7596),
.Y(n_7981)
);

INVx5_ASAP7_75t_L g7982 ( 
.A(n_7482),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_7238),
.Y(n_7983)
);

AND2x4_ASAP7_75t_L g7984 ( 
.A(n_7412),
.B(n_5249),
.Y(n_7984)
);

AND2x4_ASAP7_75t_L g7985 ( 
.A(n_7424),
.B(n_5263),
.Y(n_7985)
);

AND2x4_ASAP7_75t_L g7986 ( 
.A(n_7445),
.B(n_7490),
.Y(n_7986)
);

BUFx12f_ASAP7_75t_L g7987 ( 
.A(n_7466),
.Y(n_7987)
);

BUFx6f_ASAP7_75t_L g7988 ( 
.A(n_7240),
.Y(n_7988)
);

INVx4_ASAP7_75t_L g7989 ( 
.A(n_7192),
.Y(n_7989)
);

INVx2_ASAP7_75t_SL g7990 ( 
.A(n_7132),
.Y(n_7990)
);

AND2x4_ASAP7_75t_L g7991 ( 
.A(n_7506),
.B(n_5270),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7241),
.Y(n_7992)
);

INVx2_ASAP7_75t_L g7993 ( 
.A(n_7242),
.Y(n_7993)
);

INVx2_ASAP7_75t_L g7994 ( 
.A(n_7245),
.Y(n_7994)
);

CKINVDCx6p67_ASAP7_75t_R g7995 ( 
.A(n_7478),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_7247),
.Y(n_7996)
);

BUFx8_ASAP7_75t_L g7997 ( 
.A(n_7289),
.Y(n_7997)
);

INVx2_ASAP7_75t_L g7998 ( 
.A(n_7248),
.Y(n_7998)
);

OAI22xp5_ASAP7_75t_SL g7999 ( 
.A1(n_7479),
.A2(n_5709),
.B1(n_5769),
.B2(n_5705),
.Y(n_7999)
);

INVx2_ASAP7_75t_L g8000 ( 
.A(n_7251),
.Y(n_8000)
);

BUFx12f_ASAP7_75t_L g8001 ( 
.A(n_7470),
.Y(n_8001)
);

AOI22xp5_ASAP7_75t_L g8002 ( 
.A1(n_7195),
.A2(n_6026),
.B1(n_6100),
.B2(n_5932),
.Y(n_8002)
);

INVx2_ASAP7_75t_L g8003 ( 
.A(n_7252),
.Y(n_8003)
);

AND2x4_ASAP7_75t_L g8004 ( 
.A(n_7543),
.B(n_5271),
.Y(n_8004)
);

HB1xp67_ASAP7_75t_L g8005 ( 
.A(n_7152),
.Y(n_8005)
);

AND2x4_ASAP7_75t_L g8006 ( 
.A(n_7253),
.B(n_5274),
.Y(n_8006)
);

INVx3_ASAP7_75t_L g8007 ( 
.A(n_7254),
.Y(n_8007)
);

AND2x4_ASAP7_75t_L g8008 ( 
.A(n_7259),
.B(n_5276),
.Y(n_8008)
);

BUFx6f_ASAP7_75t_L g8009 ( 
.A(n_7261),
.Y(n_8009)
);

INVx5_ASAP7_75t_L g8010 ( 
.A(n_7265),
.Y(n_8010)
);

AOI22xp5_ASAP7_75t_L g8011 ( 
.A1(n_7200),
.A2(n_6168),
.B1(n_6192),
.B2(n_6122),
.Y(n_8011)
);

INVx1_ASAP7_75t_L g8012 ( 
.A(n_7262),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_7263),
.Y(n_8013)
);

INVx3_ASAP7_75t_L g8014 ( 
.A(n_7266),
.Y(n_8014)
);

INVx1_ASAP7_75t_L g8015 ( 
.A(n_7267),
.Y(n_8015)
);

INVx2_ASAP7_75t_L g8016 ( 
.A(n_7268),
.Y(n_8016)
);

BUFx6f_ASAP7_75t_L g8017 ( 
.A(n_7086),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7088),
.Y(n_8018)
);

NAND2xp5_ASAP7_75t_L g8019 ( 
.A(n_7089),
.B(n_5413),
.Y(n_8019)
);

AND2x4_ASAP7_75t_L g8020 ( 
.A(n_7208),
.B(n_5278),
.Y(n_8020)
);

INVx2_ASAP7_75t_L g8021 ( 
.A(n_7090),
.Y(n_8021)
);

NOR2xp33_ASAP7_75t_L g8022 ( 
.A(n_7203),
.B(n_7215),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7091),
.B(n_5431),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_7092),
.Y(n_8024)
);

BUFx6f_ASAP7_75t_L g8025 ( 
.A(n_7094),
.Y(n_8025)
);

BUFx6f_ASAP7_75t_L g8026 ( 
.A(n_7096),
.Y(n_8026)
);

BUFx6f_ASAP7_75t_L g8027 ( 
.A(n_7100),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_7101),
.Y(n_8028)
);

INVx1_ASAP7_75t_L g8029 ( 
.A(n_7102),
.Y(n_8029)
);

CKINVDCx16_ASAP7_75t_R g8030 ( 
.A(n_7207),
.Y(n_8030)
);

INVx2_ASAP7_75t_L g8031 ( 
.A(n_7103),
.Y(n_8031)
);

INVx2_ASAP7_75t_L g8032 ( 
.A(n_7586),
.Y(n_8032)
);

INVx2_ASAP7_75t_L g8033 ( 
.A(n_7588),
.Y(n_8033)
);

INVx4_ASAP7_75t_L g8034 ( 
.A(n_7228),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_7589),
.Y(n_8035)
);

BUFx6f_ASAP7_75t_L g8036 ( 
.A(n_7592),
.Y(n_8036)
);

INVx4_ASAP7_75t_L g8037 ( 
.A(n_7249),
.Y(n_8037)
);

INVx2_ASAP7_75t_L g8038 ( 
.A(n_7595),
.Y(n_8038)
);

AOI22xp5_ASAP7_75t_L g8039 ( 
.A1(n_7250),
.A2(n_7255),
.B1(n_7272),
.B2(n_7257),
.Y(n_8039)
);

INVx3_ASAP7_75t_L g8040 ( 
.A(n_7597),
.Y(n_8040)
);

BUFx3_ASAP7_75t_L g8041 ( 
.A(n_7389),
.Y(n_8041)
);

CKINVDCx5p33_ASAP7_75t_R g8042 ( 
.A(n_7273),
.Y(n_8042)
);

BUFx6f_ASAP7_75t_L g8043 ( 
.A(n_7598),
.Y(n_8043)
);

INVx2_ASAP7_75t_L g8044 ( 
.A(n_7603),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_7606),
.Y(n_8045)
);

INVx3_ASAP7_75t_L g8046 ( 
.A(n_7609),
.Y(n_8046)
);

INVx2_ASAP7_75t_L g8047 ( 
.A(n_7610),
.Y(n_8047)
);

INVx6_ASAP7_75t_L g8048 ( 
.A(n_7225),
.Y(n_8048)
);

CKINVDCx20_ASAP7_75t_R g8049 ( 
.A(n_7113),
.Y(n_8049)
);

INVx1_ASAP7_75t_L g8050 ( 
.A(n_7246),
.Y(n_8050)
);

AND2x6_ASAP7_75t_L g8051 ( 
.A(n_7311),
.B(n_6195),
.Y(n_8051)
);

NAND2xp5_ASAP7_75t_L g8052 ( 
.A(n_7274),
.B(n_5452),
.Y(n_8052)
);

AOI22x1_ASAP7_75t_SL g8053 ( 
.A1(n_7591),
.A2(n_5813),
.B1(n_5851),
.B2(n_5790),
.Y(n_8053)
);

OAI21x1_ASAP7_75t_L g8054 ( 
.A1(n_7292),
.A2(n_5543),
.B(n_5515),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_7346),
.Y(n_8055)
);

INVx6_ASAP7_75t_L g8056 ( 
.A(n_7229),
.Y(n_8056)
);

AND2x2_ASAP7_75t_L g8057 ( 
.A(n_7363),
.B(n_5645),
.Y(n_8057)
);

INVx2_ASAP7_75t_SL g8058 ( 
.A(n_7604),
.Y(n_8058)
);

INVx5_ASAP7_75t_L g8059 ( 
.A(n_7312),
.Y(n_8059)
);

AND2x4_ASAP7_75t_L g8060 ( 
.A(n_7278),
.B(n_5280),
.Y(n_8060)
);

OA21x2_ASAP7_75t_L g8061 ( 
.A1(n_7284),
.A2(n_5282),
.B(n_5281),
.Y(n_8061)
);

BUFx2_ASAP7_75t_L g8062 ( 
.A(n_7485),
.Y(n_8062)
);

BUFx6f_ASAP7_75t_L g8063 ( 
.A(n_7474),
.Y(n_8063)
);

NAND2xp5_ASAP7_75t_L g8064 ( 
.A(n_7290),
.B(n_5559),
.Y(n_8064)
);

NOR2xp33_ASAP7_75t_SL g8065 ( 
.A(n_7484),
.B(n_5867),
.Y(n_8065)
);

INVx2_ASAP7_75t_SL g8066 ( 
.A(n_7500),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7301),
.Y(n_8067)
);

BUFx6f_ASAP7_75t_L g8068 ( 
.A(n_7501),
.Y(n_8068)
);

OA21x2_ASAP7_75t_L g8069 ( 
.A1(n_7302),
.A2(n_5286),
.B(n_5283),
.Y(n_8069)
);

INVx1_ASAP7_75t_L g8070 ( 
.A(n_7305),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7306),
.Y(n_8071)
);

HB1xp67_ASAP7_75t_L g8072 ( 
.A(n_7505),
.Y(n_8072)
);

INVx4_ASAP7_75t_L g8073 ( 
.A(n_7308),
.Y(n_8073)
);

NAND2xp5_ASAP7_75t_L g8074 ( 
.A(n_7309),
.B(n_5581),
.Y(n_8074)
);

AND2x6_ASAP7_75t_L g8075 ( 
.A(n_7422),
.B(n_6224),
.Y(n_8075)
);

BUFx3_ASAP7_75t_L g8076 ( 
.A(n_7390),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7321),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7325),
.Y(n_8078)
);

AND2x2_ASAP7_75t_L g8079 ( 
.A(n_7510),
.B(n_5645),
.Y(n_8079)
);

INVx3_ASAP7_75t_L g8080 ( 
.A(n_7514),
.Y(n_8080)
);

AND2x2_ASAP7_75t_L g8081 ( 
.A(n_7517),
.B(n_5707),
.Y(n_8081)
);

BUFx6f_ASAP7_75t_L g8082 ( 
.A(n_7518),
.Y(n_8082)
);

NAND2xp5_ASAP7_75t_L g8083 ( 
.A(n_7326),
.B(n_7330),
.Y(n_8083)
);

BUFx6f_ASAP7_75t_L g8084 ( 
.A(n_7532),
.Y(n_8084)
);

AND2x2_ASAP7_75t_L g8085 ( 
.A(n_7535),
.B(n_5707),
.Y(n_8085)
);

OA21x2_ASAP7_75t_L g8086 ( 
.A1(n_7335),
.A2(n_5293),
.B(n_5290),
.Y(n_8086)
);

INVx3_ASAP7_75t_L g8087 ( 
.A(n_7540),
.Y(n_8087)
);

AND2x4_ASAP7_75t_L g8088 ( 
.A(n_7340),
.B(n_5296),
.Y(n_8088)
);

BUFx3_ASAP7_75t_L g8089 ( 
.A(n_7409),
.Y(n_8089)
);

INVx2_ASAP7_75t_L g8090 ( 
.A(n_7348),
.Y(n_8090)
);

NAND2xp5_ASAP7_75t_L g8091 ( 
.A(n_7350),
.B(n_5616),
.Y(n_8091)
);

NAND2xp5_ASAP7_75t_L g8092 ( 
.A(n_7354),
.B(n_5646),
.Y(n_8092)
);

INVx2_ASAP7_75t_SL g8093 ( 
.A(n_7541),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_7360),
.Y(n_8094)
);

INVx1_ASAP7_75t_L g8095 ( 
.A(n_7364),
.Y(n_8095)
);

BUFx6f_ASAP7_75t_L g8096 ( 
.A(n_7545),
.Y(n_8096)
);

INVx2_ASAP7_75t_L g8097 ( 
.A(n_7365),
.Y(n_8097)
);

BUFx6f_ASAP7_75t_L g8098 ( 
.A(n_7547),
.Y(n_8098)
);

NAND2xp5_ASAP7_75t_L g8099 ( 
.A(n_7366),
.B(n_5685),
.Y(n_8099)
);

INVx2_ASAP7_75t_SL g8100 ( 
.A(n_7548),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7379),
.Y(n_8101)
);

AND2x2_ASAP7_75t_L g8102 ( 
.A(n_7549),
.B(n_7556),
.Y(n_8102)
);

INVx3_ASAP7_75t_L g8103 ( 
.A(n_7557),
.Y(n_8103)
);

BUFx2_ASAP7_75t_L g8104 ( 
.A(n_7493),
.Y(n_8104)
);

AND2x2_ASAP7_75t_L g8105 ( 
.A(n_7382),
.B(n_5751),
.Y(n_8105)
);

INVx2_ASAP7_75t_L g8106 ( 
.A(n_7385),
.Y(n_8106)
);

BUFx2_ASAP7_75t_L g8107 ( 
.A(n_7525),
.Y(n_8107)
);

AND2x4_ASAP7_75t_L g8108 ( 
.A(n_7387),
.B(n_5298),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7393),
.Y(n_8109)
);

AND2x6_ASAP7_75t_L g8110 ( 
.A(n_7436),
.B(n_6287),
.Y(n_8110)
);

AOI22x1_ASAP7_75t_SL g8111 ( 
.A1(n_7593),
.A2(n_5920),
.B1(n_5970),
.B2(n_5879),
.Y(n_8111)
);

BUFx6f_ASAP7_75t_L g8112 ( 
.A(n_7395),
.Y(n_8112)
);

BUFx6f_ASAP7_75t_L g8113 ( 
.A(n_7416),
.Y(n_8113)
);

INVx2_ASAP7_75t_L g8114 ( 
.A(n_7585),
.Y(n_8114)
);

AND2x2_ASAP7_75t_L g8115 ( 
.A(n_7594),
.B(n_7599),
.Y(n_8115)
);

NOR2x1_ASAP7_75t_L g8116 ( 
.A(n_7530),
.B(n_5862),
.Y(n_8116)
);

INVx2_ASAP7_75t_L g8117 ( 
.A(n_7600),
.Y(n_8117)
);

INVx2_ASAP7_75t_L g8118 ( 
.A(n_7602),
.Y(n_8118)
);

AND2x2_ASAP7_75t_SL g8119 ( 
.A(n_7567),
.B(n_5690),
.Y(n_8119)
);

NAND2xp5_ASAP7_75t_L g8120 ( 
.A(n_7607),
.B(n_5693),
.Y(n_8120)
);

OAI22xp5_ASAP7_75t_L g8121 ( 
.A1(n_7611),
.A2(n_5364),
.B1(n_5366),
.B2(n_5363),
.Y(n_8121)
);

AND2x2_ASAP7_75t_L g8122 ( 
.A(n_7571),
.B(n_7580),
.Y(n_8122)
);

AND2x2_ASAP7_75t_L g8123 ( 
.A(n_7582),
.B(n_5751),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_7443),
.Y(n_8124)
);

INVxp67_ASAP7_75t_L g8125 ( 
.A(n_7233),
.Y(n_8125)
);

HB1xp67_ASAP7_75t_L g8126 ( 
.A(n_7244),
.Y(n_8126)
);

INVx1_ASAP7_75t_L g8127 ( 
.A(n_7605),
.Y(n_8127)
);

NAND2xp5_ASAP7_75t_L g8128 ( 
.A(n_7608),
.B(n_5716),
.Y(n_8128)
);

OAI22x1_ASAP7_75t_SL g8129 ( 
.A1(n_7258),
.A2(n_5997),
.B1(n_5998),
.B2(n_5985),
.Y(n_8129)
);

NAND2xp5_ASAP7_75t_L g8130 ( 
.A(n_7320),
.B(n_5767),
.Y(n_8130)
);

INVx2_ASAP7_75t_L g8131 ( 
.A(n_7121),
.Y(n_8131)
);

NOR2xp33_ASAP7_75t_L g8132 ( 
.A(n_7285),
.B(n_5372),
.Y(n_8132)
);

AOI22xp5_ASAP7_75t_L g8133 ( 
.A1(n_7187),
.A2(n_6462),
.B1(n_6467),
.B2(n_6345),
.Y(n_8133)
);

OR2x2_ASAP7_75t_L g8134 ( 
.A(n_7285),
.B(n_6489),
.Y(n_8134)
);

INVx2_ASAP7_75t_SL g8135 ( 
.A(n_7573),
.Y(n_8135)
);

INVx2_ASAP7_75t_L g8136 ( 
.A(n_7121),
.Y(n_8136)
);

INVx1_ASAP7_75t_L g8137 ( 
.A(n_7313),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7121),
.Y(n_8138)
);

INVx2_ASAP7_75t_L g8139 ( 
.A(n_7121),
.Y(n_8139)
);

OA21x2_ASAP7_75t_L g8140 ( 
.A1(n_7483),
.A2(n_5302),
.B(n_5301),
.Y(n_8140)
);

BUFx6f_ASAP7_75t_L g8141 ( 
.A(n_7194),
.Y(n_8141)
);

AND2x2_ASAP7_75t_L g8142 ( 
.A(n_7572),
.B(n_5786),
.Y(n_8142)
);

AND2x4_ASAP7_75t_L g8143 ( 
.A(n_7198),
.B(n_5305),
.Y(n_8143)
);

OA21x2_ASAP7_75t_L g8144 ( 
.A1(n_7483),
.A2(n_5311),
.B(n_5309),
.Y(n_8144)
);

AND2x4_ASAP7_75t_L g8145 ( 
.A(n_7198),
.B(n_5312),
.Y(n_8145)
);

INVx1_ASAP7_75t_L g8146 ( 
.A(n_7313),
.Y(n_8146)
);

AND2x4_ASAP7_75t_L g8147 ( 
.A(n_7198),
.B(n_5314),
.Y(n_8147)
);

BUFx3_ASAP7_75t_L g8148 ( 
.A(n_7198),
.Y(n_8148)
);

INVx2_ASAP7_75t_L g8149 ( 
.A(n_7121),
.Y(n_8149)
);

OAI21x1_ASAP7_75t_L g8150 ( 
.A1(n_7483),
.A2(n_5801),
.B(n_5792),
.Y(n_8150)
);

AND2x2_ASAP7_75t_L g8151 ( 
.A(n_7572),
.B(n_5786),
.Y(n_8151)
);

BUFx6f_ASAP7_75t_L g8152 ( 
.A(n_7194),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7121),
.Y(n_8153)
);

OA21x2_ASAP7_75t_L g8154 ( 
.A1(n_7483),
.A2(n_5320),
.B(n_5316),
.Y(n_8154)
);

AND2x2_ASAP7_75t_L g8155 ( 
.A(n_7572),
.B(n_5934),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7313),
.Y(n_8156)
);

AND2x6_ASAP7_75t_L g8157 ( 
.A(n_7538),
.B(n_6497),
.Y(n_8157)
);

INVx2_ASAP7_75t_L g8158 ( 
.A(n_7121),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_7313),
.Y(n_8159)
);

INVx3_ASAP7_75t_L g8160 ( 
.A(n_7194),
.Y(n_8160)
);

INVx2_ASAP7_75t_L g8161 ( 
.A(n_7121),
.Y(n_8161)
);

AOI22x1_ASAP7_75t_SL g8162 ( 
.A1(n_7264),
.A2(n_6004),
.B1(n_6005),
.B2(n_6000),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_7121),
.Y(n_8163)
);

BUFx2_ASAP7_75t_L g8164 ( 
.A(n_7464),
.Y(n_8164)
);

OA21x2_ASAP7_75t_L g8165 ( 
.A1(n_7483),
.A2(n_5327),
.B(n_5325),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7320),
.B(n_5808),
.Y(n_8166)
);

CKINVDCx8_ASAP7_75t_R g8167 ( 
.A(n_7464),
.Y(n_8167)
);

BUFx6f_ASAP7_75t_L g8168 ( 
.A(n_7194),
.Y(n_8168)
);

INVx2_ASAP7_75t_SL g8169 ( 
.A(n_7573),
.Y(n_8169)
);

BUFx6f_ASAP7_75t_L g8170 ( 
.A(n_7194),
.Y(n_8170)
);

INVx2_ASAP7_75t_L g8171 ( 
.A(n_7121),
.Y(n_8171)
);

BUFx3_ASAP7_75t_L g8172 ( 
.A(n_7198),
.Y(n_8172)
);

CKINVDCx11_ASAP7_75t_R g8173 ( 
.A(n_7264),
.Y(n_8173)
);

INVx2_ASAP7_75t_L g8174 ( 
.A(n_7121),
.Y(n_8174)
);

BUFx12f_ASAP7_75t_L g8175 ( 
.A(n_7417),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_7313),
.Y(n_8176)
);

INVx2_ASAP7_75t_L g8177 ( 
.A(n_7121),
.Y(n_8177)
);

BUFx12f_ASAP7_75t_L g8178 ( 
.A(n_7417),
.Y(n_8178)
);

OAI22xp5_ASAP7_75t_SL g8179 ( 
.A1(n_7584),
.A2(n_6042),
.B1(n_6053),
.B2(n_6039),
.Y(n_8179)
);

BUFx2_ASAP7_75t_L g8180 ( 
.A(n_7464),
.Y(n_8180)
);

BUFx6f_ASAP7_75t_L g8181 ( 
.A(n_7194),
.Y(n_8181)
);

INVx2_ASAP7_75t_L g8182 ( 
.A(n_7121),
.Y(n_8182)
);

AOI22xp5_ASAP7_75t_L g8183 ( 
.A1(n_7187),
.A2(n_6529),
.B1(n_6537),
.B2(n_6513),
.Y(n_8183)
);

BUFx8_ASAP7_75t_L g8184 ( 
.A(n_7120),
.Y(n_8184)
);

AND2x2_ASAP7_75t_L g8185 ( 
.A(n_7572),
.B(n_5934),
.Y(n_8185)
);

OAI21x1_ASAP7_75t_L g8186 ( 
.A1(n_7483),
.A2(n_5913),
.B(n_5886),
.Y(n_8186)
);

OAI21x1_ASAP7_75t_L g8187 ( 
.A1(n_7483),
.A2(n_5978),
.B(n_5937),
.Y(n_8187)
);

HB1xp67_ASAP7_75t_L g8188 ( 
.A(n_7584),
.Y(n_8188)
);

OAI22x1_ASAP7_75t_SL g8189 ( 
.A1(n_7433),
.A2(n_6066),
.B1(n_6067),
.B2(n_6056),
.Y(n_8189)
);

AND2x2_ASAP7_75t_L g8190 ( 
.A(n_7572),
.B(n_5963),
.Y(n_8190)
);

INVx2_ASAP7_75t_SL g8191 ( 
.A(n_7573),
.Y(n_8191)
);

INVx5_ASAP7_75t_L g8192 ( 
.A(n_7143),
.Y(n_8192)
);

BUFx6f_ASAP7_75t_L g8193 ( 
.A(n_7194),
.Y(n_8193)
);

INVx2_ASAP7_75t_L g8194 ( 
.A(n_7121),
.Y(n_8194)
);

INVx3_ASAP7_75t_L g8195 ( 
.A(n_7635),
.Y(n_8195)
);

CKINVDCx20_ASAP7_75t_R g8196 ( 
.A(n_7878),
.Y(n_8196)
);

INVxp33_ASAP7_75t_L g8197 ( 
.A(n_8188),
.Y(n_8197)
);

HB1xp67_ASAP7_75t_L g8198 ( 
.A(n_7666),
.Y(n_8198)
);

AND2x4_ASAP7_75t_L g8199 ( 
.A(n_8148),
.B(n_5330),
.Y(n_8199)
);

INVx1_ASAP7_75t_L g8200 ( 
.A(n_7865),
.Y(n_8200)
);

CKINVDCx5p33_ASAP7_75t_R g8201 ( 
.A(n_7620),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7867),
.Y(n_8202)
);

NAND2xp5_ASAP7_75t_SL g8203 ( 
.A(n_7623),
.B(n_5375),
.Y(n_8203)
);

BUFx3_ASAP7_75t_L g8204 ( 
.A(n_8172),
.Y(n_8204)
);

INVx2_ASAP7_75t_L g8205 ( 
.A(n_7721),
.Y(n_8205)
);

AND2x2_ASAP7_75t_L g8206 ( 
.A(n_7691),
.B(n_5963),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7726),
.Y(n_8207)
);

CKINVDCx20_ASAP7_75t_R g8208 ( 
.A(n_7690),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_7880),
.Y(n_8209)
);

CKINVDCx5p33_ASAP7_75t_R g8210 ( 
.A(n_7742),
.Y(n_8210)
);

CKINVDCx5p33_ASAP7_75t_R g8211 ( 
.A(n_7787),
.Y(n_8211)
);

INVxp67_ASAP7_75t_L g8212 ( 
.A(n_8134),
.Y(n_8212)
);

CKINVDCx5p33_ASAP7_75t_R g8213 ( 
.A(n_7842),
.Y(n_8213)
);

CKINVDCx5p33_ASAP7_75t_R g8214 ( 
.A(n_7847),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_7886),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7889),
.Y(n_8216)
);

CKINVDCx5p33_ASAP7_75t_R g8217 ( 
.A(n_7851),
.Y(n_8217)
);

INVx1_ASAP7_75t_L g8218 ( 
.A(n_7890),
.Y(n_8218)
);

CKINVDCx20_ASAP7_75t_R g8219 ( 
.A(n_7761),
.Y(n_8219)
);

INVx1_ASAP7_75t_L g8220 ( 
.A(n_7899),
.Y(n_8220)
);

HB1xp67_ASAP7_75t_L g8221 ( 
.A(n_7631),
.Y(n_8221)
);

INVx1_ASAP7_75t_L g8222 ( 
.A(n_7901),
.Y(n_8222)
);

INVx1_ASAP7_75t_L g8223 ( 
.A(n_7908),
.Y(n_8223)
);

INVx2_ASAP7_75t_L g8224 ( 
.A(n_7738),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7921),
.Y(n_8225)
);

BUFx6f_ASAP7_75t_L g8226 ( 
.A(n_7630),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7931),
.Y(n_8227)
);

CKINVDCx5p33_ASAP7_75t_R g8228 ( 
.A(n_7907),
.Y(n_8228)
);

NAND2xp5_ASAP7_75t_SL g8229 ( 
.A(n_7657),
.B(n_5379),
.Y(n_8229)
);

BUFx2_ASAP7_75t_L g8230 ( 
.A(n_7654),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_7632),
.B(n_5384),
.Y(n_8231)
);

CKINVDCx5p33_ASAP7_75t_R g8232 ( 
.A(n_7920),
.Y(n_8232)
);

BUFx6f_ASAP7_75t_L g8233 ( 
.A(n_7636),
.Y(n_8233)
);

INVx3_ASAP7_75t_L g8234 ( 
.A(n_7659),
.Y(n_8234)
);

INVx2_ASAP7_75t_L g8235 ( 
.A(n_7743),
.Y(n_8235)
);

NAND2xp5_ASAP7_75t_L g8236 ( 
.A(n_7621),
.B(n_5385),
.Y(n_8236)
);

CKINVDCx5p33_ASAP7_75t_R g8237 ( 
.A(n_7946),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7932),
.Y(n_8238)
);

INVx3_ASAP7_75t_L g8239 ( 
.A(n_7671),
.Y(n_8239)
);

NOR2xp33_ASAP7_75t_L g8240 ( 
.A(n_7700),
.B(n_6553),
.Y(n_8240)
);

NAND2xp5_ASAP7_75t_L g8241 ( 
.A(n_7625),
.B(n_5386),
.Y(n_8241)
);

INVx2_ASAP7_75t_L g8242 ( 
.A(n_7702),
.Y(n_8242)
);

CKINVDCx5p33_ASAP7_75t_R g8243 ( 
.A(n_8042),
.Y(n_8243)
);

INVx2_ASAP7_75t_L g8244 ( 
.A(n_7780),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_7938),
.Y(n_8245)
);

INVx1_ASAP7_75t_L g8246 ( 
.A(n_7940),
.Y(n_8246)
);

OA21x2_ASAP7_75t_L g8247 ( 
.A1(n_7642),
.A2(n_5347),
.B(n_5346),
.Y(n_8247)
);

AND2x6_ASAP7_75t_L g8248 ( 
.A(n_7701),
.B(n_5356),
.Y(n_8248)
);

CKINVDCx20_ASAP7_75t_R g8249 ( 
.A(n_7775),
.Y(n_8249)
);

CKINVDCx5p33_ASAP7_75t_R g8250 ( 
.A(n_7669),
.Y(n_8250)
);

INVx1_ASAP7_75t_L g8251 ( 
.A(n_7951),
.Y(n_8251)
);

INVx2_ASAP7_75t_L g8252 ( 
.A(n_7693),
.Y(n_8252)
);

CKINVDCx5p33_ASAP7_75t_R g8253 ( 
.A(n_8173),
.Y(n_8253)
);

INVx2_ASAP7_75t_L g8254 ( 
.A(n_7706),
.Y(n_8254)
);

NAND2xp33_ASAP7_75t_R g8255 ( 
.A(n_7683),
.B(n_7703),
.Y(n_8255)
);

INVx2_ASAP7_75t_L g8256 ( 
.A(n_7718),
.Y(n_8256)
);

CKINVDCx5p33_ASAP7_75t_R g8257 ( 
.A(n_7643),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7967),
.Y(n_8258)
);

CKINVDCx20_ASAP7_75t_R g8259 ( 
.A(n_7845),
.Y(n_8259)
);

CKINVDCx20_ASAP7_75t_R g8260 ( 
.A(n_8049),
.Y(n_8260)
);

BUFx6f_ASAP7_75t_L g8261 ( 
.A(n_7641),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_7971),
.Y(n_8262)
);

CKINVDCx5p33_ASAP7_75t_R g8263 ( 
.A(n_7648),
.Y(n_8263)
);

CKINVDCx5p33_ASAP7_75t_R g8264 ( 
.A(n_7692),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_7974),
.Y(n_8265)
);

CKINVDCx20_ASAP7_75t_R g8266 ( 
.A(n_8030),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_7992),
.Y(n_8267)
);

CKINVDCx20_ASAP7_75t_R g8268 ( 
.A(n_7913),
.Y(n_8268)
);

INVx1_ASAP7_75t_L g8269 ( 
.A(n_7996),
.Y(n_8269)
);

BUFx6f_ASAP7_75t_L g8270 ( 
.A(n_7616),
.Y(n_8270)
);

INVx2_ASAP7_75t_L g8271 ( 
.A(n_8021),
.Y(n_8271)
);

INVx2_ASAP7_75t_L g8272 ( 
.A(n_8031),
.Y(n_8272)
);

CKINVDCx5p33_ASAP7_75t_R g8273 ( 
.A(n_7723),
.Y(n_8273)
);

NOR2xp33_ASAP7_75t_L g8274 ( 
.A(n_8132),
.B(n_5387),
.Y(n_8274)
);

INVx2_ASAP7_75t_L g8275 ( 
.A(n_8032),
.Y(n_8275)
);

CKINVDCx5p33_ASAP7_75t_R g8276 ( 
.A(n_7741),
.Y(n_8276)
);

NAND2xp5_ASAP7_75t_L g8277 ( 
.A(n_7629),
.B(n_5390),
.Y(n_8277)
);

CKINVDCx20_ASAP7_75t_R g8278 ( 
.A(n_7961),
.Y(n_8278)
);

INVx3_ASAP7_75t_L g8279 ( 
.A(n_7685),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_8012),
.Y(n_8280)
);

INVx1_ASAP7_75t_L g8281 ( 
.A(n_8013),
.Y(n_8281)
);

NAND2xp5_ASAP7_75t_L g8282 ( 
.A(n_7633),
.B(n_5391),
.Y(n_8282)
);

NOR2xp33_ASAP7_75t_SL g8283 ( 
.A(n_7759),
.B(n_6112),
.Y(n_8283)
);

CKINVDCx5p33_ASAP7_75t_R g8284 ( 
.A(n_7795),
.Y(n_8284)
);

CKINVDCx20_ASAP7_75t_R g8285 ( 
.A(n_7995),
.Y(n_8285)
);

CKINVDCx5p33_ASAP7_75t_R g8286 ( 
.A(n_7829),
.Y(n_8286)
);

INVx2_ASAP7_75t_L g8287 ( 
.A(n_8033),
.Y(n_8287)
);

INVx1_ASAP7_75t_L g8288 ( 
.A(n_8015),
.Y(n_8288)
);

INVx3_ASAP7_75t_L g8289 ( 
.A(n_7663),
.Y(n_8289)
);

INVx1_ASAP7_75t_L g8290 ( 
.A(n_7841),
.Y(n_8290)
);

INVx2_ASAP7_75t_L g8291 ( 
.A(n_8038),
.Y(n_8291)
);

CKINVDCx5p33_ASAP7_75t_R g8292 ( 
.A(n_7893),
.Y(n_8292)
);

AND2x4_ASAP7_75t_L g8293 ( 
.A(n_7650),
.B(n_5362),
.Y(n_8293)
);

CKINVDCx20_ASAP7_75t_R g8294 ( 
.A(n_7957),
.Y(n_8294)
);

CKINVDCx5p33_ASAP7_75t_R g8295 ( 
.A(n_7987),
.Y(n_8295)
);

CKINVDCx5p33_ASAP7_75t_R g8296 ( 
.A(n_8001),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7844),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_7853),
.Y(n_8298)
);

BUFx10_ASAP7_75t_L g8299 ( 
.A(n_8022),
.Y(n_8299)
);

INVx2_ASAP7_75t_L g8300 ( 
.A(n_8044),
.Y(n_8300)
);

INVx2_ASAP7_75t_L g8301 ( 
.A(n_8047),
.Y(n_8301)
);

CKINVDCx5p33_ASAP7_75t_R g8302 ( 
.A(n_8175),
.Y(n_8302)
);

BUFx6f_ASAP7_75t_L g8303 ( 
.A(n_7619),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_7855),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_7861),
.Y(n_8305)
);

CKINVDCx5p33_ASAP7_75t_R g8306 ( 
.A(n_8178),
.Y(n_8306)
);

CKINVDCx20_ASAP7_75t_R g8307 ( 
.A(n_8167),
.Y(n_8307)
);

NAND2xp5_ASAP7_75t_L g8308 ( 
.A(n_7638),
.B(n_5396),
.Y(n_8308)
);

BUFx3_ASAP7_75t_L g8309 ( 
.A(n_8048),
.Y(n_8309)
);

CKINVDCx5p33_ASAP7_75t_R g8310 ( 
.A(n_8063),
.Y(n_8310)
);

CKINVDCx5p33_ASAP7_75t_R g8311 ( 
.A(n_8068),
.Y(n_8311)
);

CKINVDCx5p33_ASAP7_75t_R g8312 ( 
.A(n_8082),
.Y(n_8312)
);

AND2x4_ASAP7_75t_L g8313 ( 
.A(n_8143),
.B(n_5377),
.Y(n_8313)
);

INVx2_ASAP7_75t_L g8314 ( 
.A(n_7781),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_7646),
.Y(n_8315)
);

CKINVDCx5p33_ASAP7_75t_R g8316 ( 
.A(n_8084),
.Y(n_8316)
);

INVx2_ASAP7_75t_L g8317 ( 
.A(n_7799),
.Y(n_8317)
);

CKINVDCx5p33_ASAP7_75t_R g8318 ( 
.A(n_8096),
.Y(n_8318)
);

INVx1_ASAP7_75t_L g8319 ( 
.A(n_7652),
.Y(n_8319)
);

INVx2_ASAP7_75t_L g8320 ( 
.A(n_7803),
.Y(n_8320)
);

INVx2_ASAP7_75t_L g8321 ( 
.A(n_7811),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7656),
.Y(n_8322)
);

BUFx2_ASAP7_75t_L g8323 ( 
.A(n_8164),
.Y(n_8323)
);

CKINVDCx5p33_ASAP7_75t_R g8324 ( 
.A(n_8098),
.Y(n_8324)
);

INVx2_ASAP7_75t_L g8325 ( 
.A(n_7812),
.Y(n_8325)
);

NAND2xp5_ASAP7_75t_L g8326 ( 
.A(n_7660),
.B(n_5399),
.Y(n_8326)
);

INVx3_ASAP7_75t_L g8327 ( 
.A(n_8017),
.Y(n_8327)
);

HB1xp67_ASAP7_75t_L g8328 ( 
.A(n_8180),
.Y(n_8328)
);

NOR2xp33_ASAP7_75t_R g8329 ( 
.A(n_8080),
.B(n_6127),
.Y(n_8329)
);

CKINVDCx5p33_ASAP7_75t_R g8330 ( 
.A(n_8112),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_7673),
.Y(n_8331)
);

CKINVDCx5p33_ASAP7_75t_R g8332 ( 
.A(n_8113),
.Y(n_8332)
);

NAND2xp33_ASAP7_75t_L g8333 ( 
.A(n_7758),
.B(n_5400),
.Y(n_8333)
);

AND2x4_ASAP7_75t_L g8334 ( 
.A(n_8145),
.B(n_5380),
.Y(n_8334)
);

NAND2xp5_ASAP7_75t_L g8335 ( 
.A(n_7676),
.B(n_5401),
.Y(n_8335)
);

AND2x2_ASAP7_75t_L g8336 ( 
.A(n_8142),
.B(n_5981),
.Y(n_8336)
);

INVx1_ASAP7_75t_L g8337 ( 
.A(n_7684),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_7696),
.Y(n_8338)
);

NOR2xp33_ASAP7_75t_L g8339 ( 
.A(n_8052),
.B(n_5407),
.Y(n_8339)
);

AND2x2_ASAP7_75t_L g8340 ( 
.A(n_8151),
.B(n_5981),
.Y(n_8340)
);

CKINVDCx20_ASAP7_75t_R g8341 ( 
.A(n_7734),
.Y(n_8341)
);

CKINVDCx5p33_ASAP7_75t_R g8342 ( 
.A(n_8056),
.Y(n_8342)
);

INVx2_ASAP7_75t_L g8343 ( 
.A(n_7815),
.Y(n_8343)
);

CKINVDCx16_ASAP7_75t_R g8344 ( 
.A(n_8065),
.Y(n_8344)
);

CKINVDCx5p33_ASAP7_75t_R g8345 ( 
.A(n_7695),
.Y(n_8345)
);

INVx2_ASAP7_75t_L g8346 ( 
.A(n_7816),
.Y(n_8346)
);

BUFx6f_ASAP7_75t_L g8347 ( 
.A(n_8141),
.Y(n_8347)
);

INVx3_ASAP7_75t_L g8348 ( 
.A(n_8025),
.Y(n_8348)
);

CKINVDCx20_ASAP7_75t_R g8349 ( 
.A(n_7707),
.Y(n_8349)
);

NOR2xp33_ASAP7_75t_L g8350 ( 
.A(n_8064),
.B(n_5408),
.Y(n_8350)
);

CKINVDCx5p33_ASAP7_75t_R g8351 ( 
.A(n_7735),
.Y(n_8351)
);

BUFx2_ASAP7_75t_L g8352 ( 
.A(n_7751),
.Y(n_8352)
);

BUFx6f_ASAP7_75t_L g8353 ( 
.A(n_8152),
.Y(n_8353)
);

CKINVDCx5p33_ASAP7_75t_R g8354 ( 
.A(n_7739),
.Y(n_8354)
);

INVx1_ASAP7_75t_L g8355 ( 
.A(n_7699),
.Y(n_8355)
);

CKINVDCx5p33_ASAP7_75t_R g8356 ( 
.A(n_7755),
.Y(n_8356)
);

AND2x2_ASAP7_75t_L g8357 ( 
.A(n_8155),
.B(n_6017),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_7818),
.Y(n_8358)
);

BUFx10_ASAP7_75t_L g8359 ( 
.A(n_7789),
.Y(n_8359)
);

HB1xp67_ASAP7_75t_L g8360 ( 
.A(n_7622),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_7705),
.Y(n_8361)
);

INVx2_ASAP7_75t_SL g8362 ( 
.A(n_7637),
.Y(n_8362)
);

OR2x2_ASAP7_75t_L g8363 ( 
.A(n_8128),
.B(n_6095),
.Y(n_8363)
);

AND2x2_ASAP7_75t_L g8364 ( 
.A(n_8185),
.B(n_6017),
.Y(n_8364)
);

INVx1_ASAP7_75t_L g8365 ( 
.A(n_7708),
.Y(n_8365)
);

INVx2_ASAP7_75t_L g8366 ( 
.A(n_7831),
.Y(n_8366)
);

NOR2xp33_ASAP7_75t_R g8367 ( 
.A(n_8087),
.B(n_6147),
.Y(n_8367)
);

INVx1_ASAP7_75t_L g8368 ( 
.A(n_7711),
.Y(n_8368)
);

CKINVDCx5p33_ASAP7_75t_R g8369 ( 
.A(n_7772),
.Y(n_8369)
);

CKINVDCx5p33_ASAP7_75t_R g8370 ( 
.A(n_7857),
.Y(n_8370)
);

BUFx6f_ASAP7_75t_L g8371 ( 
.A(n_8168),
.Y(n_8371)
);

INVx2_ASAP7_75t_L g8372 ( 
.A(n_7834),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7712),
.Y(n_8373)
);

CKINVDCx5p33_ASAP7_75t_R g8374 ( 
.A(n_7881),
.Y(n_8374)
);

INVx3_ASAP7_75t_L g8375 ( 
.A(n_8026),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7715),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_7720),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_7722),
.Y(n_8378)
);

CKINVDCx20_ASAP7_75t_R g8379 ( 
.A(n_7914),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7724),
.Y(n_8380)
);

NAND2xp5_ASAP7_75t_L g8381 ( 
.A(n_7725),
.B(n_5415),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_7728),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_7732),
.Y(n_8383)
);

CKINVDCx20_ASAP7_75t_R g8384 ( 
.A(n_7966),
.Y(n_8384)
);

INVx2_ASAP7_75t_L g8385 ( 
.A(n_7836),
.Y(n_8385)
);

INVx3_ASAP7_75t_L g8386 ( 
.A(n_8027),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7748),
.Y(n_8387)
);

NOR2xp33_ASAP7_75t_L g8388 ( 
.A(n_8074),
.B(n_5416),
.Y(n_8388)
);

BUFx2_ASAP7_75t_L g8389 ( 
.A(n_7762),
.Y(n_8389)
);

CKINVDCx20_ASAP7_75t_R g8390 ( 
.A(n_8041),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_7749),
.Y(n_8391)
);

NOR2xp33_ASAP7_75t_R g8392 ( 
.A(n_8103),
.B(n_6154),
.Y(n_8392)
);

INVx3_ASAP7_75t_L g8393 ( 
.A(n_8036),
.Y(n_8393)
);

INVxp67_ASAP7_75t_L g8394 ( 
.A(n_7698),
.Y(n_8394)
);

CKINVDCx5p33_ASAP7_75t_R g8395 ( 
.A(n_8076),
.Y(n_8395)
);

NAND2xp5_ASAP7_75t_SL g8396 ( 
.A(n_7627),
.B(n_5417),
.Y(n_8396)
);

OR2x6_ASAP7_75t_L g8397 ( 
.A(n_7820),
.B(n_5383),
.Y(n_8397)
);

CKINVDCx5p33_ASAP7_75t_R g8398 ( 
.A(n_8089),
.Y(n_8398)
);

BUFx6f_ASAP7_75t_L g8399 ( 
.A(n_8170),
.Y(n_8399)
);

CKINVDCx5p33_ASAP7_75t_R g8400 ( 
.A(n_8039),
.Y(n_8400)
);

NAND2xp5_ASAP7_75t_L g8401 ( 
.A(n_7752),
.B(n_5418),
.Y(n_8401)
);

CKINVDCx5p33_ASAP7_75t_R g8402 ( 
.A(n_7817),
.Y(n_8402)
);

CKINVDCx5p33_ASAP7_75t_R g8403 ( 
.A(n_7837),
.Y(n_8403)
);

INVx2_ASAP7_75t_L g8404 ( 
.A(n_7839),
.Y(n_8404)
);

CKINVDCx5p33_ASAP7_75t_R g8405 ( 
.A(n_7885),
.Y(n_8405)
);

INVx1_ASAP7_75t_L g8406 ( 
.A(n_7757),
.Y(n_8406)
);

INVx3_ASAP7_75t_L g8407 ( 
.A(n_8043),
.Y(n_8407)
);

HB1xp67_ASAP7_75t_L g8408 ( 
.A(n_7821),
.Y(n_8408)
);

CKINVDCx5p33_ASAP7_75t_R g8409 ( 
.A(n_7909),
.Y(n_8409)
);

AND2x2_ASAP7_75t_L g8410 ( 
.A(n_8190),
.B(n_6038),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_7763),
.Y(n_8411)
);

AOI22xp5_ASAP7_75t_L g8412 ( 
.A1(n_7758),
.A2(n_6190),
.B1(n_6218),
.B2(n_6175),
.Y(n_8412)
);

CKINVDCx20_ASAP7_75t_R g8413 ( 
.A(n_7773),
.Y(n_8413)
);

CKINVDCx20_ASAP7_75t_R g8414 ( 
.A(n_7868),
.Y(n_8414)
);

BUFx6f_ASAP7_75t_L g8415 ( 
.A(n_8181),
.Y(n_8415)
);

INVx2_ASAP7_75t_L g8416 ( 
.A(n_7848),
.Y(n_8416)
);

INVxp67_ASAP7_75t_L g8417 ( 
.A(n_7710),
.Y(n_8417)
);

INVx3_ASAP7_75t_L g8418 ( 
.A(n_8193),
.Y(n_8418)
);

CKINVDCx5p33_ASAP7_75t_R g8419 ( 
.A(n_7989),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_7764),
.Y(n_8420)
);

CKINVDCx5p33_ASAP7_75t_R g8421 ( 
.A(n_8034),
.Y(n_8421)
);

INVx2_ASAP7_75t_L g8422 ( 
.A(n_7850),
.Y(n_8422)
);

INVx3_ASAP7_75t_L g8423 ( 
.A(n_7791),
.Y(n_8423)
);

HB1xp67_ASAP7_75t_L g8424 ( 
.A(n_7828),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_7778),
.B(n_5421),
.Y(n_8425)
);

INVx1_ASAP7_75t_L g8426 ( 
.A(n_7779),
.Y(n_8426)
);

CKINVDCx5p33_ASAP7_75t_R g8427 ( 
.A(n_8037),
.Y(n_8427)
);

INVx1_ASAP7_75t_L g8428 ( 
.A(n_7788),
.Y(n_8428)
);

HB1xp67_ASAP7_75t_L g8429 ( 
.A(n_7840),
.Y(n_8429)
);

INVx4_ASAP7_75t_L g8430 ( 
.A(n_7982),
.Y(n_8430)
);

NOR2xp33_ASAP7_75t_R g8431 ( 
.A(n_7618),
.B(n_6285),
.Y(n_8431)
);

INVx1_ASAP7_75t_L g8432 ( 
.A(n_7792),
.Y(n_8432)
);

AND2x2_ASAP7_75t_SL g8433 ( 
.A(n_8119),
.B(n_6007),
.Y(n_8433)
);

INVx1_ASAP7_75t_L g8434 ( 
.A(n_7793),
.Y(n_8434)
);

CKINVDCx20_ASAP7_75t_R g8435 ( 
.A(n_7917),
.Y(n_8435)
);

AND2x2_ASAP7_75t_SL g8436 ( 
.A(n_7753),
.B(n_6031),
.Y(n_8436)
);

INVx2_ASAP7_75t_SL g8437 ( 
.A(n_7651),
.Y(n_8437)
);

CKINVDCx5p33_ASAP7_75t_R g8438 ( 
.A(n_8073),
.Y(n_8438)
);

OAI21x1_ASAP7_75t_L g8439 ( 
.A1(n_7806),
.A2(n_6128),
.B(n_6091),
.Y(n_8439)
);

CKINVDCx5p33_ASAP7_75t_R g8440 ( 
.A(n_7997),
.Y(n_8440)
);

OR2x2_ASAP7_75t_L g8441 ( 
.A(n_8135),
.B(n_5423),
.Y(n_8441)
);

INVx2_ASAP7_75t_L g8442 ( 
.A(n_7856),
.Y(n_8442)
);

INVx3_ASAP7_75t_L g8443 ( 
.A(n_7822),
.Y(n_8443)
);

INVx2_ASAP7_75t_L g8444 ( 
.A(n_7860),
.Y(n_8444)
);

INVx2_ASAP7_75t_L g8445 ( 
.A(n_7863),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_7798),
.Y(n_8446)
);

NOR2x1_ASAP7_75t_L g8447 ( 
.A(n_8083),
.B(n_6286),
.Y(n_8447)
);

AND2x2_ASAP7_75t_L g8448 ( 
.A(n_7801),
.B(n_6038),
.Y(n_8448)
);

BUFx6f_ASAP7_75t_L g8449 ( 
.A(n_7870),
.Y(n_8449)
);

NAND2xp5_ASAP7_75t_L g8450 ( 
.A(n_7800),
.B(n_5428),
.Y(n_8450)
);

CKINVDCx5p33_ASAP7_75t_R g8451 ( 
.A(n_7963),
.Y(n_8451)
);

CKINVDCx20_ASAP7_75t_R g8452 ( 
.A(n_8062),
.Y(n_8452)
);

AND2x2_ASAP7_75t_L g8453 ( 
.A(n_8169),
.B(n_6109),
.Y(n_8453)
);

INVx2_ASAP7_75t_L g8454 ( 
.A(n_7873),
.Y(n_8454)
);

INVx3_ASAP7_75t_L g8455 ( 
.A(n_7823),
.Y(n_8455)
);

CKINVDCx20_ASAP7_75t_R g8456 ( 
.A(n_8104),
.Y(n_8456)
);

NAND2xp5_ASAP7_75t_SL g8457 ( 
.A(n_8191),
.B(n_5433),
.Y(n_8457)
);

BUFx2_ASAP7_75t_L g8458 ( 
.A(n_8157),
.Y(n_8458)
);

CKINVDCx16_ASAP7_75t_R g8459 ( 
.A(n_7854),
.Y(n_8459)
);

INVxp67_ASAP7_75t_L g8460 ( 
.A(n_7713),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_7804),
.Y(n_8461)
);

NAND2xp5_ASAP7_75t_L g8462 ( 
.A(n_7813),
.B(n_5439),
.Y(n_8462)
);

BUFx6f_ASAP7_75t_L g8463 ( 
.A(n_7877),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_7824),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7830),
.Y(n_8465)
);

INVxp67_ASAP7_75t_L g8466 ( 
.A(n_7827),
.Y(n_8466)
);

HB1xp67_ASAP7_75t_L g8467 ( 
.A(n_7879),
.Y(n_8467)
);

CKINVDCx20_ASAP7_75t_R g8468 ( 
.A(n_8107),
.Y(n_8468)
);

AND2x2_ASAP7_75t_L g8469 ( 
.A(n_7677),
.B(n_6109),
.Y(n_8469)
);

CKINVDCx5p33_ASAP7_75t_R g8470 ( 
.A(n_8102),
.Y(n_8470)
);

AND2x2_ASAP7_75t_L g8471 ( 
.A(n_7765),
.B(n_6142),
.Y(n_8471)
);

AND2x2_ASAP7_75t_L g8472 ( 
.A(n_7717),
.B(n_6142),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_8137),
.B(n_5440),
.Y(n_8473)
);

BUFx10_ASAP7_75t_L g8474 ( 
.A(n_7874),
.Y(n_8474)
);

INVx2_ASAP7_75t_L g8475 ( 
.A(n_7884),
.Y(n_8475)
);

INVx1_ASAP7_75t_L g8476 ( 
.A(n_8146),
.Y(n_8476)
);

CKINVDCx5p33_ASAP7_75t_R g8477 ( 
.A(n_8115),
.Y(n_8477)
);

INVx2_ASAP7_75t_L g8478 ( 
.A(n_7898),
.Y(n_8478)
);

INVx1_ASAP7_75t_L g8479 ( 
.A(n_8156),
.Y(n_8479)
);

OAI21x1_ASAP7_75t_L g8480 ( 
.A1(n_7807),
.A2(n_6160),
.B(n_6136),
.Y(n_8480)
);

INVx3_ASAP7_75t_L g8481 ( 
.A(n_7832),
.Y(n_8481)
);

CKINVDCx5p33_ASAP7_75t_R g8482 ( 
.A(n_8072),
.Y(n_8482)
);

CKINVDCx5p33_ASAP7_75t_R g8483 ( 
.A(n_7979),
.Y(n_8483)
);

CKINVDCx5p33_ASAP7_75t_R g8484 ( 
.A(n_7981),
.Y(n_8484)
);

OAI22xp5_ASAP7_75t_SL g8485 ( 
.A1(n_7999),
.A2(n_6380),
.B1(n_6382),
.B2(n_6365),
.Y(n_8485)
);

CKINVDCx5p33_ASAP7_75t_R g8486 ( 
.A(n_8010),
.Y(n_8486)
);

AND2x4_ASAP7_75t_L g8487 ( 
.A(n_8147),
.B(n_5388),
.Y(n_8487)
);

BUFx6f_ASAP7_75t_L g8488 ( 
.A(n_8006),
.Y(n_8488)
);

INVx1_ASAP7_75t_L g8489 ( 
.A(n_8159),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_8176),
.Y(n_8490)
);

CKINVDCx5p33_ASAP7_75t_R g8491 ( 
.A(n_8059),
.Y(n_8491)
);

BUFx2_ASAP7_75t_L g8492 ( 
.A(n_8157),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_8018),
.Y(n_8493)
);

INVx1_ASAP7_75t_L g8494 ( 
.A(n_8024),
.Y(n_8494)
);

CKINVDCx20_ASAP7_75t_R g8495 ( 
.A(n_7678),
.Y(n_8495)
);

CKINVDCx20_ASAP7_75t_R g8496 ( 
.A(n_8184),
.Y(n_8496)
);

CKINVDCx5p33_ASAP7_75t_R g8497 ( 
.A(n_7649),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_8028),
.Y(n_8498)
);

INVx1_ASAP7_75t_L g8499 ( 
.A(n_8029),
.Y(n_8499)
);

INVx2_ASAP7_75t_L g8500 ( 
.A(n_7910),
.Y(n_8500)
);

NAND2xp5_ASAP7_75t_L g8501 ( 
.A(n_8130),
.B(n_5441),
.Y(n_8501)
);

BUFx10_ASAP7_75t_L g8502 ( 
.A(n_8051),
.Y(n_8502)
);

INVx1_ASAP7_75t_L g8503 ( 
.A(n_8035),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_8045),
.Y(n_8504)
);

AND2x2_ASAP7_75t_L g8505 ( 
.A(n_7770),
.B(n_6277),
.Y(n_8505)
);

BUFx6f_ASAP7_75t_L g8506 ( 
.A(n_8008),
.Y(n_8506)
);

AND2x2_ASAP7_75t_L g8507 ( 
.A(n_7662),
.B(n_6277),
.Y(n_8507)
);

OAI22xp5_ASAP7_75t_SL g8508 ( 
.A1(n_8179),
.A2(n_6431),
.B1(n_6434),
.B2(n_6410),
.Y(n_8508)
);

AND2x2_ASAP7_75t_L g8509 ( 
.A(n_7838),
.B(n_6293),
.Y(n_8509)
);

CKINVDCx5p33_ASAP7_75t_R g8510 ( 
.A(n_7687),
.Y(n_8510)
);

AND2x2_ASAP7_75t_L g8511 ( 
.A(n_7887),
.B(n_6293),
.Y(n_8511)
);

INVx2_ASAP7_75t_L g8512 ( 
.A(n_7919),
.Y(n_8512)
);

NAND2xp33_ASAP7_75t_SL g8513 ( 
.A(n_8079),
.B(n_6469),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_7928),
.Y(n_8514)
);

INVx2_ASAP7_75t_L g8515 ( 
.A(n_7937),
.Y(n_8515)
);

AND2x4_ASAP7_75t_L g8516 ( 
.A(n_7681),
.B(n_7686),
.Y(n_8516)
);

BUFx6f_ASAP7_75t_L g8517 ( 
.A(n_7833),
.Y(n_8517)
);

BUFx8_ASAP7_75t_L g8518 ( 
.A(n_8051),
.Y(n_8518)
);

CKINVDCx5p33_ASAP7_75t_R g8519 ( 
.A(n_7746),
.Y(n_8519)
);

INVx2_ASAP7_75t_L g8520 ( 
.A(n_7941),
.Y(n_8520)
);

NAND2xp5_ASAP7_75t_L g8521 ( 
.A(n_8166),
.B(n_5445),
.Y(n_8521)
);

BUFx6f_ASAP7_75t_L g8522 ( 
.A(n_7843),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_7944),
.Y(n_8523)
);

CKINVDCx20_ASAP7_75t_R g8524 ( 
.A(n_8192),
.Y(n_8524)
);

INVx2_ASAP7_75t_L g8525 ( 
.A(n_7949),
.Y(n_8525)
);

NAND2xp5_ASAP7_75t_L g8526 ( 
.A(n_7859),
.B(n_7670),
.Y(n_8526)
);

NOR2xp33_ASAP7_75t_SL g8527 ( 
.A(n_7808),
.B(n_6483),
.Y(n_8527)
);

INVx1_ASAP7_75t_L g8528 ( 
.A(n_7950),
.Y(n_8528)
);

INVx2_ASAP7_75t_L g8529 ( 
.A(n_7958),
.Y(n_8529)
);

OA21x2_ASAP7_75t_L g8530 ( 
.A1(n_8150),
.A2(n_8187),
.B(n_8186),
.Y(n_8530)
);

INVx1_ASAP7_75t_L g8531 ( 
.A(n_7960),
.Y(n_8531)
);

NAND2xp5_ASAP7_75t_L g8532 ( 
.A(n_7754),
.B(n_5448),
.Y(n_8532)
);

AND2x2_ASAP7_75t_L g8533 ( 
.A(n_7905),
.B(n_6359),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_SL g8534 ( 
.A(n_8091),
.B(n_8092),
.Y(n_8534)
);

BUFx2_ASAP7_75t_L g8535 ( 
.A(n_7875),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_7964),
.Y(n_8536)
);

AND2x2_ASAP7_75t_L g8537 ( 
.A(n_7945),
.B(n_6359),
.Y(n_8537)
);

CKINVDCx5p33_ASAP7_75t_R g8538 ( 
.A(n_8066),
.Y(n_8538)
);

NAND2xp5_ASAP7_75t_L g8539 ( 
.A(n_7784),
.B(n_5449),
.Y(n_8539)
);

INVx1_ASAP7_75t_L g8540 ( 
.A(n_7976),
.Y(n_8540)
);

INVx1_ASAP7_75t_SL g8541 ( 
.A(n_7900),
.Y(n_8541)
);

CKINVDCx5p33_ASAP7_75t_R g8542 ( 
.A(n_8093),
.Y(n_8542)
);

NAND2xp5_ASAP7_75t_SL g8543 ( 
.A(n_8099),
.B(n_5451),
.Y(n_8543)
);

CKINVDCx20_ASAP7_75t_R g8544 ( 
.A(n_7776),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_7977),
.Y(n_8545)
);

INVx3_ASAP7_75t_L g8546 ( 
.A(n_7760),
.Y(n_8546)
);

CKINVDCx20_ASAP7_75t_R g8547 ( 
.A(n_8126),
.Y(n_8547)
);

AND2x2_ASAP7_75t_L g8548 ( 
.A(n_7972),
.B(n_6394),
.Y(n_8548)
);

NAND2xp5_ASAP7_75t_L g8549 ( 
.A(n_7894),
.B(n_5453),
.Y(n_8549)
);

INVxp67_ASAP7_75t_L g8550 ( 
.A(n_7930),
.Y(n_8550)
);

INVx1_ASAP7_75t_L g8551 ( 
.A(n_7983),
.Y(n_8551)
);

INVx2_ASAP7_75t_L g8552 ( 
.A(n_7993),
.Y(n_8552)
);

INVx2_ASAP7_75t_L g8553 ( 
.A(n_7994),
.Y(n_8553)
);

NOR2xp33_ASAP7_75t_R g8554 ( 
.A(n_8124),
.B(n_6496),
.Y(n_8554)
);

CKINVDCx20_ASAP7_75t_R g8555 ( 
.A(n_7729),
.Y(n_8555)
);

CKINVDCx5p33_ASAP7_75t_R g8556 ( 
.A(n_8100),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_7998),
.Y(n_8557)
);

INVx2_ASAP7_75t_L g8558 ( 
.A(n_8000),
.Y(n_8558)
);

CKINVDCx5p33_ASAP7_75t_R g8559 ( 
.A(n_8122),
.Y(n_8559)
);

INVx1_ASAP7_75t_L g8560 ( 
.A(n_8003),
.Y(n_8560)
);

BUFx6f_ASAP7_75t_L g8561 ( 
.A(n_7689),
.Y(n_8561)
);

INVx1_ASAP7_75t_L g8562 ( 
.A(n_8016),
.Y(n_8562)
);

NAND2xp5_ASAP7_75t_L g8563 ( 
.A(n_7896),
.B(n_7916),
.Y(n_8563)
);

CKINVDCx5p33_ASAP7_75t_R g8564 ( 
.A(n_8090),
.Y(n_8564)
);

NOR2xp33_ASAP7_75t_L g8565 ( 
.A(n_8120),
.B(n_5458),
.Y(n_8565)
);

NAND2xp5_ASAP7_75t_L g8566 ( 
.A(n_7953),
.B(n_7876),
.Y(n_8566)
);

BUFx6f_ASAP7_75t_L g8567 ( 
.A(n_7694),
.Y(n_8567)
);

INVx2_ASAP7_75t_L g8568 ( 
.A(n_7634),
.Y(n_8568)
);

NOR2xp33_ASAP7_75t_L g8569 ( 
.A(n_7615),
.B(n_5459),
.Y(n_8569)
);

NAND2xp5_ASAP7_75t_L g8570 ( 
.A(n_7730),
.B(n_7733),
.Y(n_8570)
);

INVx2_ASAP7_75t_L g8571 ( 
.A(n_7644),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_8040),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_8046),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_7645),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_7658),
.Y(n_8575)
);

CKINVDCx5p33_ASAP7_75t_R g8576 ( 
.A(n_8097),
.Y(n_8576)
);

CKINVDCx5p33_ASAP7_75t_R g8577 ( 
.A(n_8106),
.Y(n_8577)
);

CKINVDCx5p33_ASAP7_75t_R g8578 ( 
.A(n_8109),
.Y(n_8578)
);

HB1xp67_ASAP7_75t_L g8579 ( 
.A(n_8061),
.Y(n_8579)
);

CKINVDCx5p33_ASAP7_75t_R g8580 ( 
.A(n_8114),
.Y(n_8580)
);

INVx2_ASAP7_75t_L g8581 ( 
.A(n_7672),
.Y(n_8581)
);

INVx1_ASAP7_75t_L g8582 ( 
.A(n_7675),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_7680),
.Y(n_8583)
);

INVx2_ASAP7_75t_L g8584 ( 
.A(n_8131),
.Y(n_8584)
);

OAI22xp5_ASAP7_75t_SL g8585 ( 
.A1(n_7943),
.A2(n_6566),
.B1(n_6577),
.B2(n_6560),
.Y(n_8585)
);

AND2x4_ASAP7_75t_L g8586 ( 
.A(n_7688),
.B(n_5389),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_8136),
.Y(n_8587)
);

INVx1_ASAP7_75t_L g8588 ( 
.A(n_8138),
.Y(n_8588)
);

INVx1_ASAP7_75t_L g8589 ( 
.A(n_8139),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_8149),
.Y(n_8590)
);

CKINVDCx5p33_ASAP7_75t_R g8591 ( 
.A(n_8117),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_8153),
.Y(n_8592)
);

INVx1_ASAP7_75t_L g8593 ( 
.A(n_8158),
.Y(n_8593)
);

CKINVDCx5p33_ASAP7_75t_R g8594 ( 
.A(n_8118),
.Y(n_8594)
);

CKINVDCx20_ASAP7_75t_R g8595 ( 
.A(n_8125),
.Y(n_8595)
);

AND2x6_ASAP7_75t_L g8596 ( 
.A(n_8067),
.B(n_5393),
.Y(n_8596)
);

CKINVDCx20_ASAP7_75t_R g8597 ( 
.A(n_7947),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_8161),
.Y(n_8598)
);

NAND2xp5_ASAP7_75t_L g8599 ( 
.A(n_7737),
.B(n_5465),
.Y(n_8599)
);

INVx2_ASAP7_75t_L g8600 ( 
.A(n_8163),
.Y(n_8600)
);

NOR2xp33_ASAP7_75t_L g8601 ( 
.A(n_7794),
.B(n_5466),
.Y(n_8601)
);

CKINVDCx20_ASAP7_75t_R g8602 ( 
.A(n_8005),
.Y(n_8602)
);

NAND2xp5_ASAP7_75t_L g8603 ( 
.A(n_7767),
.B(n_5472),
.Y(n_8603)
);

AND2x4_ASAP7_75t_L g8604 ( 
.A(n_7709),
.B(n_7714),
.Y(n_8604)
);

INVx1_ASAP7_75t_L g8605 ( 
.A(n_8171),
.Y(n_8605)
);

NAND2xp33_ASAP7_75t_R g8606 ( 
.A(n_8069),
.B(n_5474),
.Y(n_8606)
);

NAND2xp5_ASAP7_75t_L g8607 ( 
.A(n_7785),
.B(n_5475),
.Y(n_8607)
);

INVx2_ASAP7_75t_L g8608 ( 
.A(n_8174),
.Y(n_8608)
);

INVx3_ASAP7_75t_L g8609 ( 
.A(n_7777),
.Y(n_8609)
);

INVx1_ASAP7_75t_L g8610 ( 
.A(n_8177),
.Y(n_8610)
);

CKINVDCx20_ASAP7_75t_R g8611 ( 
.A(n_8127),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_8182),
.Y(n_8612)
);

INVx1_ASAP7_75t_L g8613 ( 
.A(n_8194),
.Y(n_8613)
);

BUFx6f_ASAP7_75t_L g8614 ( 
.A(n_7697),
.Y(n_8614)
);

INVx2_ASAP7_75t_L g8615 ( 
.A(n_7745),
.Y(n_8615)
);

INVx1_ASAP7_75t_L g8616 ( 
.A(n_7750),
.Y(n_8616)
);

INVx2_ASAP7_75t_L g8617 ( 
.A(n_7911),
.Y(n_8617)
);

INVx2_ASAP7_75t_L g8618 ( 
.A(n_7948),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_7962),
.Y(n_8619)
);

CKINVDCx5p33_ASAP7_75t_R g8620 ( 
.A(n_8070),
.Y(n_8620)
);

CKINVDCx20_ASAP7_75t_R g8621 ( 
.A(n_7906),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_7970),
.Y(n_8622)
);

INVx1_ASAP7_75t_L g8623 ( 
.A(n_7973),
.Y(n_8623)
);

AND2x2_ASAP7_75t_L g8624 ( 
.A(n_8081),
.B(n_6394),
.Y(n_8624)
);

INVx2_ASAP7_75t_L g8625 ( 
.A(n_7980),
.Y(n_8625)
);

INVx2_ASAP7_75t_L g8626 ( 
.A(n_8007),
.Y(n_8626)
);

INVx2_ASAP7_75t_L g8627 ( 
.A(n_8014),
.Y(n_8627)
);

INVx1_ASAP7_75t_L g8628 ( 
.A(n_7978),
.Y(n_8628)
);

CKINVDCx20_ASAP7_75t_R g8629 ( 
.A(n_7990),
.Y(n_8629)
);

CKINVDCx5p33_ASAP7_75t_R g8630 ( 
.A(n_8071),
.Y(n_8630)
);

INVx1_ASAP7_75t_L g8631 ( 
.A(n_8019),
.Y(n_8631)
);

HB1xp67_ASAP7_75t_L g8632 ( 
.A(n_8086),
.Y(n_8632)
);

AND2x4_ASAP7_75t_L g8633 ( 
.A(n_7653),
.B(n_7769),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_8023),
.Y(n_8634)
);

AND2x4_ASAP7_75t_L g8635 ( 
.A(n_7786),
.B(n_5395),
.Y(n_8635)
);

INVx1_ASAP7_75t_L g8636 ( 
.A(n_7802),
.Y(n_8636)
);

CKINVDCx5p33_ASAP7_75t_R g8637 ( 
.A(n_8077),
.Y(n_8637)
);

CKINVDCx5p33_ASAP7_75t_R g8638 ( 
.A(n_8078),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_8140),
.Y(n_8639)
);

INVx2_ASAP7_75t_L g8640 ( 
.A(n_7612),
.Y(n_8640)
);

INVx1_ASAP7_75t_L g8641 ( 
.A(n_8144),
.Y(n_8641)
);

INVx2_ASAP7_75t_L g8642 ( 
.A(n_8160),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_8154),
.Y(n_8643)
);

INVx3_ASAP7_75t_L g8644 ( 
.A(n_7719),
.Y(n_8644)
);

INVx2_ASAP7_75t_L g8645 ( 
.A(n_7849),
.Y(n_8645)
);

CKINVDCx5p33_ASAP7_75t_R g8646 ( 
.A(n_8094),
.Y(n_8646)
);

CKINVDCx5p33_ASAP7_75t_R g8647 ( 
.A(n_8095),
.Y(n_8647)
);

NAND2xp5_ASAP7_75t_L g8648 ( 
.A(n_7888),
.B(n_5477),
.Y(n_8648)
);

CKINVDCx20_ASAP7_75t_R g8649 ( 
.A(n_8058),
.Y(n_8649)
);

CKINVDCx5p33_ASAP7_75t_R g8650 ( 
.A(n_8101),
.Y(n_8650)
);

BUFx6f_ASAP7_75t_L g8651 ( 
.A(n_7727),
.Y(n_8651)
);

AND2x2_ASAP7_75t_L g8652 ( 
.A(n_8085),
.B(n_6397),
.Y(n_8652)
);

CKINVDCx5p33_ASAP7_75t_R g8653 ( 
.A(n_7955),
.Y(n_8653)
);

CKINVDCx5p33_ASAP7_75t_R g8654 ( 
.A(n_8075),
.Y(n_8654)
);

BUFx2_ASAP7_75t_L g8655 ( 
.A(n_7875),
.Y(n_8655)
);

BUFx6f_ASAP7_75t_L g8656 ( 
.A(n_7731),
.Y(n_8656)
);

INVxp67_ASAP7_75t_L g8657 ( 
.A(n_8105),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8165),
.Y(n_8658)
);

INVx1_ASAP7_75t_L g8659 ( 
.A(n_7852),
.Y(n_8659)
);

BUFx6f_ASAP7_75t_L g8660 ( 
.A(n_7736),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_7862),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_7897),
.Y(n_8662)
);

HB1xp67_ASAP7_75t_L g8663 ( 
.A(n_7902),
.Y(n_8663)
);

CKINVDCx8_ASAP7_75t_R g8664 ( 
.A(n_8075),
.Y(n_8664)
);

CKINVDCx20_ASAP7_75t_R g8665 ( 
.A(n_8123),
.Y(n_8665)
);

CKINVDCx5p33_ASAP7_75t_R g8666 ( 
.A(n_8110),
.Y(n_8666)
);

INVx2_ASAP7_75t_L g8667 ( 
.A(n_7864),
.Y(n_8667)
);

HB1xp67_ASAP7_75t_L g8668 ( 
.A(n_8060),
.Y(n_8668)
);

INVx4_ASAP7_75t_L g8669 ( 
.A(n_7814),
.Y(n_8669)
);

INVx1_ASAP7_75t_L g8670 ( 
.A(n_7936),
.Y(n_8670)
);

CKINVDCx5p33_ASAP7_75t_R g8671 ( 
.A(n_8110),
.Y(n_8671)
);

CKINVDCx5p33_ASAP7_75t_R g8672 ( 
.A(n_7866),
.Y(n_8672)
);

NAND2xp5_ASAP7_75t_L g8673 ( 
.A(n_7892),
.B(n_5478),
.Y(n_8673)
);

INVx1_ASAP7_75t_L g8674 ( 
.A(n_7810),
.Y(n_8674)
);

INVx2_ASAP7_75t_L g8675 ( 
.A(n_7871),
.Y(n_8675)
);

INVx3_ASAP7_75t_L g8676 ( 
.A(n_7744),
.Y(n_8676)
);

CKINVDCx5p33_ASAP7_75t_R g8677 ( 
.A(n_7866),
.Y(n_8677)
);

BUFx6f_ASAP7_75t_L g8678 ( 
.A(n_7882),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_SL g8679 ( 
.A(n_7639),
.B(n_5480),
.Y(n_8679)
);

NAND2xp5_ASAP7_75t_L g8680 ( 
.A(n_7895),
.B(n_5487),
.Y(n_8680)
);

CKINVDCx5p33_ASAP7_75t_R g8681 ( 
.A(n_8121),
.Y(n_8681)
);

CKINVDCx5p33_ASAP7_75t_R g8682 ( 
.A(n_7986),
.Y(n_8682)
);

CKINVDCx20_ASAP7_75t_R g8683 ( 
.A(n_7704),
.Y(n_8683)
);

BUFx2_ASAP7_75t_L g8684 ( 
.A(n_7891),
.Y(n_8684)
);

INVx4_ASAP7_75t_L g8685 ( 
.A(n_7883),
.Y(n_8685)
);

INVx1_ASAP7_75t_L g8686 ( 
.A(n_7819),
.Y(n_8686)
);

CKINVDCx20_ASAP7_75t_R g8687 ( 
.A(n_8050),
.Y(n_8687)
);

NAND2xp5_ASAP7_75t_L g8688 ( 
.A(n_7903),
.B(n_7923),
.Y(n_8688)
);

INVx1_ASAP7_75t_SL g8689 ( 
.A(n_8088),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_7825),
.Y(n_8690)
);

INVx1_ASAP7_75t_L g8691 ( 
.A(n_7835),
.Y(n_8691)
);

INVx1_ASAP7_75t_L g8692 ( 
.A(n_7679),
.Y(n_8692)
);

CKINVDCx5p33_ASAP7_75t_R g8693 ( 
.A(n_7617),
.Y(n_8693)
);

INVx2_ASAP7_75t_L g8694 ( 
.A(n_7915),
.Y(n_8694)
);

INVx2_ASAP7_75t_L g8695 ( 
.A(n_7925),
.Y(n_8695)
);

NAND2xp5_ASAP7_75t_L g8696 ( 
.A(n_7933),
.B(n_5491),
.Y(n_8696)
);

CKINVDCx5p33_ASAP7_75t_R g8697 ( 
.A(n_7617),
.Y(n_8697)
);

NAND2xp33_ASAP7_75t_R g8698 ( 
.A(n_8108),
.B(n_5492),
.Y(n_8698)
);

INVx3_ASAP7_75t_L g8699 ( 
.A(n_7927),
.Y(n_8699)
);

CKINVDCx5p33_ASAP7_75t_R g8700 ( 
.A(n_7665),
.Y(n_8700)
);

AND2x4_ASAP7_75t_L g8701 ( 
.A(n_7805),
.B(n_5404),
.Y(n_8701)
);

INVx3_ASAP7_75t_L g8702 ( 
.A(n_7939),
.Y(n_8702)
);

INVx2_ASAP7_75t_L g8703 ( 
.A(n_7942),
.Y(n_8703)
);

NAND2xp5_ASAP7_75t_L g8704 ( 
.A(n_7968),
.B(n_5493),
.Y(n_8704)
);

CKINVDCx20_ASAP7_75t_R g8705 ( 
.A(n_8055),
.Y(n_8705)
);

CKINVDCx20_ASAP7_75t_R g8706 ( 
.A(n_8057),
.Y(n_8706)
);

BUFx6f_ASAP7_75t_L g8707 ( 
.A(n_7952),
.Y(n_8707)
);

INVx2_ASAP7_75t_L g8708 ( 
.A(n_7965),
.Y(n_8708)
);

INVx1_ASAP7_75t_L g8709 ( 
.A(n_7926),
.Y(n_8709)
);

NOR2xp33_ASAP7_75t_L g8710 ( 
.A(n_7959),
.B(n_5494),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_7969),
.Y(n_8711)
);

CKINVDCx20_ASAP7_75t_R g8712 ( 
.A(n_7826),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_7975),
.Y(n_8713)
);

INVx1_ASAP7_75t_L g8714 ( 
.A(n_7988),
.Y(n_8714)
);

AND2x2_ASAP7_75t_L g8715 ( 
.A(n_8133),
.B(n_6397),
.Y(n_8715)
);

NAND2xp5_ASAP7_75t_SL g8716 ( 
.A(n_7991),
.B(n_5497),
.Y(n_8716)
);

AND2x4_ASAP7_75t_L g8717 ( 
.A(n_7846),
.B(n_7984),
.Y(n_8717)
);

NAND2xp5_ASAP7_75t_L g8718 ( 
.A(n_7790),
.B(n_5504),
.Y(n_8718)
);

CKINVDCx5p33_ASAP7_75t_R g8719 ( 
.A(n_7665),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_8009),
.Y(n_8720)
);

INVx1_ASAP7_75t_SL g8721 ( 
.A(n_8004),
.Y(n_8721)
);

NOR2xp33_ASAP7_75t_L g8722 ( 
.A(n_7664),
.B(n_5509),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_7667),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8054),
.Y(n_8724)
);

CKINVDCx5p33_ASAP7_75t_R g8725 ( 
.A(n_7924),
.Y(n_8725)
);

INVx3_ASAP7_75t_L g8726 ( 
.A(n_7768),
.Y(n_8726)
);

INVx2_ASAP7_75t_L g8727 ( 
.A(n_7716),
.Y(n_8727)
);

CKINVDCx5p33_ASAP7_75t_R g8728 ( 
.A(n_7891),
.Y(n_8728)
);

INVx2_ASAP7_75t_L g8729 ( 
.A(n_7771),
.Y(n_8729)
);

INVx2_ASAP7_75t_L g8730 ( 
.A(n_7783),
.Y(n_8730)
);

INVx1_ASAP7_75t_L g8731 ( 
.A(n_7985),
.Y(n_8731)
);

AND2x4_ASAP7_75t_L g8732 ( 
.A(n_8020),
.B(n_5406),
.Y(n_8732)
);

CKINVDCx20_ASAP7_75t_R g8733 ( 
.A(n_7904),
.Y(n_8733)
);

HB1xp67_ASAP7_75t_L g8734 ( 
.A(n_7869),
.Y(n_8734)
);

CKINVDCx5p33_ASAP7_75t_R g8735 ( 
.A(n_7647),
.Y(n_8735)
);

INVx1_ASAP7_75t_L g8736 ( 
.A(n_7872),
.Y(n_8736)
);

NAND2xp33_ASAP7_75t_L g8737 ( 
.A(n_8116),
.B(n_5511),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_7918),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_L g8739 ( 
.A(n_7796),
.B(n_5518),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_7954),
.Y(n_8740)
);

CKINVDCx20_ASAP7_75t_R g8741 ( 
.A(n_7929),
.Y(n_8741)
);

OA21x2_ASAP7_75t_L g8742 ( 
.A1(n_7655),
.A2(n_5420),
.B(n_5411),
.Y(n_8742)
);

AND2x4_ASAP7_75t_L g8743 ( 
.A(n_7614),
.B(n_5425),
.Y(n_8743)
);

INVx1_ASAP7_75t_L g8744 ( 
.A(n_7797),
.Y(n_8744)
);

INVx1_ASAP7_75t_L g8745 ( 
.A(n_7628),
.Y(n_8745)
);

INVx1_ASAP7_75t_L g8746 ( 
.A(n_7668),
.Y(n_8746)
);

INVx2_ASAP7_75t_L g8747 ( 
.A(n_7674),
.Y(n_8747)
);

CKINVDCx5p33_ASAP7_75t_R g8748 ( 
.A(n_8162),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_7682),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_7774),
.Y(n_8750)
);

INVx2_ASAP7_75t_L g8751 ( 
.A(n_7935),
.Y(n_8751)
);

AND2x2_ASAP7_75t_L g8752 ( 
.A(n_8183),
.B(n_6422),
.Y(n_8752)
);

BUFx3_ASAP7_75t_L g8753 ( 
.A(n_7809),
.Y(n_8753)
);

INVx1_ASAP7_75t_L g8754 ( 
.A(n_7740),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_7858),
.Y(n_8755)
);

CKINVDCx5p33_ASAP7_75t_R g8756 ( 
.A(n_7626),
.Y(n_8756)
);

INVx1_ASAP7_75t_L g8757 ( 
.A(n_7956),
.Y(n_8757)
);

NAND2xp5_ASAP7_75t_L g8758 ( 
.A(n_8526),
.B(n_7613),
.Y(n_8758)
);

INVx2_ASAP7_75t_L g8759 ( 
.A(n_8205),
.Y(n_8759)
);

INVx2_ASAP7_75t_L g8760 ( 
.A(n_8207),
.Y(n_8760)
);

INVx2_ASAP7_75t_L g8761 ( 
.A(n_8224),
.Y(n_8761)
);

INVx2_ASAP7_75t_L g8762 ( 
.A(n_8235),
.Y(n_8762)
);

NAND2xp5_ASAP7_75t_SL g8763 ( 
.A(n_8692),
.B(n_8002),
.Y(n_8763)
);

INVx1_ASAP7_75t_SL g8764 ( 
.A(n_8352),
.Y(n_8764)
);

AND2x4_ASAP7_75t_L g8765 ( 
.A(n_8309),
.B(n_7747),
.Y(n_8765)
);

OAI21xp5_ASAP7_75t_L g8766 ( 
.A1(n_8636),
.A2(n_7661),
.B(n_7624),
.Y(n_8766)
);

INVx1_ASAP7_75t_L g8767 ( 
.A(n_8200),
.Y(n_8767)
);

INVx2_ASAP7_75t_L g8768 ( 
.A(n_8242),
.Y(n_8768)
);

AND3x2_ASAP7_75t_L g8769 ( 
.A(n_8458),
.B(n_5432),
.C(n_5427),
.Y(n_8769)
);

NAND2xp5_ASAP7_75t_L g8770 ( 
.A(n_8570),
.B(n_7912),
.Y(n_8770)
);

INVx2_ASAP7_75t_L g8771 ( 
.A(n_8202),
.Y(n_8771)
);

INVx1_ASAP7_75t_L g8772 ( 
.A(n_8209),
.Y(n_8772)
);

INVx1_ASAP7_75t_L g8773 ( 
.A(n_8215),
.Y(n_8773)
);

BUFx2_ASAP7_75t_L g8774 ( 
.A(n_8230),
.Y(n_8774)
);

NAND2xp5_ASAP7_75t_L g8775 ( 
.A(n_8688),
.B(n_7934),
.Y(n_8775)
);

INVx1_ASAP7_75t_SL g8776 ( 
.A(n_8389),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_SL g8777 ( 
.A(n_8433),
.B(n_8011),
.Y(n_8777)
);

INVx2_ASAP7_75t_L g8778 ( 
.A(n_8216),
.Y(n_8778)
);

NAND2xp5_ASAP7_75t_SL g8779 ( 
.A(n_8195),
.B(n_7766),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_8218),
.Y(n_8780)
);

NAND3xp33_ASAP7_75t_L g8781 ( 
.A(n_8274),
.B(n_7640),
.C(n_7782),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_SL g8782 ( 
.A(n_8436),
.B(n_6612),
.Y(n_8782)
);

INVx1_ASAP7_75t_L g8783 ( 
.A(n_8220),
.Y(n_8783)
);

BUFx6f_ASAP7_75t_L g8784 ( 
.A(n_8270),
.Y(n_8784)
);

INVx1_ASAP7_75t_L g8785 ( 
.A(n_8222),
.Y(n_8785)
);

NAND2xp5_ASAP7_75t_L g8786 ( 
.A(n_8744),
.B(n_5521),
.Y(n_8786)
);

NAND2xp5_ASAP7_75t_SL g8787 ( 
.A(n_8564),
.B(n_6615),
.Y(n_8787)
);

OAI22xp5_ASAP7_75t_L g8788 ( 
.A1(n_8674),
.A2(n_5526),
.B1(n_5528),
.B2(n_5524),
.Y(n_8788)
);

AND2x2_ASAP7_75t_L g8789 ( 
.A(n_8240),
.B(n_6422),
.Y(n_8789)
);

INVx2_ASAP7_75t_L g8790 ( 
.A(n_8223),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_8225),
.Y(n_8791)
);

INVx8_ASAP7_75t_L g8792 ( 
.A(n_8484),
.Y(n_8792)
);

INVx4_ASAP7_75t_L g8793 ( 
.A(n_8310),
.Y(n_8793)
);

CKINVDCx5p33_ASAP7_75t_R g8794 ( 
.A(n_8201),
.Y(n_8794)
);

INVx6_ASAP7_75t_L g8795 ( 
.A(n_8359),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_SL g8796 ( 
.A(n_8576),
.B(n_5532),
.Y(n_8796)
);

BUFx6f_ASAP7_75t_L g8797 ( 
.A(n_8270),
.Y(n_8797)
);

INVx2_ASAP7_75t_L g8798 ( 
.A(n_8227),
.Y(n_8798)
);

INVx1_ASAP7_75t_L g8799 ( 
.A(n_8238),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_8245),
.Y(n_8800)
);

INVx2_ASAP7_75t_L g8801 ( 
.A(n_8246),
.Y(n_8801)
);

INVx2_ASAP7_75t_L g8802 ( 
.A(n_8251),
.Y(n_8802)
);

INVx2_ASAP7_75t_L g8803 ( 
.A(n_8258),
.Y(n_8803)
);

NAND2xp5_ASAP7_75t_SL g8804 ( 
.A(n_8577),
.B(n_8578),
.Y(n_8804)
);

NAND2xp5_ASAP7_75t_L g8805 ( 
.A(n_8631),
.B(n_5538),
.Y(n_8805)
);

INVx2_ASAP7_75t_L g8806 ( 
.A(n_8262),
.Y(n_8806)
);

AND3x2_ASAP7_75t_L g8807 ( 
.A(n_8492),
.B(n_8527),
.C(n_8535),
.Y(n_8807)
);

AOI22xp33_ASAP7_75t_L g8808 ( 
.A1(n_8722),
.A2(n_6291),
.B1(n_6319),
.B2(n_6229),
.Y(n_8808)
);

INVx1_ASAP7_75t_L g8809 ( 
.A(n_8265),
.Y(n_8809)
);

NAND2xp5_ASAP7_75t_SL g8810 ( 
.A(n_8580),
.B(n_5540),
.Y(n_8810)
);

BUFx3_ASAP7_75t_L g8811 ( 
.A(n_8474),
.Y(n_8811)
);

INVx3_ASAP7_75t_L g8812 ( 
.A(n_8678),
.Y(n_8812)
);

AO21x2_ASAP7_75t_L g8813 ( 
.A1(n_8724),
.A2(n_8641),
.B(n_8639),
.Y(n_8813)
);

INVx2_ASAP7_75t_L g8814 ( 
.A(n_8267),
.Y(n_8814)
);

NAND2xp5_ASAP7_75t_SL g8815 ( 
.A(n_8591),
.B(n_5541),
.Y(n_8815)
);

NAND2xp5_ASAP7_75t_L g8816 ( 
.A(n_8634),
.B(n_5544),
.Y(n_8816)
);

INVx2_ASAP7_75t_L g8817 ( 
.A(n_8269),
.Y(n_8817)
);

INVx2_ASAP7_75t_L g8818 ( 
.A(n_8280),
.Y(n_8818)
);

INVx3_ASAP7_75t_L g8819 ( 
.A(n_8678),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_SL g8820 ( 
.A(n_8594),
.B(n_5545),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_L g8821 ( 
.A(n_8563),
.B(n_5547),
.Y(n_8821)
);

NAND2xp5_ASAP7_75t_L g8822 ( 
.A(n_8339),
.B(n_8350),
.Y(n_8822)
);

INVx2_ASAP7_75t_L g8823 ( 
.A(n_8281),
.Y(n_8823)
);

INVx2_ASAP7_75t_L g8824 ( 
.A(n_8288),
.Y(n_8824)
);

INVx2_ASAP7_75t_L g8825 ( 
.A(n_8290),
.Y(n_8825)
);

AOI21x1_ASAP7_75t_L g8826 ( 
.A1(n_8566),
.A2(n_5435),
.B(n_5434),
.Y(n_8826)
);

BUFx3_ASAP7_75t_L g8827 ( 
.A(n_8226),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_8297),
.Y(n_8828)
);

INVx2_ASAP7_75t_L g8829 ( 
.A(n_8298),
.Y(n_8829)
);

INVx2_ASAP7_75t_SL g8830 ( 
.A(n_8323),
.Y(n_8830)
);

NAND2xp5_ASAP7_75t_L g8831 ( 
.A(n_8388),
.B(n_5550),
.Y(n_8831)
);

INVx2_ASAP7_75t_L g8832 ( 
.A(n_8304),
.Y(n_8832)
);

INVx1_ASAP7_75t_L g8833 ( 
.A(n_8305),
.Y(n_8833)
);

AND2x4_ASAP7_75t_L g8834 ( 
.A(n_8204),
.B(n_5442),
.Y(n_8834)
);

NAND2xp5_ASAP7_75t_SL g8835 ( 
.A(n_8344),
.B(n_5552),
.Y(n_8835)
);

OR2x6_ASAP7_75t_L g8836 ( 
.A(n_8221),
.B(n_5443),
.Y(n_8836)
);

INVx2_ASAP7_75t_L g8837 ( 
.A(n_8315),
.Y(n_8837)
);

INVx2_ASAP7_75t_SL g8838 ( 
.A(n_8328),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_8319),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_8322),
.Y(n_8840)
);

BUFx2_ASAP7_75t_L g8841 ( 
.A(n_8602),
.Y(n_8841)
);

NOR2xp33_ASAP7_75t_L g8842 ( 
.A(n_8212),
.B(n_7756),
.Y(n_8842)
);

INVx2_ASAP7_75t_L g8843 ( 
.A(n_8331),
.Y(n_8843)
);

NAND2xp5_ASAP7_75t_L g8844 ( 
.A(n_8565),
.B(n_8686),
.Y(n_8844)
);

INVx2_ASAP7_75t_L g8845 ( 
.A(n_8337),
.Y(n_8845)
);

INVx3_ASAP7_75t_L g8846 ( 
.A(n_8707),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_8338),
.Y(n_8847)
);

NAND3xp33_ASAP7_75t_L g8848 ( 
.A(n_8601),
.B(n_8111),
.C(n_8053),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_8355),
.Y(n_8849)
);

INVx2_ASAP7_75t_L g8850 ( 
.A(n_8361),
.Y(n_8850)
);

NAND2xp33_ASAP7_75t_L g8851 ( 
.A(n_8402),
.B(n_5553),
.Y(n_8851)
);

BUFx6f_ASAP7_75t_L g8852 ( 
.A(n_8303),
.Y(n_8852)
);

INVx2_ASAP7_75t_L g8853 ( 
.A(n_8365),
.Y(n_8853)
);

INVx2_ASAP7_75t_L g8854 ( 
.A(n_8368),
.Y(n_8854)
);

INVx2_ASAP7_75t_L g8855 ( 
.A(n_8373),
.Y(n_8855)
);

NAND2xp5_ASAP7_75t_L g8856 ( 
.A(n_8690),
.B(n_5554),
.Y(n_8856)
);

BUFx3_ASAP7_75t_L g8857 ( 
.A(n_8226),
.Y(n_8857)
);

INVx1_ASAP7_75t_L g8858 ( 
.A(n_8376),
.Y(n_8858)
);

NOR2xp33_ASAP7_75t_L g8859 ( 
.A(n_8197),
.B(n_7922),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_8377),
.Y(n_8860)
);

INVxp33_ASAP7_75t_SL g8861 ( 
.A(n_8210),
.Y(n_8861)
);

INVx2_ASAP7_75t_L g8862 ( 
.A(n_8378),
.Y(n_8862)
);

NOR2xp33_ASAP7_75t_L g8863 ( 
.A(n_8394),
.B(n_8129),
.Y(n_8863)
);

NAND2xp5_ASAP7_75t_SL g8864 ( 
.A(n_8538),
.B(n_8542),
.Y(n_8864)
);

INVx1_ASAP7_75t_L g8865 ( 
.A(n_8380),
.Y(n_8865)
);

INVx2_ASAP7_75t_L g8866 ( 
.A(n_8382),
.Y(n_8866)
);

INVx1_ASAP7_75t_L g8867 ( 
.A(n_8383),
.Y(n_8867)
);

INVx3_ASAP7_75t_L g8868 ( 
.A(n_8707),
.Y(n_8868)
);

INVx1_ASAP7_75t_L g8869 ( 
.A(n_8387),
.Y(n_8869)
);

INVx1_ASAP7_75t_L g8870 ( 
.A(n_8391),
.Y(n_8870)
);

INVx2_ASAP7_75t_L g8871 ( 
.A(n_8406),
.Y(n_8871)
);

NOR2xp33_ASAP7_75t_L g8872 ( 
.A(n_8417),
.B(n_8189),
.Y(n_8872)
);

INVx2_ASAP7_75t_L g8873 ( 
.A(n_8411),
.Y(n_8873)
);

NOR2xp33_ASAP7_75t_L g8874 ( 
.A(n_8460),
.B(n_5555),
.Y(n_8874)
);

NAND2xp5_ASAP7_75t_L g8875 ( 
.A(n_8691),
.B(n_5557),
.Y(n_8875)
);

INVx2_ASAP7_75t_L g8876 ( 
.A(n_8420),
.Y(n_8876)
);

INVx2_ASAP7_75t_L g8877 ( 
.A(n_8426),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_L g8878 ( 
.A(n_8534),
.B(n_5560),
.Y(n_8878)
);

INVx3_ASAP7_75t_L g8879 ( 
.A(n_8517),
.Y(n_8879)
);

NOR2xp33_ASAP7_75t_L g8880 ( 
.A(n_8550),
.B(n_5564),
.Y(n_8880)
);

INVx4_ASAP7_75t_L g8881 ( 
.A(n_8311),
.Y(n_8881)
);

NAND2xp5_ASAP7_75t_SL g8882 ( 
.A(n_8556),
.B(n_5565),
.Y(n_8882)
);

INVx2_ASAP7_75t_L g8883 ( 
.A(n_8428),
.Y(n_8883)
);

OR2x2_ASAP7_75t_L g8884 ( 
.A(n_8541),
.B(n_5566),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8432),
.Y(n_8885)
);

INVx1_ASAP7_75t_L g8886 ( 
.A(n_8434),
.Y(n_8886)
);

INVx1_ASAP7_75t_L g8887 ( 
.A(n_8446),
.Y(n_8887)
);

BUFx3_ASAP7_75t_L g8888 ( 
.A(n_8483),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8461),
.Y(n_8889)
);

INVx1_ASAP7_75t_L g8890 ( 
.A(n_8464),
.Y(n_8890)
);

CKINVDCx5p33_ASAP7_75t_R g8891 ( 
.A(n_8211),
.Y(n_8891)
);

NAND2xp5_ASAP7_75t_L g8892 ( 
.A(n_8659),
.B(n_5569),
.Y(n_8892)
);

INVxp33_ASAP7_75t_L g8893 ( 
.A(n_8431),
.Y(n_8893)
);

BUFx6f_ASAP7_75t_L g8894 ( 
.A(n_8303),
.Y(n_8894)
);

INVx2_ASAP7_75t_L g8895 ( 
.A(n_8465),
.Y(n_8895)
);

AND2x2_ASAP7_75t_L g8896 ( 
.A(n_8469),
.B(n_8471),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_8476),
.Y(n_8897)
);

INVxp67_ASAP7_75t_SL g8898 ( 
.A(n_8449),
.Y(n_8898)
);

INVx2_ASAP7_75t_SL g8899 ( 
.A(n_8408),
.Y(n_8899)
);

OAI22xp5_ASAP7_75t_L g8900 ( 
.A1(n_8746),
.A2(n_5577),
.B1(n_5578),
.B2(n_5573),
.Y(n_8900)
);

NAND2xp5_ASAP7_75t_SL g8901 ( 
.A(n_8620),
.B(n_5580),
.Y(n_8901)
);

INVx2_ASAP7_75t_L g8902 ( 
.A(n_8479),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_SL g8903 ( 
.A(n_8630),
.B(n_8637),
.Y(n_8903)
);

NAND2xp5_ASAP7_75t_SL g8904 ( 
.A(n_8638),
.B(n_5582),
.Y(n_8904)
);

INVx2_ASAP7_75t_L g8905 ( 
.A(n_8489),
.Y(n_8905)
);

INVx1_ASAP7_75t_L g8906 ( 
.A(n_8490),
.Y(n_8906)
);

BUFx6f_ASAP7_75t_L g8907 ( 
.A(n_8347),
.Y(n_8907)
);

NOR2xp33_ASAP7_75t_L g8908 ( 
.A(n_8466),
.B(n_5585),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8493),
.Y(n_8909)
);

NAND2xp33_ASAP7_75t_L g8910 ( 
.A(n_8403),
.B(n_5588),
.Y(n_8910)
);

CKINVDCx6p67_ASAP7_75t_R g8911 ( 
.A(n_8495),
.Y(n_8911)
);

NAND2xp5_ASAP7_75t_L g8912 ( 
.A(n_8501),
.B(n_5589),
.Y(n_8912)
);

NOR2xp33_ASAP7_75t_L g8913 ( 
.A(n_8198),
.B(n_5590),
.Y(n_8913)
);

NOR2xp33_ASAP7_75t_L g8914 ( 
.A(n_8360),
.B(n_5592),
.Y(n_8914)
);

NAND2xp5_ASAP7_75t_L g8915 ( 
.A(n_8521),
.B(n_5593),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_8494),
.Y(n_8916)
);

INVx2_ASAP7_75t_L g8917 ( 
.A(n_8568),
.Y(n_8917)
);

INVx2_ASAP7_75t_L g8918 ( 
.A(n_8571),
.Y(n_8918)
);

INVx2_ASAP7_75t_L g8919 ( 
.A(n_8581),
.Y(n_8919)
);

NAND2xp5_ASAP7_75t_L g8920 ( 
.A(n_8231),
.B(n_5596),
.Y(n_8920)
);

AOI22xp33_ASAP7_75t_L g8921 ( 
.A1(n_8749),
.A2(n_8755),
.B1(n_8757),
.B2(n_8754),
.Y(n_8921)
);

INVx2_ASAP7_75t_SL g8922 ( 
.A(n_8424),
.Y(n_8922)
);

NAND3xp33_ASAP7_75t_L g8923 ( 
.A(n_8569),
.B(n_8710),
.C(n_8203),
.Y(n_8923)
);

INVx2_ASAP7_75t_L g8924 ( 
.A(n_8584),
.Y(n_8924)
);

BUFx10_ASAP7_75t_L g8925 ( 
.A(n_8213),
.Y(n_8925)
);

BUFx3_ASAP7_75t_L g8926 ( 
.A(n_8597),
.Y(n_8926)
);

NOR2xp33_ASAP7_75t_L g8927 ( 
.A(n_8657),
.B(n_5597),
.Y(n_8927)
);

INVx2_ASAP7_75t_L g8928 ( 
.A(n_8592),
.Y(n_8928)
);

INVx3_ASAP7_75t_L g8929 ( 
.A(n_8517),
.Y(n_8929)
);

CKINVDCx6p67_ASAP7_75t_R g8930 ( 
.A(n_8496),
.Y(n_8930)
);

NOR2xp33_ASAP7_75t_L g8931 ( 
.A(n_8663),
.B(n_5598),
.Y(n_8931)
);

INVx1_ASAP7_75t_L g8932 ( 
.A(n_8498),
.Y(n_8932)
);

INVx2_ASAP7_75t_L g8933 ( 
.A(n_8600),
.Y(n_8933)
);

NAND2xp5_ASAP7_75t_L g8934 ( 
.A(n_8599),
.B(n_5600),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8603),
.B(n_5601),
.Y(n_8935)
);

INVx2_ASAP7_75t_L g8936 ( 
.A(n_8608),
.Y(n_8936)
);

NAND2xp5_ASAP7_75t_L g8937 ( 
.A(n_8607),
.B(n_5602),
.Y(n_8937)
);

INVx2_ASAP7_75t_L g8938 ( 
.A(n_8499),
.Y(n_8938)
);

INVx2_ASAP7_75t_L g8939 ( 
.A(n_8503),
.Y(n_8939)
);

INVx1_ASAP7_75t_L g8940 ( 
.A(n_8504),
.Y(n_8940)
);

INVx2_ASAP7_75t_L g8941 ( 
.A(n_8314),
.Y(n_8941)
);

NAND2xp5_ASAP7_75t_SL g8942 ( 
.A(n_8646),
.B(n_5607),
.Y(n_8942)
);

NAND2xp5_ASAP7_75t_L g8943 ( 
.A(n_8648),
.B(n_5608),
.Y(n_8943)
);

INVx1_ASAP7_75t_L g8944 ( 
.A(n_8514),
.Y(n_8944)
);

INVx2_ASAP7_75t_L g8945 ( 
.A(n_8317),
.Y(n_8945)
);

NOR2xp33_ASAP7_75t_L g8946 ( 
.A(n_8429),
.B(n_5609),
.Y(n_8946)
);

INVx1_ASAP7_75t_L g8947 ( 
.A(n_8523),
.Y(n_8947)
);

INVx2_ASAP7_75t_SL g8948 ( 
.A(n_8467),
.Y(n_8948)
);

INVx2_ASAP7_75t_L g8949 ( 
.A(n_8320),
.Y(n_8949)
);

OAI22xp33_ASAP7_75t_SL g8950 ( 
.A1(n_8283),
.A2(n_5447),
.B1(n_5455),
.B2(n_5444),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_SL g8951 ( 
.A(n_8647),
.B(n_5610),
.Y(n_8951)
);

BUFx10_ASAP7_75t_L g8952 ( 
.A(n_8214),
.Y(n_8952)
);

NAND2xp5_ASAP7_75t_L g8953 ( 
.A(n_8673),
.B(n_5614),
.Y(n_8953)
);

OAI22xp33_ASAP7_75t_L g8954 ( 
.A1(n_8745),
.A2(n_5625),
.B1(n_5626),
.B2(n_5622),
.Y(n_8954)
);

INVx2_ASAP7_75t_L g8955 ( 
.A(n_8321),
.Y(n_8955)
);

INVx1_ASAP7_75t_L g8956 ( 
.A(n_8528),
.Y(n_8956)
);

INVx2_ASAP7_75t_L g8957 ( 
.A(n_8325),
.Y(n_8957)
);

INVx3_ASAP7_75t_L g8958 ( 
.A(n_8522),
.Y(n_8958)
);

NAND2xp5_ASAP7_75t_SL g8959 ( 
.A(n_8650),
.B(n_5627),
.Y(n_8959)
);

INVx2_ASAP7_75t_L g8960 ( 
.A(n_8343),
.Y(n_8960)
);

NAND2xp5_ASAP7_75t_L g8961 ( 
.A(n_8680),
.B(n_5628),
.Y(n_8961)
);

BUFx10_ASAP7_75t_L g8962 ( 
.A(n_8217),
.Y(n_8962)
);

INVx2_ASAP7_75t_SL g8963 ( 
.A(n_8199),
.Y(n_8963)
);

INVx1_ASAP7_75t_L g8964 ( 
.A(n_8531),
.Y(n_8964)
);

NOR2xp33_ASAP7_75t_L g8965 ( 
.A(n_8653),
.B(n_5630),
.Y(n_8965)
);

INVx2_ASAP7_75t_L g8966 ( 
.A(n_8346),
.Y(n_8966)
);

NAND3xp33_ASAP7_75t_L g8967 ( 
.A(n_8412),
.B(n_5635),
.C(n_5633),
.Y(n_8967)
);

INVx2_ASAP7_75t_L g8968 ( 
.A(n_8358),
.Y(n_8968)
);

INVx3_ASAP7_75t_L g8969 ( 
.A(n_8522),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_8536),
.Y(n_8970)
);

NAND2xp5_ASAP7_75t_L g8971 ( 
.A(n_8696),
.B(n_5638),
.Y(n_8971)
);

INVx2_ASAP7_75t_L g8972 ( 
.A(n_8366),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8540),
.Y(n_8973)
);

AOI21x1_ASAP7_75t_L g8974 ( 
.A1(n_8643),
.A2(n_5457),
.B(n_5456),
.Y(n_8974)
);

INVx1_ASAP7_75t_L g8975 ( 
.A(n_8545),
.Y(n_8975)
);

INVx2_ASAP7_75t_L g8976 ( 
.A(n_8372),
.Y(n_8976)
);

INVx2_ASAP7_75t_L g8977 ( 
.A(n_8385),
.Y(n_8977)
);

INVx2_ASAP7_75t_L g8978 ( 
.A(n_8404),
.Y(n_8978)
);

BUFx6f_ASAP7_75t_L g8979 ( 
.A(n_8347),
.Y(n_8979)
);

INVx2_ASAP7_75t_SL g8980 ( 
.A(n_8453),
.Y(n_8980)
);

NAND3xp33_ASAP7_75t_L g8981 ( 
.A(n_8363),
.B(n_5642),
.C(n_5641),
.Y(n_8981)
);

BUFx10_ASAP7_75t_L g8982 ( 
.A(n_8228),
.Y(n_8982)
);

INVx2_ASAP7_75t_L g8983 ( 
.A(n_8416),
.Y(n_8983)
);

NAND2xp5_ASAP7_75t_SL g8984 ( 
.A(n_8405),
.B(n_5643),
.Y(n_8984)
);

INVx2_ASAP7_75t_L g8985 ( 
.A(n_8422),
.Y(n_8985)
);

AND2x2_ASAP7_75t_L g8986 ( 
.A(n_8336),
.B(n_6435),
.Y(n_8986)
);

INVx5_ASAP7_75t_L g8987 ( 
.A(n_8397),
.Y(n_8987)
);

INVx3_ASAP7_75t_L g8988 ( 
.A(n_8561),
.Y(n_8988)
);

OR2x6_ASAP7_75t_L g8989 ( 
.A(n_8430),
.B(n_5460),
.Y(n_8989)
);

BUFx3_ASAP7_75t_L g8990 ( 
.A(n_8349),
.Y(n_8990)
);

INVx2_ASAP7_75t_L g8991 ( 
.A(n_8442),
.Y(n_8991)
);

BUFx3_ASAP7_75t_L g8992 ( 
.A(n_8379),
.Y(n_8992)
);

NAND2xp5_ASAP7_75t_SL g8993 ( 
.A(n_8409),
.B(n_5649),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8444),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_8551),
.Y(n_8995)
);

INVx2_ASAP7_75t_L g8996 ( 
.A(n_8445),
.Y(n_8996)
);

INVx2_ASAP7_75t_L g8997 ( 
.A(n_8454),
.Y(n_8997)
);

BUFx3_ASAP7_75t_L g8998 ( 
.A(n_8384),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_8557),
.Y(n_8999)
);

INVx1_ASAP7_75t_L g9000 ( 
.A(n_8560),
.Y(n_9000)
);

NAND2xp5_ASAP7_75t_L g9001 ( 
.A(n_8704),
.B(n_5652),
.Y(n_9001)
);

NAND2xp5_ASAP7_75t_L g9002 ( 
.A(n_8718),
.B(n_5660),
.Y(n_9002)
);

INVx2_ASAP7_75t_SL g9003 ( 
.A(n_8293),
.Y(n_9003)
);

INVx2_ASAP7_75t_L g9004 ( 
.A(n_8475),
.Y(n_9004)
);

BUFx6f_ASAP7_75t_L g9005 ( 
.A(n_8353),
.Y(n_9005)
);

CKINVDCx5p33_ASAP7_75t_R g9006 ( 
.A(n_8232),
.Y(n_9006)
);

INVx1_ASAP7_75t_L g9007 ( 
.A(n_8562),
.Y(n_9007)
);

NOR2xp33_ASAP7_75t_L g9008 ( 
.A(n_8548),
.B(n_5661),
.Y(n_9008)
);

INVx3_ASAP7_75t_L g9009 ( 
.A(n_8561),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8574),
.Y(n_9010)
);

INVx2_ASAP7_75t_L g9011 ( 
.A(n_8478),
.Y(n_9011)
);

INVx2_ASAP7_75t_L g9012 ( 
.A(n_8500),
.Y(n_9012)
);

INVx2_ASAP7_75t_L g9013 ( 
.A(n_8512),
.Y(n_9013)
);

NOR2xp33_ASAP7_75t_L g9014 ( 
.A(n_8229),
.B(n_5666),
.Y(n_9014)
);

BUFx10_ASAP7_75t_L g9015 ( 
.A(n_8237),
.Y(n_9015)
);

INVx2_ASAP7_75t_L g9016 ( 
.A(n_8515),
.Y(n_9016)
);

INVx2_ASAP7_75t_L g9017 ( 
.A(n_8520),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_8575),
.Y(n_9018)
);

INVx2_ASAP7_75t_L g9019 ( 
.A(n_8525),
.Y(n_9019)
);

INVx2_ASAP7_75t_SL g9020 ( 
.A(n_8507),
.Y(n_9020)
);

NAND3xp33_ASAP7_75t_L g9021 ( 
.A(n_8206),
.B(n_5671),
.C(n_5667),
.Y(n_9021)
);

AND3x2_ASAP7_75t_L g9022 ( 
.A(n_8655),
.B(n_5463),
.C(n_5462),
.Y(n_9022)
);

INVx1_ASAP7_75t_L g9023 ( 
.A(n_8582),
.Y(n_9023)
);

INVx3_ASAP7_75t_L g9024 ( 
.A(n_8567),
.Y(n_9024)
);

INVx2_ASAP7_75t_L g9025 ( 
.A(n_8529),
.Y(n_9025)
);

INVx1_ASAP7_75t_L g9026 ( 
.A(n_8583),
.Y(n_9026)
);

INVx2_ASAP7_75t_L g9027 ( 
.A(n_8552),
.Y(n_9027)
);

AND2x6_ASAP7_75t_L g9028 ( 
.A(n_8662),
.B(n_5467),
.Y(n_9028)
);

INVx2_ASAP7_75t_L g9029 ( 
.A(n_8553),
.Y(n_9029)
);

INVx2_ASAP7_75t_L g9030 ( 
.A(n_8558),
.Y(n_9030)
);

INVxp67_ASAP7_75t_SL g9031 ( 
.A(n_8449),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8587),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_8588),
.Y(n_9033)
);

NAND2xp5_ASAP7_75t_L g9034 ( 
.A(n_8739),
.B(n_5674),
.Y(n_9034)
);

AND2x2_ASAP7_75t_L g9035 ( 
.A(n_8340),
.B(n_6435),
.Y(n_9035)
);

INVx2_ASAP7_75t_L g9036 ( 
.A(n_8244),
.Y(n_9036)
);

INVxp33_ASAP7_75t_L g9037 ( 
.A(n_8448),
.Y(n_9037)
);

INVx2_ASAP7_75t_L g9038 ( 
.A(n_8271),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8589),
.Y(n_9039)
);

NAND2xp5_ASAP7_75t_SL g9040 ( 
.A(n_8419),
.B(n_5681),
.Y(n_9040)
);

INVx2_ASAP7_75t_SL g9041 ( 
.A(n_8353),
.Y(n_9041)
);

NAND2xp5_ASAP7_75t_SL g9042 ( 
.A(n_8421),
.B(n_5686),
.Y(n_9042)
);

INVx2_ASAP7_75t_L g9043 ( 
.A(n_8272),
.Y(n_9043)
);

INVx11_ASAP7_75t_L g9044 ( 
.A(n_8518),
.Y(n_9044)
);

NAND2xp5_ASAP7_75t_L g9045 ( 
.A(n_8357),
.B(n_8364),
.Y(n_9045)
);

BUFx3_ASAP7_75t_L g9046 ( 
.A(n_8390),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8590),
.Y(n_9047)
);

INVx2_ASAP7_75t_L g9048 ( 
.A(n_8275),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_8287),
.Y(n_9049)
);

NAND2xp33_ASAP7_75t_L g9050 ( 
.A(n_8427),
.B(n_5694),
.Y(n_9050)
);

INVx2_ASAP7_75t_L g9051 ( 
.A(n_8291),
.Y(n_9051)
);

INVx1_ASAP7_75t_L g9052 ( 
.A(n_8593),
.Y(n_9052)
);

BUFx10_ASAP7_75t_L g9053 ( 
.A(n_8243),
.Y(n_9053)
);

OAI22xp33_ASAP7_75t_L g9054 ( 
.A1(n_8681),
.A2(n_5699),
.B1(n_5701),
.B2(n_5697),
.Y(n_9054)
);

INVx2_ASAP7_75t_L g9055 ( 
.A(n_8300),
.Y(n_9055)
);

AND2x4_ASAP7_75t_L g9056 ( 
.A(n_8516),
.B(n_5470),
.Y(n_9056)
);

NAND2xp5_ASAP7_75t_L g9057 ( 
.A(n_8410),
.B(n_5708),
.Y(n_9057)
);

INVx3_ASAP7_75t_L g9058 ( 
.A(n_8567),
.Y(n_9058)
);

NAND2xp5_ASAP7_75t_SL g9059 ( 
.A(n_8438),
.B(n_5713),
.Y(n_9059)
);

BUFx3_ASAP7_75t_L g9060 ( 
.A(n_8342),
.Y(n_9060)
);

INVx1_ASAP7_75t_L g9061 ( 
.A(n_8598),
.Y(n_9061)
);

NAND2xp5_ASAP7_75t_SL g9062 ( 
.A(n_8689),
.B(n_5715),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_SL g9063 ( 
.A(n_8617),
.B(n_8618),
.Y(n_9063)
);

INVxp67_ASAP7_75t_SL g9064 ( 
.A(n_8463),
.Y(n_9064)
);

INVx1_ASAP7_75t_L g9065 ( 
.A(n_8605),
.Y(n_9065)
);

BUFx6f_ASAP7_75t_L g9066 ( 
.A(n_8371),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8610),
.Y(n_9067)
);

INVx2_ASAP7_75t_L g9068 ( 
.A(n_8301),
.Y(n_9068)
);

NAND2xp5_ASAP7_75t_SL g9069 ( 
.A(n_8625),
.B(n_5718),
.Y(n_9069)
);

INVx1_ASAP7_75t_L g9070 ( 
.A(n_8612),
.Y(n_9070)
);

INVx1_ASAP7_75t_L g9071 ( 
.A(n_8613),
.Y(n_9071)
);

INVx2_ASAP7_75t_L g9072 ( 
.A(n_8615),
.Y(n_9072)
);

AOI22xp5_ASAP7_75t_L g9073 ( 
.A1(n_8447),
.A2(n_5723),
.B1(n_5724),
.B2(n_5720),
.Y(n_9073)
);

INVx2_ASAP7_75t_L g9074 ( 
.A(n_8616),
.Y(n_9074)
);

INVx3_ASAP7_75t_L g9075 ( 
.A(n_8614),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8252),
.Y(n_9076)
);

NAND2xp5_ASAP7_75t_SL g9077 ( 
.A(n_8626),
.B(n_5725),
.Y(n_9077)
);

INVx1_ASAP7_75t_L g9078 ( 
.A(n_8254),
.Y(n_9078)
);

NAND2xp5_ASAP7_75t_L g9079 ( 
.A(n_8532),
.B(n_5728),
.Y(n_9079)
);

INVx3_ASAP7_75t_L g9080 ( 
.A(n_8614),
.Y(n_9080)
);

INVx2_ASAP7_75t_L g9081 ( 
.A(n_8463),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8256),
.Y(n_9082)
);

BUFx4f_ASAP7_75t_L g9083 ( 
.A(n_8596),
.Y(n_9083)
);

INVx3_ASAP7_75t_L g9084 ( 
.A(n_8651),
.Y(n_9084)
);

AOI21x1_ASAP7_75t_L g9085 ( 
.A1(n_8658),
.A2(n_5473),
.B(n_5471),
.Y(n_9085)
);

NAND2xp5_ASAP7_75t_L g9086 ( 
.A(n_8539),
.B(n_5729),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8572),
.Y(n_9087)
);

INVx2_ASAP7_75t_L g9088 ( 
.A(n_8627),
.Y(n_9088)
);

NAND2xp5_ASAP7_75t_SL g9089 ( 
.A(n_8721),
.B(n_5731),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_8573),
.Y(n_9090)
);

BUFx2_ASAP7_75t_L g9091 ( 
.A(n_8621),
.Y(n_9091)
);

INVx2_ASAP7_75t_L g9092 ( 
.A(n_8628),
.Y(n_9092)
);

INVx1_ASAP7_75t_L g9093 ( 
.A(n_8619),
.Y(n_9093)
);

INVx2_ASAP7_75t_L g9094 ( 
.A(n_8640),
.Y(n_9094)
);

INVx2_ASAP7_75t_L g9095 ( 
.A(n_8642),
.Y(n_9095)
);

AND2x4_ASAP7_75t_L g9096 ( 
.A(n_8633),
.B(n_5481),
.Y(n_9096)
);

BUFx3_ASAP7_75t_L g9097 ( 
.A(n_8219),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8622),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_8623),
.Y(n_9099)
);

INVx1_ASAP7_75t_SL g9100 ( 
.A(n_8629),
.Y(n_9100)
);

INVx2_ASAP7_75t_L g9101 ( 
.A(n_8670),
.Y(n_9101)
);

INVxp67_ASAP7_75t_L g9102 ( 
.A(n_8472),
.Y(n_9102)
);

INVx2_ASAP7_75t_L g9103 ( 
.A(n_8723),
.Y(n_9103)
);

INVxp67_ASAP7_75t_L g9104 ( 
.A(n_8505),
.Y(n_9104)
);

INVx1_ASAP7_75t_L g9105 ( 
.A(n_8236),
.Y(n_9105)
);

NAND2xp5_ASAP7_75t_SL g9106 ( 
.A(n_8624),
.B(n_5736),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8241),
.Y(n_9107)
);

NOR2xp33_ASAP7_75t_L g9108 ( 
.A(n_8299),
.B(n_5743),
.Y(n_9108)
);

OR2x6_ASAP7_75t_L g9109 ( 
.A(n_8397),
.B(n_5483),
.Y(n_9109)
);

BUFx6f_ASAP7_75t_L g9110 ( 
.A(n_8371),
.Y(n_9110)
);

AND2x2_ASAP7_75t_L g9111 ( 
.A(n_8509),
.B(n_6532),
.Y(n_9111)
);

BUFx6f_ASAP7_75t_L g9112 ( 
.A(n_8399),
.Y(n_9112)
);

BUFx6f_ASAP7_75t_L g9113 ( 
.A(n_8399),
.Y(n_9113)
);

INVx1_ASAP7_75t_L g9114 ( 
.A(n_8277),
.Y(n_9114)
);

NAND2xp5_ASAP7_75t_SL g9115 ( 
.A(n_8652),
.B(n_5745),
.Y(n_9115)
);

NAND3xp33_ASAP7_75t_L g9116 ( 
.A(n_8482),
.B(n_5749),
.C(n_5748),
.Y(n_9116)
);

INVx1_ASAP7_75t_L g9117 ( 
.A(n_8282),
.Y(n_9117)
);

INVx2_ASAP7_75t_SL g9118 ( 
.A(n_8415),
.Y(n_9118)
);

INVx1_ASAP7_75t_L g9119 ( 
.A(n_8308),
.Y(n_9119)
);

INVx2_ASAP7_75t_SL g9120 ( 
.A(n_8415),
.Y(n_9120)
);

INVx1_ASAP7_75t_L g9121 ( 
.A(n_8326),
.Y(n_9121)
);

OR2x6_ASAP7_75t_L g9122 ( 
.A(n_8668),
.B(n_5488),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_8727),
.Y(n_9123)
);

NAND2xp33_ASAP7_75t_L g9124 ( 
.A(n_8596),
.B(n_5753),
.Y(n_9124)
);

NAND2xp5_ASAP7_75t_L g9125 ( 
.A(n_8549),
.B(n_5756),
.Y(n_9125)
);

NOR2xp33_ASAP7_75t_L g9126 ( 
.A(n_8400),
.B(n_5759),
.Y(n_9126)
);

INVx2_ASAP7_75t_SL g9127 ( 
.A(n_8586),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_SL g9128 ( 
.A(n_8329),
.B(n_5760),
.Y(n_9128)
);

INVx1_ASAP7_75t_L g9129 ( 
.A(n_8335),
.Y(n_9129)
);

INVx1_ASAP7_75t_SL g9130 ( 
.A(n_8649),
.Y(n_9130)
);

NAND2xp33_ASAP7_75t_L g9131 ( 
.A(n_8596),
.B(n_5761),
.Y(n_9131)
);

INVx2_ASAP7_75t_L g9132 ( 
.A(n_8729),
.Y(n_9132)
);

INVx2_ASAP7_75t_L g9133 ( 
.A(n_8730),
.Y(n_9133)
);

NAND2xp5_ASAP7_75t_L g9134 ( 
.A(n_8511),
.B(n_5764),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8709),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_8381),
.Y(n_9136)
);

NOR2xp33_ASAP7_75t_L g9137 ( 
.A(n_8684),
.B(n_5768),
.Y(n_9137)
);

INVx2_ASAP7_75t_L g9138 ( 
.A(n_8645),
.Y(n_9138)
);

NAND2xp5_ASAP7_75t_SL g9139 ( 
.A(n_8367),
.B(n_5771),
.Y(n_9139)
);

INVx2_ASAP7_75t_L g9140 ( 
.A(n_8661),
.Y(n_9140)
);

BUFx3_ASAP7_75t_L g9141 ( 
.A(n_8249),
.Y(n_9141)
);

INVx1_ASAP7_75t_L g9142 ( 
.A(n_8401),
.Y(n_9142)
);

INVx2_ASAP7_75t_SL g9143 ( 
.A(n_8651),
.Y(n_9143)
);

BUFx2_ASAP7_75t_L g9144 ( 
.A(n_8341),
.Y(n_9144)
);

INVx2_ASAP7_75t_L g9145 ( 
.A(n_8667),
.Y(n_9145)
);

INVx1_ASAP7_75t_L g9146 ( 
.A(n_8425),
.Y(n_9146)
);

INVx2_ASAP7_75t_L g9147 ( 
.A(n_8675),
.Y(n_9147)
);

NAND2xp5_ASAP7_75t_SL g9148 ( 
.A(n_8392),
.B(n_8726),
.Y(n_9148)
);

BUFx10_ASAP7_75t_L g9149 ( 
.A(n_8440),
.Y(n_9149)
);

INVxp67_ASAP7_75t_L g9150 ( 
.A(n_8255),
.Y(n_9150)
);

OAI22xp5_ASAP7_75t_L g9151 ( 
.A1(n_8579),
.A2(n_8632),
.B1(n_8437),
.B2(n_8362),
.Y(n_9151)
);

INVx1_ASAP7_75t_SL g9152 ( 
.A(n_8413),
.Y(n_9152)
);

INVx2_ASAP7_75t_L g9153 ( 
.A(n_8694),
.Y(n_9153)
);

NAND3x1_ASAP7_75t_L g9154 ( 
.A(n_8715),
.B(n_5498),
.C(n_5496),
.Y(n_9154)
);

INVx2_ASAP7_75t_L g9155 ( 
.A(n_8695),
.Y(n_9155)
);

INVx2_ASAP7_75t_L g9156 ( 
.A(n_8703),
.Y(n_9156)
);

INVx2_ASAP7_75t_L g9157 ( 
.A(n_8708),
.Y(n_9157)
);

NAND2xp5_ASAP7_75t_SL g9158 ( 
.A(n_8488),
.B(n_5772),
.Y(n_9158)
);

NAND2xp5_ASAP7_75t_L g9159 ( 
.A(n_8533),
.B(n_8537),
.Y(n_9159)
);

INVx2_ASAP7_75t_L g9160 ( 
.A(n_8530),
.Y(n_9160)
);

AND2x2_ASAP7_75t_L g9161 ( 
.A(n_8289),
.B(n_6532),
.Y(n_9161)
);

AND2x2_ASAP7_75t_L g9162 ( 
.A(n_8441),
.B(n_5775),
.Y(n_9162)
);

INVx3_ASAP7_75t_L g9163 ( 
.A(n_8656),
.Y(n_9163)
);

INVx4_ASAP7_75t_L g9164 ( 
.A(n_8312),
.Y(n_9164)
);

INVx2_ASAP7_75t_L g9165 ( 
.A(n_8439),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_8480),
.Y(n_9166)
);

BUFx3_ASAP7_75t_L g9167 ( 
.A(n_8259),
.Y(n_9167)
);

NAND2xp5_ASAP7_75t_SL g9168 ( 
.A(n_8488),
.B(n_5776),
.Y(n_9168)
);

INVx1_ASAP7_75t_L g9169 ( 
.A(n_8450),
.Y(n_9169)
);

AND3x2_ASAP7_75t_L g9170 ( 
.A(n_8752),
.B(n_5500),
.C(n_5499),
.Y(n_9170)
);

AND2x2_ASAP7_75t_L g9171 ( 
.A(n_8470),
.B(n_8477),
.Y(n_9171)
);

INVx2_ASAP7_75t_L g9172 ( 
.A(n_8711),
.Y(n_9172)
);

NOR2x1p5_ASAP7_75t_L g9173 ( 
.A(n_8316),
.B(n_5779),
.Y(n_9173)
);

BUFx6f_ASAP7_75t_L g9174 ( 
.A(n_8233),
.Y(n_9174)
);

INVx2_ASAP7_75t_L g9175 ( 
.A(n_8713),
.Y(n_9175)
);

INVx3_ASAP7_75t_L g9176 ( 
.A(n_8656),
.Y(n_9176)
);

INVx2_ASAP7_75t_L g9177 ( 
.A(n_8714),
.Y(n_9177)
);

INVx2_ASAP7_75t_L g9178 ( 
.A(n_8720),
.Y(n_9178)
);

BUFx6f_ASAP7_75t_SL g9179 ( 
.A(n_8502),
.Y(n_9179)
);

INVx1_ASAP7_75t_L g9180 ( 
.A(n_8462),
.Y(n_9180)
);

BUFx3_ASAP7_75t_L g9181 ( 
.A(n_8260),
.Y(n_9181)
);

NAND2xp5_ASAP7_75t_SL g9182 ( 
.A(n_8506),
.B(n_5785),
.Y(n_9182)
);

NAND2xp5_ASAP7_75t_L g9183 ( 
.A(n_8473),
.B(n_5788),
.Y(n_9183)
);

NOR2xp33_ASAP7_75t_L g9184 ( 
.A(n_8679),
.B(n_5791),
.Y(n_9184)
);

NOR2x1p5_ASAP7_75t_L g9185 ( 
.A(n_8318),
.B(n_5796),
.Y(n_9185)
);

AO21x2_ASAP7_75t_L g9186 ( 
.A1(n_8747),
.A2(n_5506),
.B(n_5503),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_L g9187 ( 
.A(n_8743),
.B(n_5797),
.Y(n_9187)
);

INVx2_ASAP7_75t_L g9188 ( 
.A(n_8423),
.Y(n_9188)
);

INVx2_ASAP7_75t_L g9189 ( 
.A(n_8443),
.Y(n_9189)
);

INVx1_ASAP7_75t_L g9190 ( 
.A(n_8731),
.Y(n_9190)
);

INVx2_ASAP7_75t_L g9191 ( 
.A(n_8455),
.Y(n_9191)
);

INVx2_ASAP7_75t_L g9192 ( 
.A(n_8481),
.Y(n_9192)
);

INVx1_ASAP7_75t_L g9193 ( 
.A(n_8313),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_8660),
.Y(n_9194)
);

OAI22x1_ASAP7_75t_L g9195 ( 
.A1(n_8728),
.A2(n_8666),
.B1(n_8671),
.B2(n_8654),
.Y(n_9195)
);

BUFx10_ASAP7_75t_L g9196 ( 
.A(n_8257),
.Y(n_9196)
);

BUFx3_ASAP7_75t_L g9197 ( 
.A(n_8324),
.Y(n_9197)
);

AOI22xp33_ASAP7_75t_L g9198 ( 
.A1(n_8751),
.A2(n_6436),
.B1(n_6552),
.B2(n_6417),
.Y(n_9198)
);

HB1xp67_ASAP7_75t_L g9199 ( 
.A(n_8682),
.Y(n_9199)
);

AND2x2_ASAP7_75t_L g9200 ( 
.A(n_8559),
.B(n_5799),
.Y(n_9200)
);

CKINVDCx20_ASAP7_75t_R g9201 ( 
.A(n_8196),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8334),
.Y(n_9202)
);

INVx11_ASAP7_75t_L g9203 ( 
.A(n_8248),
.Y(n_9203)
);

INVx2_ASAP7_75t_L g9204 ( 
.A(n_8660),
.Y(n_9204)
);

INVx2_ASAP7_75t_L g9205 ( 
.A(n_8487),
.Y(n_9205)
);

NAND2xp5_ASAP7_75t_SL g9206 ( 
.A(n_8506),
.B(n_5800),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_8635),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_8327),
.Y(n_9208)
);

INVx1_ASAP7_75t_SL g9209 ( 
.A(n_8414),
.Y(n_9209)
);

INVx2_ASAP7_75t_L g9210 ( 
.A(n_8348),
.Y(n_9210)
);

INVx1_ASAP7_75t_SL g9211 ( 
.A(n_8435),
.Y(n_9211)
);

INVx4_ASAP7_75t_L g9212 ( 
.A(n_8330),
.Y(n_9212)
);

NAND2xp5_ASAP7_75t_SL g9213 ( 
.A(n_8332),
.B(n_8672),
.Y(n_9213)
);

INVx2_ASAP7_75t_L g9214 ( 
.A(n_8375),
.Y(n_9214)
);

INVx8_ASAP7_75t_L g9215 ( 
.A(n_8248),
.Y(n_9215)
);

INVx8_ASAP7_75t_L g9216 ( 
.A(n_8248),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_8701),
.Y(n_9217)
);

INVx2_ASAP7_75t_L g9218 ( 
.A(n_8386),
.Y(n_9218)
);

AO21x2_ASAP7_75t_L g9219 ( 
.A1(n_8750),
.A2(n_5513),
.B(n_5507),
.Y(n_9219)
);

INVx2_ASAP7_75t_L g9220 ( 
.A(n_8393),
.Y(n_9220)
);

NOR2xp33_ASAP7_75t_L g9221 ( 
.A(n_8543),
.B(n_5803),
.Y(n_9221)
);

INVx2_ASAP7_75t_L g9222 ( 
.A(n_8407),
.Y(n_9222)
);

BUFx3_ASAP7_75t_L g9223 ( 
.A(n_8524),
.Y(n_9223)
);

AND2x2_ASAP7_75t_L g9224 ( 
.A(n_8732),
.B(n_5805),
.Y(n_9224)
);

AND2x2_ASAP7_75t_L g9225 ( 
.A(n_8699),
.B(n_5806),
.Y(n_9225)
);

BUFx10_ASAP7_75t_L g9226 ( 
.A(n_8263),
.Y(n_9226)
);

INVx1_ASAP7_75t_L g9227 ( 
.A(n_8702),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_8546),
.Y(n_9228)
);

INVx2_ASAP7_75t_L g9229 ( 
.A(n_8609),
.Y(n_9229)
);

NOR2xp33_ASAP7_75t_L g9230 ( 
.A(n_8345),
.B(n_5810),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_8247),
.Y(n_9231)
);

INVx1_ASAP7_75t_L g9232 ( 
.A(n_8644),
.Y(n_9232)
);

INVx2_ASAP7_75t_SL g9233 ( 
.A(n_8604),
.Y(n_9233)
);

NAND2xp5_ASAP7_75t_SL g9234 ( 
.A(n_8677),
.B(n_5815),
.Y(n_9234)
);

AO21x2_ASAP7_75t_L g9235 ( 
.A1(n_8333),
.A2(n_8457),
.B(n_8396),
.Y(n_9235)
);

INVx4_ASAP7_75t_L g9236 ( 
.A(n_8685),
.Y(n_9236)
);

INVx2_ASAP7_75t_L g9237 ( 
.A(n_8234),
.Y(n_9237)
);

INVx2_ASAP7_75t_L g9238 ( 
.A(n_8239),
.Y(n_9238)
);

AND2x2_ASAP7_75t_L g9239 ( 
.A(n_8717),
.B(n_5817),
.Y(n_9239)
);

INVx2_ASAP7_75t_L g9240 ( 
.A(n_8279),
.Y(n_9240)
);

AND2x2_ASAP7_75t_L g9241 ( 
.A(n_8734),
.B(n_8736),
.Y(n_9241)
);

NAND2xp5_ASAP7_75t_L g9242 ( 
.A(n_8738),
.B(n_5818),
.Y(n_9242)
);

AND3x2_ASAP7_75t_L g9243 ( 
.A(n_8740),
.B(n_5519),
.C(n_5514),
.Y(n_9243)
);

AOI22xp33_ASAP7_75t_L g9244 ( 
.A1(n_8753),
.A2(n_6573),
.B1(n_6574),
.B2(n_6555),
.Y(n_9244)
);

HB1xp67_ASAP7_75t_L g9245 ( 
.A(n_8687),
.Y(n_9245)
);

NAND2xp5_ASAP7_75t_SL g9246 ( 
.A(n_8693),
.B(n_5821),
.Y(n_9246)
);

INVx2_ASAP7_75t_L g9247 ( 
.A(n_8676),
.Y(n_9247)
);

INVx2_ASAP7_75t_L g9248 ( 
.A(n_8233),
.Y(n_9248)
);

INVx2_ASAP7_75t_L g9249 ( 
.A(n_8261),
.Y(n_9249)
);

NAND2xp5_ASAP7_75t_SL g9250 ( 
.A(n_8697),
.B(n_5822),
.Y(n_9250)
);

INVx4_ASAP7_75t_L g9251 ( 
.A(n_8351),
.Y(n_9251)
);

INVxp67_ASAP7_75t_SL g9252 ( 
.A(n_8261),
.Y(n_9252)
);

INVx2_ASAP7_75t_L g9253 ( 
.A(n_8742),
.Y(n_9253)
);

AND2x2_ASAP7_75t_L g9254 ( 
.A(n_8554),
.B(n_5829),
.Y(n_9254)
);

AOI22xp33_ASAP7_75t_L g9255 ( 
.A1(n_8508),
.A2(n_6600),
.B1(n_6605),
.B2(n_6579),
.Y(n_9255)
);

BUFx10_ASAP7_75t_L g9256 ( 
.A(n_8264),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_8418),
.Y(n_9257)
);

INVx2_ASAP7_75t_L g9258 ( 
.A(n_8716),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_8737),
.Y(n_9259)
);

INVx1_ASAP7_75t_L g9260 ( 
.A(n_8705),
.Y(n_9260)
);

BUFx10_ASAP7_75t_L g9261 ( 
.A(n_8273),
.Y(n_9261)
);

NAND2xp5_ASAP7_75t_L g9262 ( 
.A(n_8700),
.B(n_5832),
.Y(n_9262)
);

INVx4_ASAP7_75t_L g9263 ( 
.A(n_8354),
.Y(n_9263)
);

AND2x2_ASAP7_75t_L g9264 ( 
.A(n_8356),
.B(n_5833),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_8683),
.Y(n_9265)
);

INVx1_ASAP7_75t_L g9266 ( 
.A(n_8611),
.Y(n_9266)
);

NOR2x1p5_ASAP7_75t_L g9267 ( 
.A(n_8719),
.B(n_5835),
.Y(n_9267)
);

NAND2xp5_ASAP7_75t_L g9268 ( 
.A(n_8513),
.B(n_5837),
.Y(n_9268)
);

INVx2_ASAP7_75t_L g9269 ( 
.A(n_8369),
.Y(n_9269)
);

INVx5_ASAP7_75t_L g9270 ( 
.A(n_8669),
.Y(n_9270)
);

CKINVDCx5p33_ASAP7_75t_R g9271 ( 
.A(n_8208),
.Y(n_9271)
);

INVx3_ASAP7_75t_L g9272 ( 
.A(n_8451),
.Y(n_9272)
);

INVx1_ASAP7_75t_L g9273 ( 
.A(n_8370),
.Y(n_9273)
);

INVx1_ASAP7_75t_L g9274 ( 
.A(n_8374),
.Y(n_9274)
);

NOR2xp33_ASAP7_75t_L g9275 ( 
.A(n_8395),
.B(n_5838),
.Y(n_9275)
);

INVx1_ASAP7_75t_L g9276 ( 
.A(n_8398),
.Y(n_9276)
);

NOR2xp33_ASAP7_75t_L g9277 ( 
.A(n_8665),
.B(n_5839),
.Y(n_9277)
);

NAND2xp5_ASAP7_75t_SL g9278 ( 
.A(n_8664),
.B(n_5841),
.Y(n_9278)
);

INVx2_ASAP7_75t_L g9279 ( 
.A(n_8595),
.Y(n_9279)
);

NAND2xp33_ASAP7_75t_SL g9280 ( 
.A(n_8706),
.B(n_5843),
.Y(n_9280)
);

NAND2xp5_ASAP7_75t_L g9281 ( 
.A(n_8486),
.B(n_5844),
.Y(n_9281)
);

INVx2_ASAP7_75t_SL g9282 ( 
.A(n_8547),
.Y(n_9282)
);

INVx1_ASAP7_75t_SL g9283 ( 
.A(n_8452),
.Y(n_9283)
);

INVx2_ASAP7_75t_L g9284 ( 
.A(n_8497),
.Y(n_9284)
);

AO22x2_ASAP7_75t_L g9285 ( 
.A1(n_8485),
.A2(n_5525),
.B1(n_5527),
.B2(n_5522),
.Y(n_9285)
);

BUFx6f_ASAP7_75t_L g9286 ( 
.A(n_8510),
.Y(n_9286)
);

INVx2_ASAP7_75t_L g9287 ( 
.A(n_8519),
.Y(n_9287)
);

INVx2_ASAP7_75t_L g9288 ( 
.A(n_8491),
.Y(n_9288)
);

INVx2_ASAP7_75t_L g9289 ( 
.A(n_8456),
.Y(n_9289)
);

NOR2x1p5_ASAP7_75t_L g9290 ( 
.A(n_8276),
.B(n_5845),
.Y(n_9290)
);

INVx2_ASAP7_75t_L g9291 ( 
.A(n_8468),
.Y(n_9291)
);

NAND2xp5_ASAP7_75t_L g9292 ( 
.A(n_8459),
.B(n_5846),
.Y(n_9292)
);

INVx1_ASAP7_75t_L g9293 ( 
.A(n_8585),
.Y(n_9293)
);

INVx4_ASAP7_75t_L g9294 ( 
.A(n_8284),
.Y(n_9294)
);

INVx3_ASAP7_75t_L g9295 ( 
.A(n_8250),
.Y(n_9295)
);

NAND2xp5_ASAP7_75t_L g9296 ( 
.A(n_8307),
.B(n_5848),
.Y(n_9296)
);

NOR2xp33_ASAP7_75t_L g9297 ( 
.A(n_8266),
.B(n_5854),
.Y(n_9297)
);

AND2x6_ASAP7_75t_L g9298 ( 
.A(n_8606),
.B(n_5533),
.Y(n_9298)
);

NAND2xp5_ASAP7_75t_L g9299 ( 
.A(n_8268),
.B(n_5857),
.Y(n_9299)
);

AND2x4_ASAP7_75t_L g9300 ( 
.A(n_8278),
.B(n_5535),
.Y(n_9300)
);

INVx4_ASAP7_75t_L g9301 ( 
.A(n_8286),
.Y(n_9301)
);

OR2x6_ASAP7_75t_L g9302 ( 
.A(n_8544),
.B(n_5536),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_8292),
.Y(n_9303)
);

NAND2xp5_ASAP7_75t_SL g9304 ( 
.A(n_8295),
.B(n_8296),
.Y(n_9304)
);

INVx2_ASAP7_75t_L g9305 ( 
.A(n_8302),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_8306),
.Y(n_9306)
);

NAND2xp5_ASAP7_75t_SL g9307 ( 
.A(n_8253),
.B(n_5860),
.Y(n_9307)
);

INVx2_ASAP7_75t_L g9308 ( 
.A(n_8285),
.Y(n_9308)
);

INVx1_ASAP7_75t_L g9309 ( 
.A(n_8725),
.Y(n_9309)
);

NOR2xp33_ASAP7_75t_L g9310 ( 
.A(n_8294),
.B(n_5861),
.Y(n_9310)
);

NAND2xp5_ASAP7_75t_SL g9311 ( 
.A(n_8698),
.B(n_5864),
.Y(n_9311)
);

BUFx6f_ASAP7_75t_L g9312 ( 
.A(n_8735),
.Y(n_9312)
);

AND2x6_ASAP7_75t_L g9313 ( 
.A(n_8896),
.B(n_5539),
.Y(n_9313)
);

BUFx2_ASAP7_75t_L g9314 ( 
.A(n_8774),
.Y(n_9314)
);

NOR2xp33_ASAP7_75t_L g9315 ( 
.A(n_8822),
.B(n_8756),
.Y(n_9315)
);

OAI22xp33_ASAP7_75t_L g9316 ( 
.A1(n_8844),
.A2(n_8770),
.B1(n_8775),
.B2(n_9045),
.Y(n_9316)
);

INVx1_ASAP7_75t_L g9317 ( 
.A(n_8767),
.Y(n_9317)
);

INVx3_ASAP7_75t_L g9318 ( 
.A(n_8795),
.Y(n_9318)
);

BUFx2_ASAP7_75t_L g9319 ( 
.A(n_8830),
.Y(n_9319)
);

AOI22xp33_ASAP7_75t_L g9320 ( 
.A1(n_8781),
.A2(n_6617),
.B1(n_5563),
.B2(n_5567),
.Y(n_9320)
);

AND2x4_ASAP7_75t_L g9321 ( 
.A(n_8811),
.B(n_8555),
.Y(n_9321)
);

NAND2xp5_ASAP7_75t_L g9322 ( 
.A(n_8758),
.B(n_5865),
.Y(n_9322)
);

BUFx6f_ASAP7_75t_L g9323 ( 
.A(n_8784),
.Y(n_9323)
);

INVx3_ASAP7_75t_L g9324 ( 
.A(n_9197),
.Y(n_9324)
);

INVx1_ASAP7_75t_L g9325 ( 
.A(n_8772),
.Y(n_9325)
);

INVx2_ASAP7_75t_L g9326 ( 
.A(n_9103),
.Y(n_9326)
);

INVx3_ASAP7_75t_L g9327 ( 
.A(n_9174),
.Y(n_9327)
);

AND2x6_ASAP7_75t_L g9328 ( 
.A(n_9105),
.B(n_5548),
.Y(n_9328)
);

INVxp67_ASAP7_75t_L g9329 ( 
.A(n_8899),
.Y(n_9329)
);

AND2x6_ASAP7_75t_L g9330 ( 
.A(n_9107),
.B(n_5571),
.Y(n_9330)
);

NAND2x1p5_ASAP7_75t_L g9331 ( 
.A(n_8793),
.B(n_8881),
.Y(n_9331)
);

BUFx2_ASAP7_75t_L g9332 ( 
.A(n_8764),
.Y(n_9332)
);

OR2x2_ASAP7_75t_L g9333 ( 
.A(n_8776),
.B(n_8748),
.Y(n_9333)
);

INVx1_ASAP7_75t_L g9334 ( 
.A(n_8773),
.Y(n_9334)
);

BUFx2_ASAP7_75t_SL g9335 ( 
.A(n_8888),
.Y(n_9335)
);

AND2x2_ASAP7_75t_L g9336 ( 
.A(n_8789),
.B(n_5868),
.Y(n_9336)
);

BUFx3_ASAP7_75t_L g9337 ( 
.A(n_8792),
.Y(n_9337)
);

AND2x6_ASAP7_75t_L g9338 ( 
.A(n_9114),
.B(n_5572),
.Y(n_9338)
);

OAI22xp33_ASAP7_75t_L g9339 ( 
.A1(n_9159),
.A2(n_5870),
.B1(n_5871),
.B2(n_5869),
.Y(n_9339)
);

OR2x2_ASAP7_75t_L g9340 ( 
.A(n_9152),
.B(n_5872),
.Y(n_9340)
);

NAND2xp5_ASAP7_75t_SL g9341 ( 
.A(n_8923),
.B(n_5876),
.Y(n_9341)
);

INVx4_ASAP7_75t_L g9342 ( 
.A(n_8792),
.Y(n_9342)
);

NOR2xp33_ASAP7_75t_L g9343 ( 
.A(n_9126),
.B(n_9117),
.Y(n_9343)
);

INVx2_ASAP7_75t_L g9344 ( 
.A(n_9123),
.Y(n_9344)
);

BUFx4f_ASAP7_75t_L g9345 ( 
.A(n_9286),
.Y(n_9345)
);

NOR2xp33_ASAP7_75t_SL g9346 ( 
.A(n_8861),
.B(n_8712),
.Y(n_9346)
);

AND2x6_ASAP7_75t_L g9347 ( 
.A(n_9119),
.B(n_5574),
.Y(n_9347)
);

NOR2xp33_ASAP7_75t_L g9348 ( 
.A(n_9121),
.B(n_5877),
.Y(n_9348)
);

NAND2xp5_ASAP7_75t_L g9349 ( 
.A(n_9129),
.B(n_5878),
.Y(n_9349)
);

AOI22xp33_ASAP7_75t_L g9350 ( 
.A1(n_9298),
.A2(n_5576),
.B1(n_5583),
.B2(n_5575),
.Y(n_9350)
);

INVx1_ASAP7_75t_L g9351 ( 
.A(n_8780),
.Y(n_9351)
);

INVx2_ASAP7_75t_L g9352 ( 
.A(n_9132),
.Y(n_9352)
);

INVx1_ASAP7_75t_L g9353 ( 
.A(n_8783),
.Y(n_9353)
);

NAND2xp5_ASAP7_75t_SL g9354 ( 
.A(n_9136),
.B(n_5880),
.Y(n_9354)
);

NOR2xp33_ASAP7_75t_L g9355 ( 
.A(n_9142),
.B(n_5884),
.Y(n_9355)
);

INVx1_ASAP7_75t_L g9356 ( 
.A(n_8785),
.Y(n_9356)
);

INVx1_ASAP7_75t_L g9357 ( 
.A(n_8791),
.Y(n_9357)
);

CKINVDCx5p33_ASAP7_75t_R g9358 ( 
.A(n_8794),
.Y(n_9358)
);

NAND2xp5_ASAP7_75t_L g9359 ( 
.A(n_9146),
.B(n_5887),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_9169),
.B(n_5892),
.Y(n_9360)
);

INVx2_ASAP7_75t_L g9361 ( 
.A(n_9133),
.Y(n_9361)
);

BUFx3_ASAP7_75t_L g9362 ( 
.A(n_9174),
.Y(n_9362)
);

NOR2xp33_ASAP7_75t_L g9363 ( 
.A(n_9180),
.B(n_5893),
.Y(n_9363)
);

NAND2xp5_ASAP7_75t_L g9364 ( 
.A(n_8921),
.B(n_5899),
.Y(n_9364)
);

BUFx4f_ASAP7_75t_L g9365 ( 
.A(n_9286),
.Y(n_9365)
);

BUFx10_ASAP7_75t_L g9366 ( 
.A(n_9230),
.Y(n_9366)
);

BUFx6f_ASAP7_75t_L g9367 ( 
.A(n_8784),
.Y(n_9367)
);

CKINVDCx5p33_ASAP7_75t_R g9368 ( 
.A(n_8891),
.Y(n_9368)
);

OR2x2_ASAP7_75t_L g9369 ( 
.A(n_9209),
.B(n_5900),
.Y(n_9369)
);

INVx3_ASAP7_75t_L g9370 ( 
.A(n_8827),
.Y(n_9370)
);

NAND2xp5_ASAP7_75t_SL g9371 ( 
.A(n_9083),
.B(n_5902),
.Y(n_9371)
);

AND2x4_ASAP7_75t_L g9372 ( 
.A(n_9236),
.B(n_8733),
.Y(n_9372)
);

INVx1_ASAP7_75t_L g9373 ( 
.A(n_8799),
.Y(n_9373)
);

AND2x2_ASAP7_75t_L g9374 ( 
.A(n_8986),
.B(n_5903),
.Y(n_9374)
);

NAND2xp5_ASAP7_75t_L g9375 ( 
.A(n_8821),
.B(n_5904),
.Y(n_9375)
);

BUFx4f_ASAP7_75t_L g9376 ( 
.A(n_8797),
.Y(n_9376)
);

BUFx4f_ASAP7_75t_L g9377 ( 
.A(n_8797),
.Y(n_9377)
);

AND2x2_ASAP7_75t_L g9378 ( 
.A(n_9035),
.B(n_5905),
.Y(n_9378)
);

INVx3_ASAP7_75t_L g9379 ( 
.A(n_8857),
.Y(n_9379)
);

NOR2xp33_ASAP7_75t_L g9380 ( 
.A(n_9150),
.B(n_5906),
.Y(n_9380)
);

INVx1_ASAP7_75t_L g9381 ( 
.A(n_8800),
.Y(n_9381)
);

OAI21xp5_ASAP7_75t_L g9382 ( 
.A1(n_9092),
.A2(n_5587),
.B(n_5586),
.Y(n_9382)
);

AND2x2_ASAP7_75t_L g9383 ( 
.A(n_9200),
.B(n_5908),
.Y(n_9383)
);

AND2x4_ASAP7_75t_SL g9384 ( 
.A(n_9164),
.B(n_8741),
.Y(n_9384)
);

INVx4_ASAP7_75t_L g9385 ( 
.A(n_8852),
.Y(n_9385)
);

INVx1_ASAP7_75t_L g9386 ( 
.A(n_8809),
.Y(n_9386)
);

AND2x6_ASAP7_75t_L g9387 ( 
.A(n_9171),
.B(n_5594),
.Y(n_9387)
);

NAND2xp5_ASAP7_75t_L g9388 ( 
.A(n_8831),
.B(n_8934),
.Y(n_9388)
);

INVx2_ASAP7_75t_L g9389 ( 
.A(n_8771),
.Y(n_9389)
);

AND2x4_ASAP7_75t_L g9390 ( 
.A(n_9060),
.B(n_8963),
.Y(n_9390)
);

INVx2_ASAP7_75t_L g9391 ( 
.A(n_8778),
.Y(n_9391)
);

NOR2xp33_ASAP7_75t_L g9392 ( 
.A(n_9008),
.B(n_5909),
.Y(n_9392)
);

CKINVDCx5p33_ASAP7_75t_R g9393 ( 
.A(n_9006),
.Y(n_9393)
);

HB1xp67_ASAP7_75t_L g9394 ( 
.A(n_8838),
.Y(n_9394)
);

INVx1_ASAP7_75t_L g9395 ( 
.A(n_8833),
.Y(n_9395)
);

INVx3_ASAP7_75t_L g9396 ( 
.A(n_9212),
.Y(n_9396)
);

BUFx6f_ASAP7_75t_L g9397 ( 
.A(n_8852),
.Y(n_9397)
);

INVx4_ASAP7_75t_L g9398 ( 
.A(n_8894),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_L g9399 ( 
.A(n_8935),
.B(n_8937),
.Y(n_9399)
);

INVx5_ASAP7_75t_L g9400 ( 
.A(n_8894),
.Y(n_9400)
);

BUFx3_ASAP7_75t_L g9401 ( 
.A(n_8907),
.Y(n_9401)
);

CKINVDCx20_ASAP7_75t_R g9402 ( 
.A(n_9201),
.Y(n_9402)
);

NOR2xp33_ASAP7_75t_L g9403 ( 
.A(n_8782),
.B(n_5910),
.Y(n_9403)
);

INVx1_ASAP7_75t_L g9404 ( 
.A(n_8847),
.Y(n_9404)
);

AND2x2_ASAP7_75t_L g9405 ( 
.A(n_9111),
.B(n_5912),
.Y(n_9405)
);

AND2x6_ASAP7_75t_L g9406 ( 
.A(n_9258),
.B(n_5595),
.Y(n_9406)
);

NAND2xp33_ASAP7_75t_L g9407 ( 
.A(n_9215),
.B(n_5916),
.Y(n_9407)
);

NOR2xp33_ASAP7_75t_L g9408 ( 
.A(n_8777),
.B(n_5917),
.Y(n_9408)
);

BUFx2_ASAP7_75t_L g9409 ( 
.A(n_8841),
.Y(n_9409)
);

INVx1_ASAP7_75t_L g9410 ( 
.A(n_8858),
.Y(n_9410)
);

AND2x4_ASAP7_75t_L g9411 ( 
.A(n_9127),
.B(n_5603),
.Y(n_9411)
);

BUFx3_ASAP7_75t_L g9412 ( 
.A(n_8907),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8860),
.Y(n_9413)
);

OAI22xp33_ASAP7_75t_L g9414 ( 
.A1(n_9037),
.A2(n_5919),
.B1(n_5922),
.B2(n_5918),
.Y(n_9414)
);

AND2x4_ASAP7_75t_L g9415 ( 
.A(n_9003),
.B(n_5604),
.Y(n_9415)
);

CKINVDCx16_ASAP7_75t_R g9416 ( 
.A(n_8990),
.Y(n_9416)
);

AOI22xp5_ASAP7_75t_L g9417 ( 
.A1(n_8763),
.A2(n_5925),
.B1(n_5926),
.B2(n_5923),
.Y(n_9417)
);

BUFx3_ASAP7_75t_L g9418 ( 
.A(n_8979),
.Y(n_9418)
);

INVx2_ASAP7_75t_L g9419 ( 
.A(n_8790),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_8865),
.Y(n_9420)
);

AND3x4_ASAP7_75t_L g9421 ( 
.A(n_9279),
.B(n_5928),
.C(n_5927),
.Y(n_9421)
);

OR2x2_ASAP7_75t_L g9422 ( 
.A(n_9211),
.B(n_5929),
.Y(n_9422)
);

AND2x2_ASAP7_75t_L g9423 ( 
.A(n_9162),
.B(n_5933),
.Y(n_9423)
);

OR2x2_ASAP7_75t_SL g9424 ( 
.A(n_8848),
.B(n_5605),
.Y(n_9424)
);

INVx8_ASAP7_75t_L g9425 ( 
.A(n_8979),
.Y(n_9425)
);

INVx4_ASAP7_75t_L g9426 ( 
.A(n_9005),
.Y(n_9426)
);

NAND2xp5_ASAP7_75t_SL g9427 ( 
.A(n_8980),
.B(n_5939),
.Y(n_9427)
);

AND2x6_ASAP7_75t_L g9428 ( 
.A(n_9293),
.B(n_5617),
.Y(n_9428)
);

AND2x6_ASAP7_75t_L g9429 ( 
.A(n_9005),
.B(n_5621),
.Y(n_9429)
);

BUFx3_ASAP7_75t_L g9430 ( 
.A(n_9066),
.Y(n_9430)
);

NAND2xp5_ASAP7_75t_SL g9431 ( 
.A(n_9102),
.B(n_5944),
.Y(n_9431)
);

INVxp33_ASAP7_75t_SL g9432 ( 
.A(n_9271),
.Y(n_9432)
);

AOI22xp33_ASAP7_75t_L g9433 ( 
.A1(n_9298),
.A2(n_5631),
.B1(n_5636),
.B2(n_5623),
.Y(n_9433)
);

INVx2_ASAP7_75t_L g9434 ( 
.A(n_8798),
.Y(n_9434)
);

AND2x6_ASAP7_75t_L g9435 ( 
.A(n_9066),
.B(n_5639),
.Y(n_9435)
);

INVx2_ASAP7_75t_L g9436 ( 
.A(n_8801),
.Y(n_9436)
);

NOR2xp33_ASAP7_75t_L g9437 ( 
.A(n_8804),
.B(n_5947),
.Y(n_9437)
);

CKINVDCx5p33_ASAP7_75t_R g9438 ( 
.A(n_8925),
.Y(n_9438)
);

NOR2xp33_ASAP7_75t_L g9439 ( 
.A(n_8787),
.B(n_5955),
.Y(n_9439)
);

INVx2_ASAP7_75t_L g9440 ( 
.A(n_8802),
.Y(n_9440)
);

INVx2_ASAP7_75t_L g9441 ( 
.A(n_8803),
.Y(n_9441)
);

INVx4_ASAP7_75t_L g9442 ( 
.A(n_9110),
.Y(n_9442)
);

INVx1_ASAP7_75t_L g9443 ( 
.A(n_8867),
.Y(n_9443)
);

AND2x6_ASAP7_75t_L g9444 ( 
.A(n_9110),
.B(n_5644),
.Y(n_9444)
);

INVx3_ASAP7_75t_L g9445 ( 
.A(n_9112),
.Y(n_9445)
);

NAND2xp5_ASAP7_75t_SL g9446 ( 
.A(n_8922),
.B(n_5956),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_8869),
.Y(n_9447)
);

NAND2xp5_ASAP7_75t_SL g9448 ( 
.A(n_8948),
.B(n_5957),
.Y(n_9448)
);

CKINVDCx5p33_ASAP7_75t_R g9449 ( 
.A(n_8952),
.Y(n_9449)
);

NOR2xp33_ASAP7_75t_L g9450 ( 
.A(n_8903),
.B(n_5959),
.Y(n_9450)
);

INVx1_ASAP7_75t_L g9451 ( 
.A(n_8870),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_8885),
.Y(n_9452)
);

INVxp67_ASAP7_75t_SL g9453 ( 
.A(n_9081),
.Y(n_9453)
);

AND2x6_ASAP7_75t_L g9454 ( 
.A(n_9112),
.B(n_5647),
.Y(n_9454)
);

CKINVDCx5p33_ASAP7_75t_R g9455 ( 
.A(n_8962),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_8886),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_8887),
.Y(n_9457)
);

NAND2xp5_ASAP7_75t_L g9458 ( 
.A(n_8912),
.B(n_5960),
.Y(n_9458)
);

AOI22xp5_ASAP7_75t_L g9459 ( 
.A1(n_9014),
.A2(n_5962),
.B1(n_5964),
.B2(n_5961),
.Y(n_9459)
);

BUFx3_ASAP7_75t_L g9460 ( 
.A(n_9113),
.Y(n_9460)
);

NAND2xp5_ASAP7_75t_SL g9461 ( 
.A(n_9104),
.B(n_5968),
.Y(n_9461)
);

INVx2_ASAP7_75t_L g9462 ( 
.A(n_8806),
.Y(n_9462)
);

INVx4_ASAP7_75t_SL g9463 ( 
.A(n_9179),
.Y(n_9463)
);

INVx4_ASAP7_75t_L g9464 ( 
.A(n_9113),
.Y(n_9464)
);

AND2x6_ASAP7_75t_L g9465 ( 
.A(n_9273),
.B(n_5655),
.Y(n_9465)
);

BUFx3_ASAP7_75t_L g9466 ( 
.A(n_8992),
.Y(n_9466)
);

INVx2_ASAP7_75t_L g9467 ( 
.A(n_8814),
.Y(n_9467)
);

CKINVDCx20_ASAP7_75t_R g9468 ( 
.A(n_8911),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_SL g9469 ( 
.A(n_8817),
.B(n_5969),
.Y(n_9469)
);

INVx5_ASAP7_75t_L g9470 ( 
.A(n_8982),
.Y(n_9470)
);

INVx2_ASAP7_75t_SL g9471 ( 
.A(n_9248),
.Y(n_9471)
);

BUFx3_ASAP7_75t_L g9472 ( 
.A(n_8998),
.Y(n_9472)
);

AOI22xp33_ASAP7_75t_L g9473 ( 
.A1(n_9298),
.A2(n_5658),
.B1(n_5662),
.B2(n_5656),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_SL g9474 ( 
.A(n_8818),
.B(n_5972),
.Y(n_9474)
);

INVx4_ASAP7_75t_SL g9475 ( 
.A(n_9312),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_8823),
.Y(n_9476)
);

AND2x2_ASAP7_75t_SL g9477 ( 
.A(n_9144),
.B(n_5668),
.Y(n_9477)
);

AOI21x1_ASAP7_75t_L g9478 ( 
.A1(n_9253),
.A2(n_5675),
.B(n_5669),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_8889),
.Y(n_9479)
);

INVx1_ASAP7_75t_SL g9480 ( 
.A(n_9283),
.Y(n_9480)
);

AOI22xp5_ASAP7_75t_L g9481 ( 
.A1(n_9184),
.A2(n_5974),
.B1(n_5975),
.B2(n_5973),
.Y(n_9481)
);

AOI22xp33_ASAP7_75t_L g9482 ( 
.A1(n_8766),
.A2(n_8825),
.B1(n_8828),
.B2(n_8824),
.Y(n_9482)
);

BUFx6f_ASAP7_75t_L g9483 ( 
.A(n_9046),
.Y(n_9483)
);

NOR2xp33_ASAP7_75t_L g9484 ( 
.A(n_9296),
.B(n_5976),
.Y(n_9484)
);

INVx2_ASAP7_75t_L g9485 ( 
.A(n_8829),
.Y(n_9485)
);

INVx1_ASAP7_75t_L g9486 ( 
.A(n_8890),
.Y(n_9486)
);

NOR2xp33_ASAP7_75t_L g9487 ( 
.A(n_9275),
.B(n_5977),
.Y(n_9487)
);

INVxp67_ASAP7_75t_SL g9488 ( 
.A(n_8898),
.Y(n_9488)
);

BUFx3_ASAP7_75t_L g9489 ( 
.A(n_9097),
.Y(n_9489)
);

INVx1_ASAP7_75t_L g9490 ( 
.A(n_8897),
.Y(n_9490)
);

AND2x2_ASAP7_75t_L g9491 ( 
.A(n_9254),
.B(n_9161),
.Y(n_9491)
);

INVx5_ASAP7_75t_L g9492 ( 
.A(n_9015),
.Y(n_9492)
);

INVx2_ASAP7_75t_L g9493 ( 
.A(n_8832),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_8906),
.Y(n_9494)
);

INVx1_ASAP7_75t_L g9495 ( 
.A(n_8909),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_8916),
.Y(n_9496)
);

INVx4_ASAP7_75t_L g9497 ( 
.A(n_9270),
.Y(n_9497)
);

NOR2xp33_ASAP7_75t_L g9498 ( 
.A(n_9299),
.B(n_5983),
.Y(n_9498)
);

INVx2_ASAP7_75t_L g9499 ( 
.A(n_8837),
.Y(n_9499)
);

NOR2xp33_ASAP7_75t_L g9500 ( 
.A(n_8965),
.B(n_9079),
.Y(n_9500)
);

OR2x6_ASAP7_75t_L g9501 ( 
.A(n_9215),
.B(n_5677),
.Y(n_9501)
);

INVx1_ASAP7_75t_L g9502 ( 
.A(n_8932),
.Y(n_9502)
);

INVx3_ASAP7_75t_L g9503 ( 
.A(n_9053),
.Y(n_9503)
);

INVx2_ASAP7_75t_L g9504 ( 
.A(n_8839),
.Y(n_9504)
);

INVx1_ASAP7_75t_L g9505 ( 
.A(n_8940),
.Y(n_9505)
);

BUFx6f_ASAP7_75t_L g9506 ( 
.A(n_9041),
.Y(n_9506)
);

NOR2xp33_ASAP7_75t_L g9507 ( 
.A(n_9086),
.B(n_5984),
.Y(n_9507)
);

INVx2_ASAP7_75t_L g9508 ( 
.A(n_8840),
.Y(n_9508)
);

INVx2_ASAP7_75t_L g9509 ( 
.A(n_8843),
.Y(n_9509)
);

NOR2xp33_ASAP7_75t_L g9510 ( 
.A(n_9125),
.B(n_5986),
.Y(n_9510)
);

NAND2xp5_ASAP7_75t_SL g9511 ( 
.A(n_8845),
.B(n_5987),
.Y(n_9511)
);

AND2x4_ASAP7_75t_L g9512 ( 
.A(n_9205),
.B(n_5679),
.Y(n_9512)
);

INVx1_ASAP7_75t_L g9513 ( 
.A(n_8849),
.Y(n_9513)
);

BUFx4f_ASAP7_75t_L g9514 ( 
.A(n_9312),
.Y(n_9514)
);

NAND2xp5_ASAP7_75t_SL g9515 ( 
.A(n_8850),
.B(n_5988),
.Y(n_9515)
);

INVx3_ASAP7_75t_L g9516 ( 
.A(n_8812),
.Y(n_9516)
);

INVx2_ASAP7_75t_L g9517 ( 
.A(n_8853),
.Y(n_9517)
);

INVx1_ASAP7_75t_L g9518 ( 
.A(n_8854),
.Y(n_9518)
);

INVx2_ASAP7_75t_L g9519 ( 
.A(n_8855),
.Y(n_9519)
);

NOR2xp33_ASAP7_75t_L g9520 ( 
.A(n_8915),
.B(n_5989),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8862),
.Y(n_9521)
);

INVx5_ASAP7_75t_L g9522 ( 
.A(n_9196),
.Y(n_9522)
);

NOR2xp33_ASAP7_75t_L g9523 ( 
.A(n_8893),
.B(n_5990),
.Y(n_9523)
);

AND2x4_ASAP7_75t_L g9524 ( 
.A(n_9233),
.B(n_5684),
.Y(n_9524)
);

AND2x6_ASAP7_75t_L g9525 ( 
.A(n_9274),
.B(n_5689),
.Y(n_9525)
);

INVx3_ASAP7_75t_L g9526 ( 
.A(n_8819),
.Y(n_9526)
);

INVx1_ASAP7_75t_L g9527 ( 
.A(n_8866),
.Y(n_9527)
);

NAND2xp5_ASAP7_75t_L g9528 ( 
.A(n_9002),
.B(n_5991),
.Y(n_9528)
);

AND2x4_ASAP7_75t_L g9529 ( 
.A(n_9241),
.B(n_5691),
.Y(n_9529)
);

INVx1_ASAP7_75t_L g9530 ( 
.A(n_8871),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_8873),
.Y(n_9531)
);

INVx3_ASAP7_75t_L g9532 ( 
.A(n_8846),
.Y(n_9532)
);

AND2x4_ASAP7_75t_L g9533 ( 
.A(n_8868),
.B(n_5695),
.Y(n_9533)
);

NOR2xp33_ASAP7_75t_L g9534 ( 
.A(n_8920),
.B(n_5993),
.Y(n_9534)
);

AND2x2_ASAP7_75t_L g9535 ( 
.A(n_9264),
.B(n_5994),
.Y(n_9535)
);

NAND2xp5_ASAP7_75t_SL g9536 ( 
.A(n_8876),
.B(n_5996),
.Y(n_9536)
);

AND2x6_ASAP7_75t_L g9537 ( 
.A(n_9276),
.B(n_5698),
.Y(n_9537)
);

INVx4_ASAP7_75t_SL g9538 ( 
.A(n_9109),
.Y(n_9538)
);

INVx2_ASAP7_75t_SL g9539 ( 
.A(n_9249),
.Y(n_9539)
);

AND2x6_ASAP7_75t_L g9540 ( 
.A(n_9309),
.B(n_5704),
.Y(n_9540)
);

AND2x6_ASAP7_75t_L g9541 ( 
.A(n_9269),
.B(n_5706),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_8877),
.Y(n_9542)
);

NAND2xp5_ASAP7_75t_SL g9543 ( 
.A(n_8883),
.B(n_6001),
.Y(n_9543)
);

OAI22xp33_ASAP7_75t_L g9544 ( 
.A1(n_9057),
.A2(n_6009),
.B1(n_6010),
.B2(n_6003),
.Y(n_9544)
);

INVx1_ASAP7_75t_L g9545 ( 
.A(n_8895),
.Y(n_9545)
);

INVx3_ASAP7_75t_L g9546 ( 
.A(n_8879),
.Y(n_9546)
);

INVx2_ASAP7_75t_SL g9547 ( 
.A(n_9143),
.Y(n_9547)
);

INVx1_ASAP7_75t_L g9548 ( 
.A(n_8902),
.Y(n_9548)
);

BUFx3_ASAP7_75t_L g9549 ( 
.A(n_9141),
.Y(n_9549)
);

NAND2xp5_ASAP7_75t_SL g9550 ( 
.A(n_8905),
.B(n_6011),
.Y(n_9550)
);

NAND2xp5_ASAP7_75t_SL g9551 ( 
.A(n_8938),
.B(n_8939),
.Y(n_9551)
);

NAND2xp5_ASAP7_75t_SL g9552 ( 
.A(n_8786),
.B(n_6012),
.Y(n_9552)
);

INVx1_ASAP7_75t_L g9553 ( 
.A(n_9010),
.Y(n_9553)
);

BUFx6f_ASAP7_75t_L g9554 ( 
.A(n_9118),
.Y(n_9554)
);

INVxp67_ASAP7_75t_L g9555 ( 
.A(n_9245),
.Y(n_9555)
);

INVx2_ASAP7_75t_L g9556 ( 
.A(n_9101),
.Y(n_9556)
);

BUFx6f_ASAP7_75t_SL g9557 ( 
.A(n_9226),
.Y(n_9557)
);

AND2x6_ASAP7_75t_L g9558 ( 
.A(n_9193),
.B(n_5717),
.Y(n_9558)
);

BUFx2_ASAP7_75t_L g9559 ( 
.A(n_9289),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_9018),
.Y(n_9560)
);

BUFx8_ASAP7_75t_SL g9561 ( 
.A(n_9091),
.Y(n_9561)
);

INVx4_ASAP7_75t_L g9562 ( 
.A(n_9270),
.Y(n_9562)
);

INVx1_ASAP7_75t_L g9563 ( 
.A(n_9023),
.Y(n_9563)
);

INVx2_ASAP7_75t_L g9564 ( 
.A(n_9135),
.Y(n_9564)
);

NOR2xp33_ASAP7_75t_L g9565 ( 
.A(n_8943),
.B(n_6013),
.Y(n_9565)
);

NAND2xp5_ASAP7_75t_L g9566 ( 
.A(n_9034),
.B(n_6014),
.Y(n_9566)
);

NAND2xp5_ASAP7_75t_L g9567 ( 
.A(n_8953),
.B(n_6015),
.Y(n_9567)
);

INVx1_ASAP7_75t_SL g9568 ( 
.A(n_9100),
.Y(n_9568)
);

AND2x6_ASAP7_75t_L g9569 ( 
.A(n_9202),
.B(n_9207),
.Y(n_9569)
);

INVx3_ASAP7_75t_L g9570 ( 
.A(n_8929),
.Y(n_9570)
);

AND2x2_ASAP7_75t_L g9571 ( 
.A(n_8931),
.B(n_6016),
.Y(n_9571)
);

INVx4_ASAP7_75t_L g9572 ( 
.A(n_8958),
.Y(n_9572)
);

BUFx10_ASAP7_75t_L g9573 ( 
.A(n_9277),
.Y(n_9573)
);

NAND2xp5_ASAP7_75t_L g9574 ( 
.A(n_8961),
.B(n_6020),
.Y(n_9574)
);

INVx1_ASAP7_75t_L g9575 ( 
.A(n_9026),
.Y(n_9575)
);

AND2x2_ASAP7_75t_SL g9576 ( 
.A(n_9251),
.B(n_5719),
.Y(n_9576)
);

NAND2xp5_ASAP7_75t_SL g9577 ( 
.A(n_8856),
.B(n_6022),
.Y(n_9577)
);

INVx2_ASAP7_75t_SL g9578 ( 
.A(n_9194),
.Y(n_9578)
);

INVx4_ASAP7_75t_L g9579 ( 
.A(n_8969),
.Y(n_9579)
);

NOR2xp33_ASAP7_75t_L g9580 ( 
.A(n_8971),
.B(n_6023),
.Y(n_9580)
);

INVx3_ASAP7_75t_L g9581 ( 
.A(n_8988),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_9032),
.Y(n_9582)
);

INVx1_ASAP7_75t_L g9583 ( 
.A(n_9033),
.Y(n_9583)
);

INVx1_ASAP7_75t_L g9584 ( 
.A(n_9039),
.Y(n_9584)
);

INVx1_ASAP7_75t_L g9585 ( 
.A(n_9047),
.Y(n_9585)
);

INVx3_ASAP7_75t_L g9586 ( 
.A(n_9009),
.Y(n_9586)
);

AOI22xp5_ASAP7_75t_L g9587 ( 
.A1(n_9221),
.A2(n_6027),
.B1(n_6029),
.B2(n_6024),
.Y(n_9587)
);

AND2x6_ASAP7_75t_L g9588 ( 
.A(n_9217),
.B(n_5721),
.Y(n_9588)
);

INVx1_ASAP7_75t_L g9589 ( 
.A(n_9052),
.Y(n_9589)
);

NAND2xp5_ASAP7_75t_L g9590 ( 
.A(n_9001),
.B(n_6030),
.Y(n_9590)
);

INVx2_ASAP7_75t_L g9591 ( 
.A(n_8759),
.Y(n_9591)
);

NOR2xp33_ASAP7_75t_L g9592 ( 
.A(n_9108),
.B(n_6033),
.Y(n_9592)
);

INVx4_ASAP7_75t_L g9593 ( 
.A(n_9024),
.Y(n_9593)
);

INVx1_ASAP7_75t_L g9594 ( 
.A(n_9061),
.Y(n_9594)
);

BUFx3_ASAP7_75t_L g9595 ( 
.A(n_9167),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_9065),
.Y(n_9596)
);

NAND2xp33_ASAP7_75t_L g9597 ( 
.A(n_9216),
.B(n_6040),
.Y(n_9597)
);

INVx1_ASAP7_75t_L g9598 ( 
.A(n_9067),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_8760),
.Y(n_9599)
);

INVx1_ASAP7_75t_L g9600 ( 
.A(n_9070),
.Y(n_9600)
);

INVx2_ASAP7_75t_L g9601 ( 
.A(n_8761),
.Y(n_9601)
);

NAND2xp5_ASAP7_75t_SL g9602 ( 
.A(n_8875),
.B(n_8805),
.Y(n_9602)
);

NOR2x1p5_ASAP7_75t_L g9603 ( 
.A(n_8930),
.B(n_6043),
.Y(n_9603)
);

AND2x4_ASAP7_75t_L g9604 ( 
.A(n_9058),
.B(n_5730),
.Y(n_9604)
);

INVx2_ASAP7_75t_SL g9605 ( 
.A(n_9204),
.Y(n_9605)
);

INVx2_ASAP7_75t_L g9606 ( 
.A(n_8762),
.Y(n_9606)
);

AND2x4_ASAP7_75t_L g9607 ( 
.A(n_9075),
.B(n_9080),
.Y(n_9607)
);

INVx2_ASAP7_75t_L g9608 ( 
.A(n_8768),
.Y(n_9608)
);

CKINVDCx20_ASAP7_75t_R g9609 ( 
.A(n_9181),
.Y(n_9609)
);

INVx1_ASAP7_75t_SL g9610 ( 
.A(n_9130),
.Y(n_9610)
);

OR2x2_ASAP7_75t_L g9611 ( 
.A(n_9265),
.B(n_6044),
.Y(n_9611)
);

AOI22xp33_ASAP7_75t_L g9612 ( 
.A1(n_8967),
.A2(n_9074),
.B1(n_9028),
.B2(n_8945),
.Y(n_9612)
);

INVx1_ASAP7_75t_L g9613 ( 
.A(n_9071),
.Y(n_9613)
);

INVx1_ASAP7_75t_L g9614 ( 
.A(n_8944),
.Y(n_9614)
);

INVx1_ASAP7_75t_L g9615 ( 
.A(n_8947),
.Y(n_9615)
);

INVx1_ASAP7_75t_L g9616 ( 
.A(n_8956),
.Y(n_9616)
);

INVx2_ASAP7_75t_L g9617 ( 
.A(n_8917),
.Y(n_9617)
);

INVx1_ASAP7_75t_L g9618 ( 
.A(n_8964),
.Y(n_9618)
);

INVx4_ASAP7_75t_L g9619 ( 
.A(n_9084),
.Y(n_9619)
);

AND2x4_ASAP7_75t_L g9620 ( 
.A(n_9163),
.B(n_5734),
.Y(n_9620)
);

NAND2xp5_ASAP7_75t_L g9621 ( 
.A(n_8816),
.B(n_6046),
.Y(n_9621)
);

BUFx2_ASAP7_75t_L g9622 ( 
.A(n_9291),
.Y(n_9622)
);

INVx1_ASAP7_75t_L g9623 ( 
.A(n_8970),
.Y(n_9623)
);

BUFx4f_ASAP7_75t_L g9624 ( 
.A(n_9260),
.Y(n_9624)
);

INVx1_ASAP7_75t_L g9625 ( 
.A(n_8973),
.Y(n_9625)
);

NOR2x1p5_ASAP7_75t_L g9626 ( 
.A(n_9294),
.B(n_6055),
.Y(n_9626)
);

INVx2_ASAP7_75t_L g9627 ( 
.A(n_8918),
.Y(n_9627)
);

BUFx6f_ASAP7_75t_L g9628 ( 
.A(n_9120),
.Y(n_9628)
);

INVx2_ASAP7_75t_L g9629 ( 
.A(n_8919),
.Y(n_9629)
);

INVx4_ASAP7_75t_L g9630 ( 
.A(n_9176),
.Y(n_9630)
);

INVx1_ASAP7_75t_L g9631 ( 
.A(n_8975),
.Y(n_9631)
);

NOR2xp33_ASAP7_75t_L g9632 ( 
.A(n_9262),
.B(n_6057),
.Y(n_9632)
);

HB1xp67_ASAP7_75t_L g9633 ( 
.A(n_9282),
.Y(n_9633)
);

NOR2xp33_ASAP7_75t_L g9634 ( 
.A(n_9183),
.B(n_6059),
.Y(n_9634)
);

BUFx2_ASAP7_75t_L g9635 ( 
.A(n_9266),
.Y(n_9635)
);

BUFx6f_ASAP7_75t_L g9636 ( 
.A(n_8926),
.Y(n_9636)
);

INVx1_ASAP7_75t_SL g9637 ( 
.A(n_9199),
.Y(n_9637)
);

NOR2xp33_ASAP7_75t_L g9638 ( 
.A(n_9134),
.B(n_6061),
.Y(n_9638)
);

NAND2xp5_ASAP7_75t_SL g9639 ( 
.A(n_8950),
.B(n_6064),
.Y(n_9639)
);

INVx3_ASAP7_75t_L g9640 ( 
.A(n_9263),
.Y(n_9640)
);

NOR2x1p5_ASAP7_75t_L g9641 ( 
.A(n_9301),
.B(n_6068),
.Y(n_9641)
);

BUFx3_ASAP7_75t_L g9642 ( 
.A(n_9223),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_8995),
.Y(n_9643)
);

BUFx10_ASAP7_75t_L g9644 ( 
.A(n_9310),
.Y(n_9644)
);

AND2x2_ASAP7_75t_L g9645 ( 
.A(n_8913),
.B(n_6070),
.Y(n_9645)
);

INVx1_ASAP7_75t_L g9646 ( 
.A(n_8999),
.Y(n_9646)
);

INVxp67_ASAP7_75t_L g9647 ( 
.A(n_8884),
.Y(n_9647)
);

BUFx3_ASAP7_75t_L g9648 ( 
.A(n_9272),
.Y(n_9648)
);

AND2x6_ASAP7_75t_L g9649 ( 
.A(n_9259),
.B(n_5737),
.Y(n_9649)
);

INVx2_ASAP7_75t_L g9650 ( 
.A(n_8924),
.Y(n_9650)
);

INVx3_ASAP7_75t_L g9651 ( 
.A(n_9256),
.Y(n_9651)
);

INVx1_ASAP7_75t_L g9652 ( 
.A(n_9000),
.Y(n_9652)
);

AOI22xp5_ASAP7_75t_SL g9653 ( 
.A1(n_8842),
.A2(n_6073),
.B1(n_6075),
.B2(n_6071),
.Y(n_9653)
);

NOR2xp33_ASAP7_75t_L g9654 ( 
.A(n_8864),
.B(n_6077),
.Y(n_9654)
);

OR2x2_ASAP7_75t_L g9655 ( 
.A(n_8892),
.B(n_6078),
.Y(n_9655)
);

INVx2_ASAP7_75t_L g9656 ( 
.A(n_8928),
.Y(n_9656)
);

AOI22xp33_ASAP7_75t_L g9657 ( 
.A1(n_9028),
.A2(n_5740),
.B1(n_5746),
.B2(n_5739),
.Y(n_9657)
);

INVx3_ASAP7_75t_L g9658 ( 
.A(n_9261),
.Y(n_9658)
);

NAND2xp5_ASAP7_75t_L g9659 ( 
.A(n_9031),
.B(n_6079),
.Y(n_9659)
);

AND2x4_ASAP7_75t_L g9660 ( 
.A(n_9252),
.B(n_5750),
.Y(n_9660)
);

INVx4_ASAP7_75t_L g9661 ( 
.A(n_8987),
.Y(n_9661)
);

INVx3_ASAP7_75t_L g9662 ( 
.A(n_9237),
.Y(n_9662)
);

NAND2xp5_ASAP7_75t_SL g9663 ( 
.A(n_8987),
.B(n_6083),
.Y(n_9663)
);

NOR2xp33_ASAP7_75t_L g9664 ( 
.A(n_8880),
.B(n_6084),
.Y(n_9664)
);

OR2x2_ASAP7_75t_L g9665 ( 
.A(n_9187),
.B(n_6085),
.Y(n_9665)
);

AOI22xp33_ASAP7_75t_L g9666 ( 
.A1(n_9028),
.A2(n_5754),
.B1(n_5763),
.B2(n_5752),
.Y(n_9666)
);

AND2x6_ASAP7_75t_L g9667 ( 
.A(n_9224),
.B(n_5765),
.Y(n_9667)
);

AOI22xp33_ASAP7_75t_L g9668 ( 
.A1(n_8941),
.A2(n_5781),
.B1(n_5782),
.B2(n_5766),
.Y(n_9668)
);

AOI22xp33_ASAP7_75t_L g9669 ( 
.A1(n_8949),
.A2(n_5787),
.B1(n_5789),
.B2(n_5783),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_SL g9670 ( 
.A(n_9021),
.B(n_6086),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_9007),
.Y(n_9671)
);

INVx1_ASAP7_75t_SL g9672 ( 
.A(n_9300),
.Y(n_9672)
);

INVx2_ASAP7_75t_SL g9673 ( 
.A(n_8834),
.Y(n_9673)
);

INVxp67_ASAP7_75t_SL g9674 ( 
.A(n_9064),
.Y(n_9674)
);

AND2x4_ASAP7_75t_L g9675 ( 
.A(n_9020),
.B(n_5793),
.Y(n_9675)
);

INVx1_ASAP7_75t_L g9676 ( 
.A(n_9190),
.Y(n_9676)
);

AND2x4_ASAP7_75t_L g9677 ( 
.A(n_9188),
.B(n_5794),
.Y(n_9677)
);

AND2x4_ASAP7_75t_L g9678 ( 
.A(n_9189),
.B(n_5795),
.Y(n_9678)
);

NOR2xp33_ASAP7_75t_L g9679 ( 
.A(n_9297),
.B(n_6088),
.Y(n_9679)
);

NAND2xp5_ASAP7_75t_L g9680 ( 
.A(n_8878),
.B(n_8955),
.Y(n_9680)
);

INVxp67_ASAP7_75t_SL g9681 ( 
.A(n_9087),
.Y(n_9681)
);

INVx2_ASAP7_75t_L g9682 ( 
.A(n_8933),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_8936),
.Y(n_9683)
);

CKINVDCx20_ASAP7_75t_R g9684 ( 
.A(n_9149),
.Y(n_9684)
);

INVx1_ASAP7_75t_L g9685 ( 
.A(n_8957),
.Y(n_9685)
);

NAND2xp33_ASAP7_75t_L g9686 ( 
.A(n_9216),
.B(n_6089),
.Y(n_9686)
);

INVx1_ASAP7_75t_L g9687 ( 
.A(n_8960),
.Y(n_9687)
);

NOR2xp33_ASAP7_75t_L g9688 ( 
.A(n_9137),
.B(n_6097),
.Y(n_9688)
);

INVx1_ASAP7_75t_L g9689 ( 
.A(n_8966),
.Y(n_9689)
);

OAI22xp5_ASAP7_75t_L g9690 ( 
.A1(n_9090),
.A2(n_6104),
.B1(n_6105),
.B2(n_6102),
.Y(n_9690)
);

NAND2xp5_ASAP7_75t_SL g9691 ( 
.A(n_8981),
.B(n_6107),
.Y(n_9691)
);

NOR2xp33_ASAP7_75t_L g9692 ( 
.A(n_9054),
.B(n_6110),
.Y(n_9692)
);

NOR2xp33_ASAP7_75t_L g9693 ( 
.A(n_8946),
.B(n_6114),
.Y(n_9693)
);

AND2x2_ASAP7_75t_L g9694 ( 
.A(n_8914),
.B(n_6115),
.Y(n_9694)
);

INVxp67_ASAP7_75t_L g9695 ( 
.A(n_8836),
.Y(n_9695)
);

NOR2xp33_ASAP7_75t_L g9696 ( 
.A(n_8901),
.B(n_8904),
.Y(n_9696)
);

NAND2xp33_ASAP7_75t_L g9697 ( 
.A(n_9151),
.B(n_9093),
.Y(n_9697)
);

INVx3_ASAP7_75t_L g9698 ( 
.A(n_9238),
.Y(n_9698)
);

AOI22xp33_ASAP7_75t_L g9699 ( 
.A1(n_8968),
.A2(n_5804),
.B1(n_5807),
.B2(n_5798),
.Y(n_9699)
);

INVx2_ASAP7_75t_SL g9700 ( 
.A(n_9240),
.Y(n_9700)
);

CKINVDCx5p33_ASAP7_75t_R g9701 ( 
.A(n_9044),
.Y(n_9701)
);

INVx4_ASAP7_75t_L g9702 ( 
.A(n_9203),
.Y(n_9702)
);

INVx2_ASAP7_75t_L g9703 ( 
.A(n_8972),
.Y(n_9703)
);

CKINVDCx5p33_ASAP7_75t_R g9704 ( 
.A(n_9195),
.Y(n_9704)
);

NAND2xp5_ASAP7_75t_SL g9705 ( 
.A(n_8765),
.B(n_6117),
.Y(n_9705)
);

INVx4_ASAP7_75t_L g9706 ( 
.A(n_8807),
.Y(n_9706)
);

BUFx3_ASAP7_75t_L g9707 ( 
.A(n_9288),
.Y(n_9707)
);

NAND2xp5_ASAP7_75t_L g9708 ( 
.A(n_8976),
.B(n_6123),
.Y(n_9708)
);

NAND2xp5_ASAP7_75t_L g9709 ( 
.A(n_8977),
.B(n_6125),
.Y(n_9709)
);

NOR2xp33_ASAP7_75t_L g9710 ( 
.A(n_8942),
.B(n_6129),
.Y(n_9710)
);

AND2x2_ASAP7_75t_L g9711 ( 
.A(n_8927),
.B(n_6132),
.Y(n_9711)
);

BUFx3_ASAP7_75t_L g9712 ( 
.A(n_9284),
.Y(n_9712)
);

BUFx3_ASAP7_75t_L g9713 ( 
.A(n_9287),
.Y(n_9713)
);

NAND2xp5_ASAP7_75t_SL g9714 ( 
.A(n_9088),
.B(n_6134),
.Y(n_9714)
);

AND2x2_ASAP7_75t_L g9715 ( 
.A(n_8908),
.B(n_6135),
.Y(n_9715)
);

NAND2xp5_ASAP7_75t_SL g9716 ( 
.A(n_9268),
.B(n_6137),
.Y(n_9716)
);

AND2x2_ASAP7_75t_L g9717 ( 
.A(n_8874),
.B(n_6138),
.Y(n_9717)
);

INVx2_ASAP7_75t_L g9718 ( 
.A(n_8978),
.Y(n_9718)
);

INVx2_ASAP7_75t_L g9719 ( 
.A(n_8983),
.Y(n_9719)
);

INVx1_ASAP7_75t_L g9720 ( 
.A(n_8985),
.Y(n_9720)
);

AND2x2_ASAP7_75t_L g9721 ( 
.A(n_9225),
.B(n_6139),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_8991),
.Y(n_9722)
);

BUFx10_ASAP7_75t_L g9723 ( 
.A(n_8859),
.Y(n_9723)
);

INVx2_ASAP7_75t_SL g9724 ( 
.A(n_9239),
.Y(n_9724)
);

INVx1_ASAP7_75t_L g9725 ( 
.A(n_8994),
.Y(n_9725)
);

INVx3_ASAP7_75t_L g9726 ( 
.A(n_9191),
.Y(n_9726)
);

INVx4_ASAP7_75t_L g9727 ( 
.A(n_9295),
.Y(n_9727)
);

INVx5_ASAP7_75t_L g9728 ( 
.A(n_8836),
.Y(n_9728)
);

INVx3_ASAP7_75t_L g9729 ( 
.A(n_9192),
.Y(n_9729)
);

AND3x4_ASAP7_75t_L g9730 ( 
.A(n_9308),
.B(n_6144),
.C(n_6140),
.Y(n_9730)
);

NOR2xp33_ASAP7_75t_L g9731 ( 
.A(n_8951),
.B(n_8959),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_8996),
.Y(n_9732)
);

AND2x2_ASAP7_75t_L g9733 ( 
.A(n_8796),
.B(n_8810),
.Y(n_9733)
);

BUFx6f_ASAP7_75t_L g9734 ( 
.A(n_9056),
.Y(n_9734)
);

INVx2_ASAP7_75t_L g9735 ( 
.A(n_8997),
.Y(n_9735)
);

INVx2_ASAP7_75t_L g9736 ( 
.A(n_9004),
.Y(n_9736)
);

NAND2xp5_ASAP7_75t_SL g9737 ( 
.A(n_9073),
.B(n_6145),
.Y(n_9737)
);

INVx2_ASAP7_75t_SL g9738 ( 
.A(n_9208),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_9011),
.Y(n_9739)
);

INVx2_ASAP7_75t_L g9740 ( 
.A(n_9012),
.Y(n_9740)
);

NAND2xp33_ASAP7_75t_L g9741 ( 
.A(n_9098),
.B(n_6146),
.Y(n_9741)
);

HB1xp67_ASAP7_75t_L g9742 ( 
.A(n_9122),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_9013),
.Y(n_9743)
);

INVx2_ASAP7_75t_L g9744 ( 
.A(n_9016),
.Y(n_9744)
);

NAND2xp33_ASAP7_75t_L g9745 ( 
.A(n_9099),
.B(n_6148),
.Y(n_9745)
);

AND2x4_ASAP7_75t_L g9746 ( 
.A(n_9210),
.B(n_5819),
.Y(n_9746)
);

INVx1_ASAP7_75t_L g9747 ( 
.A(n_9017),
.Y(n_9747)
);

NAND2xp5_ASAP7_75t_L g9748 ( 
.A(n_9019),
.B(n_6151),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_9025),
.Y(n_9749)
);

NAND2xp5_ASAP7_75t_SL g9750 ( 
.A(n_9027),
.B(n_6153),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_L g9751 ( 
.A(n_9029),
.B(n_6155),
.Y(n_9751)
);

NAND2xp5_ASAP7_75t_L g9752 ( 
.A(n_9030),
.B(n_6156),
.Y(n_9752)
);

NAND2xp5_ASAP7_75t_L g9753 ( 
.A(n_9036),
.B(n_6157),
.Y(n_9753)
);

NAND2xp5_ASAP7_75t_L g9754 ( 
.A(n_9038),
.B(n_6158),
.Y(n_9754)
);

INVx1_ASAP7_75t_L g9755 ( 
.A(n_9043),
.Y(n_9755)
);

INVxp67_ASAP7_75t_L g9756 ( 
.A(n_9122),
.Y(n_9756)
);

BUFx2_ASAP7_75t_L g9757 ( 
.A(n_9109),
.Y(n_9757)
);

NAND2xp5_ASAP7_75t_SL g9758 ( 
.A(n_9048),
.B(n_6159),
.Y(n_9758)
);

AND2x2_ASAP7_75t_L g9759 ( 
.A(n_8815),
.B(n_6161),
.Y(n_9759)
);

INVx3_ASAP7_75t_L g9760 ( 
.A(n_9214),
.Y(n_9760)
);

INVx1_ASAP7_75t_L g9761 ( 
.A(n_9049),
.Y(n_9761)
);

NOR2xp33_ASAP7_75t_L g9762 ( 
.A(n_9311),
.B(n_8820),
.Y(n_9762)
);

AND2x4_ASAP7_75t_L g9763 ( 
.A(n_9218),
.B(n_5825),
.Y(n_9763)
);

BUFx3_ASAP7_75t_L g9764 ( 
.A(n_9220),
.Y(n_9764)
);

AND2x2_ASAP7_75t_L g9765 ( 
.A(n_8835),
.B(n_6164),
.Y(n_9765)
);

NOR2xp33_ASAP7_75t_L g9766 ( 
.A(n_9281),
.B(n_6169),
.Y(n_9766)
);

INVx3_ASAP7_75t_L g9767 ( 
.A(n_9222),
.Y(n_9767)
);

CKINVDCx5p33_ASAP7_75t_R g9768 ( 
.A(n_9305),
.Y(n_9768)
);

AND2x2_ASAP7_75t_SL g9769 ( 
.A(n_9124),
.B(n_5830),
.Y(n_9769)
);

HB1xp67_ASAP7_75t_L g9770 ( 
.A(n_9096),
.Y(n_9770)
);

INVx2_ASAP7_75t_L g9771 ( 
.A(n_9051),
.Y(n_9771)
);

BUFx2_ASAP7_75t_L g9772 ( 
.A(n_9280),
.Y(n_9772)
);

INVx3_ASAP7_75t_L g9773 ( 
.A(n_9229),
.Y(n_9773)
);

INVxp67_ASAP7_75t_L g9774 ( 
.A(n_9242),
.Y(n_9774)
);

BUFx6f_ASAP7_75t_L g9775 ( 
.A(n_9247),
.Y(n_9775)
);

OAI22xp5_ASAP7_75t_SL g9776 ( 
.A1(n_9302),
.A2(n_6176),
.B1(n_6180),
.B2(n_6172),
.Y(n_9776)
);

INVx2_ASAP7_75t_L g9777 ( 
.A(n_9055),
.Y(n_9777)
);

BUFx6f_ASAP7_75t_L g9778 ( 
.A(n_8769),
.Y(n_9778)
);

INVx2_ASAP7_75t_SL g9779 ( 
.A(n_9243),
.Y(n_9779)
);

INVxp33_ASAP7_75t_L g9780 ( 
.A(n_9292),
.Y(n_9780)
);

BUFx2_ASAP7_75t_L g9781 ( 
.A(n_9138),
.Y(n_9781)
);

NAND2xp5_ASAP7_75t_L g9782 ( 
.A(n_9068),
.B(n_6181),
.Y(n_9782)
);

INVx3_ASAP7_75t_L g9783 ( 
.A(n_9172),
.Y(n_9783)
);

BUFx6f_ASAP7_75t_L g9784 ( 
.A(n_9175),
.Y(n_9784)
);

NOR2xp33_ASAP7_75t_L g9785 ( 
.A(n_8984),
.B(n_6184),
.Y(n_9785)
);

INVx1_ASAP7_75t_L g9786 ( 
.A(n_9072),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_9076),
.Y(n_9787)
);

CKINVDCx5p33_ASAP7_75t_R g9788 ( 
.A(n_9303),
.Y(n_9788)
);

AOI22xp33_ASAP7_75t_L g9789 ( 
.A1(n_9078),
.A2(n_5834),
.B1(n_5842),
.B2(n_5831),
.Y(n_9789)
);

CKINVDCx5p33_ASAP7_75t_R g9790 ( 
.A(n_9306),
.Y(n_9790)
);

INVx1_ASAP7_75t_L g9791 ( 
.A(n_9082),
.Y(n_9791)
);

INVx1_ASAP7_75t_L g9792 ( 
.A(n_9094),
.Y(n_9792)
);

INVx1_ASAP7_75t_L g9793 ( 
.A(n_9095),
.Y(n_9793)
);

OR2x2_ASAP7_75t_L g9794 ( 
.A(n_9106),
.B(n_6187),
.Y(n_9794)
);

BUFx3_ASAP7_75t_L g9795 ( 
.A(n_9257),
.Y(n_9795)
);

INVx1_ASAP7_75t_L g9796 ( 
.A(n_9140),
.Y(n_9796)
);

BUFx6f_ASAP7_75t_L g9797 ( 
.A(n_9177),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_9145),
.Y(n_9798)
);

INVx1_ASAP7_75t_L g9799 ( 
.A(n_9147),
.Y(n_9799)
);

INVx1_ASAP7_75t_L g9800 ( 
.A(n_9153),
.Y(n_9800)
);

INVx2_ASAP7_75t_L g9801 ( 
.A(n_8813),
.Y(n_9801)
);

AND2x4_ASAP7_75t_L g9802 ( 
.A(n_9178),
.B(n_5847),
.Y(n_9802)
);

INVx2_ASAP7_75t_L g9803 ( 
.A(n_9155),
.Y(n_9803)
);

NAND2xp5_ASAP7_75t_SL g9804 ( 
.A(n_9148),
.B(n_6189),
.Y(n_9804)
);

AND2x4_ASAP7_75t_L g9805 ( 
.A(n_9227),
.B(n_5849),
.Y(n_9805)
);

AND2x4_ASAP7_75t_L g9806 ( 
.A(n_9228),
.B(n_5850),
.Y(n_9806)
);

INVx1_ASAP7_75t_L g9807 ( 
.A(n_9156),
.Y(n_9807)
);

INVx1_ASAP7_75t_L g9808 ( 
.A(n_9157),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_9063),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_8974),
.Y(n_9810)
);

INVx4_ASAP7_75t_SL g9811 ( 
.A(n_8989),
.Y(n_9811)
);

AND2x4_ASAP7_75t_L g9812 ( 
.A(n_9232),
.B(n_5859),
.Y(n_9812)
);

NOR2xp33_ASAP7_75t_L g9813 ( 
.A(n_8993),
.B(n_6196),
.Y(n_9813)
);

AND2x6_ASAP7_75t_L g9814 ( 
.A(n_8863),
.B(n_5873),
.Y(n_9814)
);

OR2x6_ASAP7_75t_L g9815 ( 
.A(n_8989),
.B(n_5874),
.Y(n_9815)
);

INVx1_ASAP7_75t_SL g9816 ( 
.A(n_9213),
.Y(n_9816)
);

AOI22xp33_ASAP7_75t_L g9817 ( 
.A1(n_9235),
.A2(n_5882),
.B1(n_5885),
.B2(n_5881),
.Y(n_9817)
);

NOR2xp33_ASAP7_75t_L g9818 ( 
.A(n_9040),
.B(n_6198),
.Y(n_9818)
);

AO22x2_ASAP7_75t_L g9819 ( 
.A1(n_8779),
.A2(n_5896),
.B1(n_5901),
.B2(n_5891),
.Y(n_9819)
);

AND2x6_ASAP7_75t_L g9820 ( 
.A(n_8872),
.B(n_5907),
.Y(n_9820)
);

AOI22xp33_ASAP7_75t_L g9821 ( 
.A1(n_8808),
.A2(n_5914),
.B1(n_5921),
.B2(n_5911),
.Y(n_9821)
);

AND2x4_ASAP7_75t_L g9822 ( 
.A(n_9267),
.B(n_5935),
.Y(n_9822)
);

INVx1_ASAP7_75t_L g9823 ( 
.A(n_9085),
.Y(n_9823)
);

NOR2xp67_ASAP7_75t_L g9824 ( 
.A(n_9396),
.B(n_9116),
.Y(n_9824)
);

NAND2xp5_ASAP7_75t_L g9825 ( 
.A(n_9343),
.B(n_9115),
.Y(n_9825)
);

INVxp67_ASAP7_75t_L g9826 ( 
.A(n_9332),
.Y(n_9826)
);

NAND2xp5_ASAP7_75t_L g9827 ( 
.A(n_9500),
.B(n_8954),
.Y(n_9827)
);

NAND2xp5_ASAP7_75t_L g9828 ( 
.A(n_9316),
.B(n_8788),
.Y(n_9828)
);

NAND2xp5_ASAP7_75t_L g9829 ( 
.A(n_9399),
.B(n_8851),
.Y(n_9829)
);

INVx2_ASAP7_75t_L g9830 ( 
.A(n_9317),
.Y(n_9830)
);

INVx2_ASAP7_75t_SL g9831 ( 
.A(n_9400),
.Y(n_9831)
);

NAND2xp5_ASAP7_75t_SL g9832 ( 
.A(n_9366),
.B(n_8882),
.Y(n_9832)
);

INVx1_ASAP7_75t_L g9833 ( 
.A(n_9325),
.Y(n_9833)
);

NAND2xp5_ASAP7_75t_L g9834 ( 
.A(n_9388),
.B(n_8910),
.Y(n_9834)
);

INVx2_ASAP7_75t_L g9835 ( 
.A(n_9334),
.Y(n_9835)
);

NAND2xp5_ASAP7_75t_L g9836 ( 
.A(n_9491),
.B(n_9050),
.Y(n_9836)
);

OR2x2_ASAP7_75t_L g9837 ( 
.A(n_9480),
.B(n_9062),
.Y(n_9837)
);

NAND2xp5_ASAP7_75t_L g9838 ( 
.A(n_9507),
.B(n_9198),
.Y(n_9838)
);

NAND2xp5_ASAP7_75t_L g9839 ( 
.A(n_9510),
.B(n_9128),
.Y(n_9839)
);

BUFx3_ASAP7_75t_L g9840 ( 
.A(n_9425),
.Y(n_9840)
);

INVx1_ASAP7_75t_L g9841 ( 
.A(n_9351),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_9353),
.Y(n_9842)
);

AND2x4_ASAP7_75t_L g9843 ( 
.A(n_9318),
.B(n_9173),
.Y(n_9843)
);

NAND2xp5_ASAP7_75t_L g9844 ( 
.A(n_9520),
.B(n_9139),
.Y(n_9844)
);

AOI22xp5_ASAP7_75t_L g9845 ( 
.A1(n_9679),
.A2(n_9042),
.B1(n_9059),
.B2(n_9131),
.Y(n_9845)
);

NOR2xp33_ASAP7_75t_L g9846 ( 
.A(n_9392),
.B(n_9246),
.Y(n_9846)
);

NAND2xp5_ASAP7_75t_L g9847 ( 
.A(n_9534),
.B(n_8900),
.Y(n_9847)
);

INVx4_ASAP7_75t_L g9848 ( 
.A(n_9400),
.Y(n_9848)
);

NAND2xp5_ASAP7_75t_SL g9849 ( 
.A(n_9477),
.B(n_9089),
.Y(n_9849)
);

INVx1_ASAP7_75t_L g9850 ( 
.A(n_9356),
.Y(n_9850)
);

AOI22xp5_ASAP7_75t_L g9851 ( 
.A1(n_9487),
.A2(n_9154),
.B1(n_9307),
.B2(n_9185),
.Y(n_9851)
);

INVx1_ASAP7_75t_L g9852 ( 
.A(n_9357),
.Y(n_9852)
);

NOR2xp33_ASAP7_75t_L g9853 ( 
.A(n_9774),
.B(n_9250),
.Y(n_9853)
);

NAND2xp5_ASAP7_75t_L g9854 ( 
.A(n_9565),
.B(n_9255),
.Y(n_9854)
);

AOI22xp33_ASAP7_75t_L g9855 ( 
.A1(n_9692),
.A2(n_9285),
.B1(n_9234),
.B2(n_9168),
.Y(n_9855)
);

INVx2_ASAP7_75t_L g9856 ( 
.A(n_9373),
.Y(n_9856)
);

NOR2xp33_ASAP7_75t_L g9857 ( 
.A(n_9664),
.B(n_9278),
.Y(n_9857)
);

BUFx6f_ASAP7_75t_L g9858 ( 
.A(n_9376),
.Y(n_9858)
);

NOR3xp33_ASAP7_75t_L g9859 ( 
.A(n_9693),
.B(n_9182),
.C(n_9158),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9580),
.B(n_9244),
.Y(n_9860)
);

NAND2xp5_ASAP7_75t_L g9861 ( 
.A(n_9634),
.B(n_9322),
.Y(n_9861)
);

XOR2xp5_ASAP7_75t_L g9862 ( 
.A(n_9402),
.B(n_9304),
.Y(n_9862)
);

INVx1_ASAP7_75t_L g9863 ( 
.A(n_9381),
.Y(n_9863)
);

NAND2xp5_ASAP7_75t_L g9864 ( 
.A(n_9348),
.B(n_9206),
.Y(n_9864)
);

NOR2xp33_ASAP7_75t_L g9865 ( 
.A(n_9315),
.B(n_9069),
.Y(n_9865)
);

NOR2xp33_ASAP7_75t_L g9866 ( 
.A(n_9688),
.B(n_9077),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_9386),
.Y(n_9867)
);

NAND2xp5_ASAP7_75t_L g9868 ( 
.A(n_9355),
.B(n_9363),
.Y(n_9868)
);

INVx3_ASAP7_75t_L g9869 ( 
.A(n_9497),
.Y(n_9869)
);

HB1xp67_ASAP7_75t_L g9870 ( 
.A(n_9314),
.Y(n_9870)
);

BUFx3_ASAP7_75t_L g9871 ( 
.A(n_9377),
.Y(n_9871)
);

NAND2xp5_ASAP7_75t_L g9872 ( 
.A(n_9638),
.B(n_9170),
.Y(n_9872)
);

BUFx3_ASAP7_75t_L g9873 ( 
.A(n_9362),
.Y(n_9873)
);

INVx1_ASAP7_75t_L g9874 ( 
.A(n_9395),
.Y(n_9874)
);

AOI22xp33_ASAP7_75t_SL g9875 ( 
.A1(n_9592),
.A2(n_9302),
.B1(n_6201),
.B2(n_6204),
.Y(n_9875)
);

NAND2xp5_ASAP7_75t_L g9876 ( 
.A(n_9602),
.B(n_9160),
.Y(n_9876)
);

OAI221xp5_ASAP7_75t_L g9877 ( 
.A1(n_9439),
.A2(n_5943),
.B1(n_5945),
.B2(n_5941),
.C(n_5940),
.Y(n_9877)
);

NAND2xp5_ASAP7_75t_L g9878 ( 
.A(n_9711),
.B(n_9715),
.Y(n_9878)
);

NAND2xp5_ASAP7_75t_L g9879 ( 
.A(n_9717),
.B(n_9231),
.Y(n_9879)
);

AOI22xp5_ASAP7_75t_L g9880 ( 
.A1(n_9408),
.A2(n_9290),
.B1(n_9022),
.B2(n_9219),
.Y(n_9880)
);

AOI22xp33_ASAP7_75t_L g9881 ( 
.A1(n_9403),
.A2(n_9186),
.B1(n_5948),
.B2(n_5950),
.Y(n_9881)
);

INVx1_ASAP7_75t_L g9882 ( 
.A(n_9404),
.Y(n_9882)
);

NOR2xp33_ASAP7_75t_L g9883 ( 
.A(n_9647),
.B(n_8826),
.Y(n_9883)
);

BUFx3_ASAP7_75t_L g9884 ( 
.A(n_9401),
.Y(n_9884)
);

NAND2xp5_ASAP7_75t_SL g9885 ( 
.A(n_9624),
.B(n_6200),
.Y(n_9885)
);

INVx8_ASAP7_75t_L g9886 ( 
.A(n_9323),
.Y(n_9886)
);

NAND2xp5_ASAP7_75t_L g9887 ( 
.A(n_9632),
.B(n_5946),
.Y(n_9887)
);

INVx1_ASAP7_75t_L g9888 ( 
.A(n_9410),
.Y(n_9888)
);

AOI22xp33_ASAP7_75t_L g9889 ( 
.A1(n_9769),
.A2(n_5952),
.B1(n_5954),
.B2(n_5951),
.Y(n_9889)
);

NAND2xp5_ASAP7_75t_L g9890 ( 
.A(n_9375),
.B(n_5958),
.Y(n_9890)
);

O2A1O1Ixp33_ASAP7_75t_L g9891 ( 
.A1(n_9544),
.A2(n_5971),
.B(n_5979),
.C(n_5965),
.Y(n_9891)
);

NAND2xp5_ASAP7_75t_L g9892 ( 
.A(n_9766),
.B(n_5982),
.Y(n_9892)
);

NAND2xp5_ASAP7_75t_L g9893 ( 
.A(n_9645),
.B(n_5995),
.Y(n_9893)
);

NAND2xp5_ASAP7_75t_L g9894 ( 
.A(n_9694),
.B(n_9571),
.Y(n_9894)
);

AOI22xp5_ASAP7_75t_L g9895 ( 
.A1(n_9696),
.A2(n_6207),
.B1(n_6208),
.B2(n_6206),
.Y(n_9895)
);

INVx1_ASAP7_75t_L g9896 ( 
.A(n_9413),
.Y(n_9896)
);

INVx2_ASAP7_75t_L g9897 ( 
.A(n_9420),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_L g9898 ( 
.A(n_9458),
.B(n_5999),
.Y(n_9898)
);

INVx2_ASAP7_75t_L g9899 ( 
.A(n_9443),
.Y(n_9899)
);

NOR2xp33_ASAP7_75t_L g9900 ( 
.A(n_9568),
.B(n_6210),
.Y(n_9900)
);

NAND2xp5_ASAP7_75t_L g9901 ( 
.A(n_9528),
.B(n_6002),
.Y(n_9901)
);

NAND2xp5_ASAP7_75t_SL g9902 ( 
.A(n_9573),
.B(n_6212),
.Y(n_9902)
);

AOI21xp5_ASAP7_75t_L g9903 ( 
.A1(n_9680),
.A2(n_9166),
.B(n_9165),
.Y(n_9903)
);

NAND2xp5_ASAP7_75t_L g9904 ( 
.A(n_9566),
.B(n_6008),
.Y(n_9904)
);

NAND2xp5_ASAP7_75t_L g9905 ( 
.A(n_9567),
.B(n_6019),
.Y(n_9905)
);

O2A1O1Ixp33_ASAP7_75t_L g9906 ( 
.A1(n_9341),
.A2(n_6034),
.B(n_6035),
.C(n_6032),
.Y(n_9906)
);

BUFx8_ASAP7_75t_L g9907 ( 
.A(n_9557),
.Y(n_9907)
);

BUFx5_ASAP7_75t_L g9908 ( 
.A(n_9810),
.Y(n_9908)
);

INVx2_ASAP7_75t_L g9909 ( 
.A(n_9447),
.Y(n_9909)
);

AOI22xp33_ASAP7_75t_L g9910 ( 
.A1(n_9710),
.A2(n_6050),
.B1(n_6051),
.B2(n_6037),
.Y(n_9910)
);

NAND2xp5_ASAP7_75t_L g9911 ( 
.A(n_9574),
.B(n_6058),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_9451),
.Y(n_9912)
);

INVx2_ASAP7_75t_L g9913 ( 
.A(n_9452),
.Y(n_9913)
);

INVx1_ASAP7_75t_L g9914 ( 
.A(n_9456),
.Y(n_9914)
);

NAND2xp5_ASAP7_75t_SL g9915 ( 
.A(n_9768),
.B(n_6213),
.Y(n_9915)
);

AOI22xp5_ASAP7_75t_L g9916 ( 
.A1(n_9731),
.A2(n_6216),
.B1(n_6220),
.B2(n_6214),
.Y(n_9916)
);

NAND3xp33_ASAP7_75t_L g9917 ( 
.A(n_9459),
.B(n_6225),
.C(n_6222),
.Y(n_9917)
);

NAND2xp5_ASAP7_75t_L g9918 ( 
.A(n_9590),
.B(n_6062),
.Y(n_9918)
);

CKINVDCx5p33_ASAP7_75t_R g9919 ( 
.A(n_9358),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_9457),
.Y(n_9920)
);

NAND2xp5_ASAP7_75t_L g9921 ( 
.A(n_9621),
.B(n_6063),
.Y(n_9921)
);

NOR3xp33_ASAP7_75t_L g9922 ( 
.A(n_9523),
.B(n_6069),
.C(n_6065),
.Y(n_9922)
);

AND2x2_ASAP7_75t_L g9923 ( 
.A(n_9336),
.B(n_6226),
.Y(n_9923)
);

NAND2xp5_ASAP7_75t_L g9924 ( 
.A(n_9349),
.B(n_6072),
.Y(n_9924)
);

NAND2xp5_ASAP7_75t_SL g9925 ( 
.A(n_9576),
.B(n_6231),
.Y(n_9925)
);

NAND2xp5_ASAP7_75t_SL g9926 ( 
.A(n_9788),
.B(n_6232),
.Y(n_9926)
);

INVx1_ASAP7_75t_L g9927 ( 
.A(n_9479),
.Y(n_9927)
);

INVx2_ASAP7_75t_L g9928 ( 
.A(n_9486),
.Y(n_9928)
);

INVx1_ASAP7_75t_L g9929 ( 
.A(n_9490),
.Y(n_9929)
);

INVx1_ASAP7_75t_L g9930 ( 
.A(n_9494),
.Y(n_9930)
);

NOR3xp33_ASAP7_75t_L g9931 ( 
.A(n_9705),
.B(n_6082),
.C(n_6074),
.Y(n_9931)
);

OR2x2_ASAP7_75t_SL g9932 ( 
.A(n_9333),
.B(n_6093),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_9495),
.Y(n_9933)
);

INVx8_ASAP7_75t_L g9934 ( 
.A(n_9323),
.Y(n_9934)
);

INVx1_ASAP7_75t_SL g9935 ( 
.A(n_9319),
.Y(n_9935)
);

NAND2xp5_ASAP7_75t_L g9936 ( 
.A(n_9359),
.B(n_6101),
.Y(n_9936)
);

NAND2xp5_ASAP7_75t_L g9937 ( 
.A(n_9360),
.B(n_6106),
.Y(n_9937)
);

NAND2xp5_ASAP7_75t_L g9938 ( 
.A(n_9484),
.B(n_6108),
.Y(n_9938)
);

NOR2xp33_ASAP7_75t_L g9939 ( 
.A(n_9610),
.B(n_6233),
.Y(n_9939)
);

INVxp67_ASAP7_75t_L g9940 ( 
.A(n_9559),
.Y(n_9940)
);

INVx1_ASAP7_75t_L g9941 ( 
.A(n_9496),
.Y(n_9941)
);

NAND2xp5_ASAP7_75t_L g9942 ( 
.A(n_9681),
.B(n_6119),
.Y(n_9942)
);

INVx1_ASAP7_75t_L g9943 ( 
.A(n_9502),
.Y(n_9943)
);

NAND2xp5_ASAP7_75t_SL g9944 ( 
.A(n_9790),
.B(n_6236),
.Y(n_9944)
);

BUFx6f_ASAP7_75t_SL g9945 ( 
.A(n_9321),
.Y(n_9945)
);

NAND2xp5_ASAP7_75t_SL g9946 ( 
.A(n_9728),
.B(n_9470),
.Y(n_9946)
);

A2O1A1Ixp33_ASAP7_75t_L g9947 ( 
.A1(n_9762),
.A2(n_6121),
.B(n_6124),
.C(n_6120),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_L g9948 ( 
.A(n_9498),
.B(n_6126),
.Y(n_9948)
);

BUFx3_ASAP7_75t_L g9949 ( 
.A(n_9412),
.Y(n_9949)
);

NOR2xp33_ASAP7_75t_L g9950 ( 
.A(n_9780),
.B(n_6237),
.Y(n_9950)
);

NAND2xp5_ASAP7_75t_L g9951 ( 
.A(n_9505),
.B(n_6130),
.Y(n_9951)
);

AND2x2_ASAP7_75t_L g9952 ( 
.A(n_9383),
.B(n_6238),
.Y(n_9952)
);

NOR2xp67_ASAP7_75t_L g9953 ( 
.A(n_9640),
.B(n_4585),
.Y(n_9953)
);

NAND2xp5_ASAP7_75t_SL g9954 ( 
.A(n_9728),
.B(n_9470),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9482),
.B(n_6133),
.Y(n_9955)
);

INVx2_ASAP7_75t_L g9956 ( 
.A(n_9553),
.Y(n_9956)
);

NOR2xp67_ASAP7_75t_L g9957 ( 
.A(n_9342),
.B(n_4587),
.Y(n_9957)
);

NAND2xp5_ASAP7_75t_SL g9958 ( 
.A(n_9492),
.B(n_6240),
.Y(n_9958)
);

AOI22xp33_ASAP7_75t_L g9959 ( 
.A1(n_9785),
.A2(n_6163),
.B1(n_6171),
.B2(n_6143),
.Y(n_9959)
);

INVx2_ASAP7_75t_L g9960 ( 
.A(n_9560),
.Y(n_9960)
);

NAND2xp5_ASAP7_75t_L g9961 ( 
.A(n_9364),
.B(n_9676),
.Y(n_9961)
);

INVx2_ASAP7_75t_L g9962 ( 
.A(n_9563),
.Y(n_9962)
);

INVx1_ASAP7_75t_L g9963 ( 
.A(n_9575),
.Y(n_9963)
);

AND2x4_ASAP7_75t_SL g9964 ( 
.A(n_9324),
.B(n_6173),
.Y(n_9964)
);

AND2x4_ASAP7_75t_L g9965 ( 
.A(n_9466),
.B(n_6174),
.Y(n_9965)
);

INVx2_ASAP7_75t_L g9966 ( 
.A(n_9582),
.Y(n_9966)
);

NAND2xp5_ASAP7_75t_SL g9967 ( 
.A(n_9492),
.B(n_6242),
.Y(n_9967)
);

AO221x1_ASAP7_75t_L g9968 ( 
.A1(n_9819),
.A2(n_6183),
.B1(n_6185),
.B2(n_6182),
.C(n_6179),
.Y(n_9968)
);

NAND2xp5_ASAP7_75t_SL g9969 ( 
.A(n_9816),
.B(n_6247),
.Y(n_9969)
);

OAI22xp5_ASAP7_75t_L g9970 ( 
.A1(n_9488),
.A2(n_6249),
.B1(n_6250),
.B2(n_6248),
.Y(n_9970)
);

NAND2xp5_ASAP7_75t_L g9971 ( 
.A(n_9380),
.B(n_6188),
.Y(n_9971)
);

NAND2xp5_ASAP7_75t_SL g9972 ( 
.A(n_9727),
.B(n_6253),
.Y(n_9972)
);

INVx3_ASAP7_75t_L g9973 ( 
.A(n_9562),
.Y(n_9973)
);

NAND2xp5_ASAP7_75t_L g9974 ( 
.A(n_9513),
.B(n_6191),
.Y(n_9974)
);

NOR2xp33_ASAP7_75t_L g9975 ( 
.A(n_9555),
.B(n_6260),
.Y(n_9975)
);

AOI22xp5_ASAP7_75t_L g9976 ( 
.A1(n_9450),
.A2(n_6268),
.B1(n_6270),
.B2(n_6264),
.Y(n_9976)
);

NAND2xp5_ASAP7_75t_L g9977 ( 
.A(n_9518),
.B(n_6194),
.Y(n_9977)
);

INVx1_ASAP7_75t_L g9978 ( 
.A(n_9583),
.Y(n_9978)
);

NAND2xp5_ASAP7_75t_L g9979 ( 
.A(n_9521),
.B(n_9527),
.Y(n_9979)
);

NAND2xp5_ASAP7_75t_SL g9980 ( 
.A(n_9644),
.B(n_6271),
.Y(n_9980)
);

AOI22xp5_ASAP7_75t_L g9981 ( 
.A1(n_9724),
.A2(n_6275),
.B1(n_6276),
.B2(n_6274),
.Y(n_9981)
);

INVx2_ASAP7_75t_L g9982 ( 
.A(n_9584),
.Y(n_9982)
);

INVx2_ASAP7_75t_L g9983 ( 
.A(n_9585),
.Y(n_9983)
);

NAND2xp33_ASAP7_75t_L g9984 ( 
.A(n_9368),
.B(n_6279),
.Y(n_9984)
);

NAND2xp5_ASAP7_75t_SL g9985 ( 
.A(n_9637),
.B(n_6284),
.Y(n_9985)
);

INVxp67_ASAP7_75t_L g9986 ( 
.A(n_9622),
.Y(n_9986)
);

AOI221xp5_ASAP7_75t_L g9987 ( 
.A1(n_9339),
.A2(n_6202),
.B1(n_6205),
.B2(n_6199),
.C(n_6197),
.Y(n_9987)
);

NAND2xp5_ASAP7_75t_L g9988 ( 
.A(n_9530),
.B(n_6209),
.Y(n_9988)
);

OAI22xp5_ASAP7_75t_L g9989 ( 
.A1(n_9674),
.A2(n_6289),
.B1(n_6295),
.B2(n_6288),
.Y(n_9989)
);

NAND2xp5_ASAP7_75t_L g9990 ( 
.A(n_9531),
.B(n_6223),
.Y(n_9990)
);

NOR2xp33_ASAP7_75t_L g9991 ( 
.A(n_9706),
.B(n_6297),
.Y(n_9991)
);

INVx2_ASAP7_75t_L g9992 ( 
.A(n_9589),
.Y(n_9992)
);

AOI22xp33_ASAP7_75t_L g9993 ( 
.A1(n_9813),
.A2(n_6234),
.B1(n_6235),
.B2(n_6230),
.Y(n_9993)
);

NAND2xp5_ASAP7_75t_L g9994 ( 
.A(n_9542),
.B(n_6241),
.Y(n_9994)
);

NAND2xp5_ASAP7_75t_L g9995 ( 
.A(n_9545),
.B(n_6244),
.Y(n_9995)
);

AND2x2_ASAP7_75t_L g9996 ( 
.A(n_9535),
.B(n_6298),
.Y(n_9996)
);

INVx1_ASAP7_75t_L g9997 ( 
.A(n_9594),
.Y(n_9997)
);

INVx1_ASAP7_75t_L g9998 ( 
.A(n_9596),
.Y(n_9998)
);

AOI22xp5_ASAP7_75t_L g9999 ( 
.A1(n_9654),
.A2(n_6302),
.B1(n_6305),
.B2(n_6300),
.Y(n_9999)
);

INVx5_ASAP7_75t_L g10000 ( 
.A(n_9367),
.Y(n_10000)
);

AOI22xp5_ASAP7_75t_L g10001 ( 
.A1(n_9437),
.A2(n_6308),
.B1(n_6309),
.B2(n_6306),
.Y(n_10001)
);

INVx8_ASAP7_75t_L g10002 ( 
.A(n_9367),
.Y(n_10002)
);

AOI22xp5_ASAP7_75t_L g10003 ( 
.A1(n_9818),
.A2(n_9733),
.B1(n_9672),
.B2(n_9313),
.Y(n_10003)
);

NOR2xp33_ASAP7_75t_L g10004 ( 
.A(n_9432),
.B(n_6312),
.Y(n_10004)
);

AND2x2_ASAP7_75t_L g10005 ( 
.A(n_9423),
.B(n_9374),
.Y(n_10005)
);

NAND2xp5_ASAP7_75t_L g10006 ( 
.A(n_9548),
.B(n_6245),
.Y(n_10006)
);

INVx1_ASAP7_75t_L g10007 ( 
.A(n_9598),
.Y(n_10007)
);

NAND2xp5_ASAP7_75t_L g10008 ( 
.A(n_9600),
.B(n_6246),
.Y(n_10008)
);

AOI22xp33_ASAP7_75t_L g10009 ( 
.A1(n_9737),
.A2(n_6255),
.B1(n_6256),
.B2(n_6252),
.Y(n_10009)
);

NAND2xp5_ASAP7_75t_L g10010 ( 
.A(n_9613),
.B(n_6257),
.Y(n_10010)
);

NAND2xp5_ASAP7_75t_L g10011 ( 
.A(n_9614),
.B(n_6258),
.Y(n_10011)
);

NAND2xp5_ASAP7_75t_L g10012 ( 
.A(n_9615),
.B(n_6259),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_9616),
.Y(n_10013)
);

AOI22xp5_ASAP7_75t_L g10014 ( 
.A1(n_9313),
.A2(n_6314),
.B1(n_6316),
.B2(n_6313),
.Y(n_10014)
);

INVx1_ASAP7_75t_L g10015 ( 
.A(n_9618),
.Y(n_10015)
);

NOR2xp33_ASAP7_75t_L g10016 ( 
.A(n_9635),
.B(n_6317),
.Y(n_10016)
);

NAND2xp5_ASAP7_75t_L g10017 ( 
.A(n_9623),
.B(n_6262),
.Y(n_10017)
);

AND2x4_ASAP7_75t_L g10018 ( 
.A(n_9472),
.B(n_6263),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_9625),
.Y(n_10019)
);

AO221x1_ASAP7_75t_L g10020 ( 
.A1(n_9776),
.A2(n_9414),
.B1(n_9772),
.B2(n_9797),
.C(n_9784),
.Y(n_10020)
);

NAND2xp5_ASAP7_75t_SL g10021 ( 
.A(n_9522),
.B(n_6323),
.Y(n_10021)
);

NAND2xp5_ASAP7_75t_L g10022 ( 
.A(n_9631),
.B(n_6266),
.Y(n_10022)
);

O2A1O1Ixp5_ASAP7_75t_L g10023 ( 
.A1(n_9716),
.A2(n_6269),
.B(n_6272),
.C(n_6267),
.Y(n_10023)
);

AOI22xp33_ASAP7_75t_L g10024 ( 
.A1(n_9328),
.A2(n_6280),
.B1(n_6290),
.B2(n_6278),
.Y(n_10024)
);

OR2x6_ASAP7_75t_SL g10025 ( 
.A(n_9393),
.B(n_6326),
.Y(n_10025)
);

NAND2xp5_ASAP7_75t_L g10026 ( 
.A(n_9643),
.B(n_6292),
.Y(n_10026)
);

INVx2_ASAP7_75t_L g10027 ( 
.A(n_9646),
.Y(n_10027)
);

INVx2_ASAP7_75t_L g10028 ( 
.A(n_9652),
.Y(n_10028)
);

NOR2xp33_ASAP7_75t_L g10029 ( 
.A(n_9329),
.B(n_6328),
.Y(n_10029)
);

O2A1O1Ixp33_ASAP7_75t_L g10030 ( 
.A1(n_9354),
.A2(n_6299),
.B(n_6303),
.C(n_6296),
.Y(n_10030)
);

NOR2xp33_ASAP7_75t_L g10031 ( 
.A(n_9655),
.B(n_6333),
.Y(n_10031)
);

NAND3xp33_ASAP7_75t_L g10032 ( 
.A(n_9481),
.B(n_9587),
.C(n_9433),
.Y(n_10032)
);

AOI22xp5_ASAP7_75t_L g10033 ( 
.A1(n_9346),
.A2(n_6335),
.B1(n_6337),
.B2(n_6334),
.Y(n_10033)
);

INVx1_ASAP7_75t_L g10034 ( 
.A(n_9671),
.Y(n_10034)
);

NAND2x1p5_ASAP7_75t_L g10035 ( 
.A(n_9345),
.B(n_6304),
.Y(n_10035)
);

NAND2xp5_ASAP7_75t_L g10036 ( 
.A(n_9389),
.B(n_6315),
.Y(n_10036)
);

AOI22xp5_ASAP7_75t_L g10037 ( 
.A1(n_9328),
.A2(n_6346),
.B1(n_6347),
.B2(n_6341),
.Y(n_10037)
);

INVx1_ASAP7_75t_L g10038 ( 
.A(n_9556),
.Y(n_10038)
);

NAND2xp5_ASAP7_75t_L g10039 ( 
.A(n_9391),
.B(n_6324),
.Y(n_10039)
);

INVx1_ASAP7_75t_L g10040 ( 
.A(n_9326),
.Y(n_10040)
);

OR2x2_ASAP7_75t_L g10041 ( 
.A(n_9409),
.B(n_6348),
.Y(n_10041)
);

INVx1_ASAP7_75t_L g10042 ( 
.A(n_9344),
.Y(n_10042)
);

INVx1_ASAP7_75t_L g10043 ( 
.A(n_9352),
.Y(n_10043)
);

NAND2xp5_ASAP7_75t_L g10044 ( 
.A(n_9419),
.B(n_6327),
.Y(n_10044)
);

NAND2xp5_ASAP7_75t_SL g10045 ( 
.A(n_9522),
.B(n_6349),
.Y(n_10045)
);

INVx2_ASAP7_75t_L g10046 ( 
.A(n_9361),
.Y(n_10046)
);

NAND2xp5_ASAP7_75t_L g10047 ( 
.A(n_9434),
.B(n_6329),
.Y(n_10047)
);

NOR2xp67_ASAP7_75t_SL g10048 ( 
.A(n_9335),
.B(n_6351),
.Y(n_10048)
);

NAND2xp5_ASAP7_75t_L g10049 ( 
.A(n_9436),
.B(n_9440),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_9564),
.Y(n_10050)
);

NOR2xp33_ASAP7_75t_L g10051 ( 
.A(n_9340),
.B(n_6353),
.Y(n_10051)
);

INVx2_ASAP7_75t_SL g10052 ( 
.A(n_9397),
.Y(n_10052)
);

NAND2xp5_ASAP7_75t_L g10053 ( 
.A(n_9441),
.B(n_6332),
.Y(n_10053)
);

BUFx4f_ASAP7_75t_L g10054 ( 
.A(n_9397),
.Y(n_10054)
);

NOR2xp33_ASAP7_75t_L g10055 ( 
.A(n_9369),
.B(n_6354),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_SL g10056 ( 
.A(n_9416),
.B(n_6356),
.Y(n_10056)
);

NAND2xp5_ASAP7_75t_L g10057 ( 
.A(n_9462),
.B(n_9467),
.Y(n_10057)
);

NAND2xp5_ASAP7_75t_L g10058 ( 
.A(n_9476),
.B(n_6336),
.Y(n_10058)
);

NAND2xp5_ASAP7_75t_L g10059 ( 
.A(n_9485),
.B(n_6339),
.Y(n_10059)
);

NAND2xp5_ASAP7_75t_L g10060 ( 
.A(n_9493),
.B(n_6340),
.Y(n_10060)
);

BUFx3_ASAP7_75t_L g10061 ( 
.A(n_9418),
.Y(n_10061)
);

NAND2xp5_ASAP7_75t_L g10062 ( 
.A(n_9499),
.B(n_6342),
.Y(n_10062)
);

INVx2_ASAP7_75t_L g10063 ( 
.A(n_9504),
.Y(n_10063)
);

INVx2_ASAP7_75t_L g10064 ( 
.A(n_9508),
.Y(n_10064)
);

OR2x6_ASAP7_75t_L g10065 ( 
.A(n_9337),
.B(n_9661),
.Y(n_10065)
);

A2O1A1Ixp33_ASAP7_75t_L g10066 ( 
.A1(n_9382),
.A2(n_6344),
.B(n_6352),
.C(n_6343),
.Y(n_10066)
);

NOR2xp33_ASAP7_75t_L g10067 ( 
.A(n_9422),
.B(n_6358),
.Y(n_10067)
);

NAND2xp5_ASAP7_75t_SL g10068 ( 
.A(n_9483),
.B(n_6363),
.Y(n_10068)
);

AOI22xp33_ASAP7_75t_L g10069 ( 
.A1(n_9330),
.A2(n_9338),
.B1(n_9347),
.B2(n_9721),
.Y(n_10069)
);

NAND2xp5_ASAP7_75t_L g10070 ( 
.A(n_9509),
.B(n_6355),
.Y(n_10070)
);

INVx1_ASAP7_75t_L g10071 ( 
.A(n_9517),
.Y(n_10071)
);

AND2x2_ASAP7_75t_L g10072 ( 
.A(n_9378),
.B(n_9405),
.Y(n_10072)
);

INVx2_ASAP7_75t_L g10073 ( 
.A(n_9519),
.Y(n_10073)
);

NOR2xp33_ASAP7_75t_L g10074 ( 
.A(n_9394),
.B(n_6367),
.Y(n_10074)
);

OR2x2_ASAP7_75t_L g10075 ( 
.A(n_9611),
.B(n_6368),
.Y(n_10075)
);

INVx2_ASAP7_75t_SL g10076 ( 
.A(n_9430),
.Y(n_10076)
);

INVx1_ASAP7_75t_L g10077 ( 
.A(n_9787),
.Y(n_10077)
);

INVx2_ASAP7_75t_L g10078 ( 
.A(n_9591),
.Y(n_10078)
);

INVx2_ASAP7_75t_SL g10079 ( 
.A(n_9460),
.Y(n_10079)
);

INVxp67_ASAP7_75t_L g10080 ( 
.A(n_9633),
.Y(n_10080)
);

NAND2xp5_ASAP7_75t_L g10081 ( 
.A(n_9330),
.B(n_6364),
.Y(n_10081)
);

INVx2_ASAP7_75t_L g10082 ( 
.A(n_9599),
.Y(n_10082)
);

NAND2xp5_ASAP7_75t_L g10083 ( 
.A(n_9338),
.B(n_6366),
.Y(n_10083)
);

NAND2xp5_ASAP7_75t_L g10084 ( 
.A(n_9347),
.B(n_6369),
.Y(n_10084)
);

NAND2xp5_ASAP7_75t_L g10085 ( 
.A(n_9659),
.B(n_6370),
.Y(n_10085)
);

OAI22xp33_ASAP7_75t_L g10086 ( 
.A1(n_9417),
.A2(n_6375),
.B1(n_6376),
.B2(n_6371),
.Y(n_10086)
);

INVx1_ASAP7_75t_L g10087 ( 
.A(n_9791),
.Y(n_10087)
);

OAI22xp5_ASAP7_75t_L g10088 ( 
.A1(n_9453),
.A2(n_6377),
.B1(n_6379),
.B2(n_6378),
.Y(n_10088)
);

NAND2xp5_ASAP7_75t_SL g10089 ( 
.A(n_9483),
.B(n_6384),
.Y(n_10089)
);

NAND2xp5_ASAP7_75t_SL g10090 ( 
.A(n_9784),
.B(n_9797),
.Y(n_10090)
);

AOI22xp5_ASAP7_75t_L g10091 ( 
.A1(n_9730),
.A2(n_6388),
.B1(n_6389),
.B2(n_6387),
.Y(n_10091)
);

NOR2xp33_ASAP7_75t_L g10092 ( 
.A(n_9665),
.B(n_6390),
.Y(n_10092)
);

INVx2_ASAP7_75t_SL g10093 ( 
.A(n_9506),
.Y(n_10093)
);

AOI22xp5_ASAP7_75t_L g10094 ( 
.A1(n_9667),
.A2(n_6393),
.B1(n_6395),
.B2(n_6391),
.Y(n_10094)
);

NOR3xp33_ASAP7_75t_L g10095 ( 
.A(n_9804),
.B(n_6385),
.C(n_6374),
.Y(n_10095)
);

NAND2xp5_ASAP7_75t_SL g10096 ( 
.A(n_9707),
.B(n_6402),
.Y(n_10096)
);

NAND2xp5_ASAP7_75t_L g10097 ( 
.A(n_9320),
.B(n_6386),
.Y(n_10097)
);

OAI22xp5_ASAP7_75t_L g10098 ( 
.A1(n_9612),
.A2(n_6406),
.B1(n_6408),
.B2(n_6405),
.Y(n_10098)
);

NAND2xp5_ASAP7_75t_SL g10099 ( 
.A(n_9712),
.B(n_6411),
.Y(n_10099)
);

NAND2xp5_ASAP7_75t_L g10100 ( 
.A(n_9759),
.B(n_6392),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_9683),
.Y(n_10101)
);

NAND3xp33_ASAP7_75t_L g10102 ( 
.A(n_9350),
.B(n_6414),
.C(n_6412),
.Y(n_10102)
);

NOR2xp33_ASAP7_75t_L g10103 ( 
.A(n_9552),
.B(n_6416),
.Y(n_10103)
);

NOR2xp33_ASAP7_75t_L g10104 ( 
.A(n_9577),
.B(n_6420),
.Y(n_10104)
);

NAND2xp5_ASAP7_75t_SL g10105 ( 
.A(n_9713),
.B(n_6423),
.Y(n_10105)
);

NAND2xp5_ASAP7_75t_L g10106 ( 
.A(n_9783),
.B(n_6398),
.Y(n_10106)
);

NAND2xp33_ASAP7_75t_L g10107 ( 
.A(n_9569),
.B(n_6426),
.Y(n_10107)
);

NOR2xp33_ASAP7_75t_L g10108 ( 
.A(n_9609),
.B(n_6427),
.Y(n_10108)
);

INVx5_ASAP7_75t_L g10109 ( 
.A(n_9561),
.Y(n_10109)
);

NAND2xp33_ASAP7_75t_L g10110 ( 
.A(n_9569),
.B(n_6429),
.Y(n_10110)
);

INVx1_ASAP7_75t_L g10111 ( 
.A(n_9685),
.Y(n_10111)
);

BUFx6f_ASAP7_75t_L g10112 ( 
.A(n_9365),
.Y(n_10112)
);

INVx2_ASAP7_75t_L g10113 ( 
.A(n_9601),
.Y(n_10113)
);

OR2x6_ASAP7_75t_L g10114 ( 
.A(n_9331),
.B(n_6399),
.Y(n_10114)
);

NOR2xp33_ASAP7_75t_L g10115 ( 
.A(n_9794),
.B(n_6430),
.Y(n_10115)
);

NAND2xp5_ASAP7_75t_L g10116 ( 
.A(n_9687),
.B(n_6400),
.Y(n_10116)
);

NAND2xp5_ASAP7_75t_L g10117 ( 
.A(n_9689),
.B(n_6413),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9720),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_9722),
.Y(n_10119)
);

INVx2_ASAP7_75t_L g10120 ( 
.A(n_9606),
.Y(n_10120)
);

NAND2xp5_ASAP7_75t_L g10121 ( 
.A(n_9725),
.B(n_6415),
.Y(n_10121)
);

O2A1O1Ixp33_ASAP7_75t_L g10122 ( 
.A1(n_9639),
.A2(n_6421),
.B(n_6425),
.C(n_6419),
.Y(n_10122)
);

NAND2xp5_ASAP7_75t_L g10123 ( 
.A(n_9732),
.B(n_6428),
.Y(n_10123)
);

AOI22xp5_ASAP7_75t_L g10124 ( 
.A1(n_9667),
.A2(n_9421),
.B1(n_9387),
.B2(n_9741),
.Y(n_10124)
);

NAND2xp5_ASAP7_75t_L g10125 ( 
.A(n_9739),
.B(n_6437),
.Y(n_10125)
);

OAI21xp5_ASAP7_75t_L g10126 ( 
.A1(n_9817),
.A2(n_6439),
.B(n_6438),
.Y(n_10126)
);

INVx3_ASAP7_75t_L g10127 ( 
.A(n_9648),
.Y(n_10127)
);

AND2x2_ASAP7_75t_L g10128 ( 
.A(n_9765),
.B(n_6433),
.Y(n_10128)
);

INVx2_ASAP7_75t_L g10129 ( 
.A(n_9608),
.Y(n_10129)
);

NAND2xp5_ASAP7_75t_L g10130 ( 
.A(n_9747),
.B(n_6441),
.Y(n_10130)
);

OAI22xp5_ASAP7_75t_L g10131 ( 
.A1(n_9809),
.A2(n_6442),
.B1(n_6445),
.B2(n_6440),
.Y(n_10131)
);

INVx1_ASAP7_75t_L g10132 ( 
.A(n_9749),
.Y(n_10132)
);

NOR2xp33_ASAP7_75t_L g10133 ( 
.A(n_9781),
.B(n_6446),
.Y(n_10133)
);

NAND2xp5_ASAP7_75t_L g10134 ( 
.A(n_9755),
.B(n_6443),
.Y(n_10134)
);

INVx2_ASAP7_75t_L g10135 ( 
.A(n_9617),
.Y(n_10135)
);

INVx3_ASAP7_75t_L g10136 ( 
.A(n_9385),
.Y(n_10136)
);

NAND2xp5_ASAP7_75t_L g10137 ( 
.A(n_9761),
.B(n_6448),
.Y(n_10137)
);

INVx1_ASAP7_75t_L g10138 ( 
.A(n_9786),
.Y(n_10138)
);

INVx1_ASAP7_75t_L g10139 ( 
.A(n_9627),
.Y(n_10139)
);

NAND2xp5_ASAP7_75t_L g10140 ( 
.A(n_9629),
.B(n_6451),
.Y(n_10140)
);

NAND2xp5_ASAP7_75t_L g10141 ( 
.A(n_9650),
.B(n_6461),
.Y(n_10141)
);

NAND2xp5_ASAP7_75t_SL g10142 ( 
.A(n_9390),
.B(n_6447),
.Y(n_10142)
);

INVx3_ASAP7_75t_L g10143 ( 
.A(n_9398),
.Y(n_10143)
);

NAND2xp5_ASAP7_75t_SL g10144 ( 
.A(n_9503),
.B(n_6449),
.Y(n_10144)
);

INVx2_ASAP7_75t_L g10145 ( 
.A(n_9656),
.Y(n_10145)
);

NOR2xp33_ASAP7_75t_L g10146 ( 
.A(n_9489),
.B(n_9549),
.Y(n_10146)
);

NAND2xp5_ASAP7_75t_SL g10147 ( 
.A(n_9734),
.B(n_6452),
.Y(n_10147)
);

NOR2xp33_ASAP7_75t_L g10148 ( 
.A(n_9595),
.B(n_6453),
.Y(n_10148)
);

INVxp33_ASAP7_75t_L g10149 ( 
.A(n_9742),
.Y(n_10149)
);

NAND2xp5_ASAP7_75t_L g10150 ( 
.A(n_9682),
.B(n_6479),
.Y(n_10150)
);

INVx2_ASAP7_75t_SL g10151 ( 
.A(n_9506),
.Y(n_10151)
);

NAND2xp5_ASAP7_75t_SL g10152 ( 
.A(n_9734),
.B(n_6454),
.Y(n_10152)
);

NAND2xp5_ASAP7_75t_L g10153 ( 
.A(n_9703),
.B(n_6484),
.Y(n_10153)
);

NOR2xp33_ASAP7_75t_L g10154 ( 
.A(n_9469),
.B(n_6455),
.Y(n_10154)
);

NAND2xp5_ASAP7_75t_SL g10155 ( 
.A(n_9775),
.B(n_6456),
.Y(n_10155)
);

NOR2xp33_ASAP7_75t_L g10156 ( 
.A(n_9474),
.B(n_6459),
.Y(n_10156)
);

NOR3xp33_ASAP7_75t_L g10157 ( 
.A(n_9371),
.B(n_6495),
.C(n_6490),
.Y(n_10157)
);

NAND2xp5_ASAP7_75t_SL g10158 ( 
.A(n_9775),
.B(n_6463),
.Y(n_10158)
);

INVx2_ASAP7_75t_L g10159 ( 
.A(n_9718),
.Y(n_10159)
);

BUFx6f_ASAP7_75t_L g10160 ( 
.A(n_9554),
.Y(n_10160)
);

NOR2xp33_ASAP7_75t_L g10161 ( 
.A(n_9511),
.B(n_6464),
.Y(n_10161)
);

NAND2xp5_ASAP7_75t_SL g10162 ( 
.A(n_9554),
.B(n_9628),
.Y(n_10162)
);

INVx3_ASAP7_75t_L g10163 ( 
.A(n_9426),
.Y(n_10163)
);

NAND2xp5_ASAP7_75t_L g10164 ( 
.A(n_9719),
.B(n_6498),
.Y(n_10164)
);

INVx2_ASAP7_75t_L g10165 ( 
.A(n_9735),
.Y(n_10165)
);

NOR2xp33_ASAP7_75t_L g10166 ( 
.A(n_9515),
.B(n_6465),
.Y(n_10166)
);

NAND2xp5_ASAP7_75t_L g10167 ( 
.A(n_9736),
.B(n_6505),
.Y(n_10167)
);

INVx2_ASAP7_75t_L g10168 ( 
.A(n_9740),
.Y(n_10168)
);

INVx1_ASAP7_75t_L g10169 ( 
.A(n_9743),
.Y(n_10169)
);

INVx1_ASAP7_75t_L g10170 ( 
.A(n_9744),
.Y(n_10170)
);

INVx2_ASAP7_75t_L g10171 ( 
.A(n_9771),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_9777),
.Y(n_10172)
);

INVx2_ASAP7_75t_SL g10173 ( 
.A(n_9628),
.Y(n_10173)
);

NAND2xp5_ASAP7_75t_SL g10174 ( 
.A(n_9756),
.B(n_9370),
.Y(n_10174)
);

INVx2_ASAP7_75t_L g10175 ( 
.A(n_9803),
.Y(n_10175)
);

NAND2xp5_ASAP7_75t_L g10176 ( 
.A(n_9551),
.B(n_9708),
.Y(n_10176)
);

NAND2xp5_ASAP7_75t_L g10177 ( 
.A(n_9709),
.B(n_6520),
.Y(n_10177)
);

INVxp67_ASAP7_75t_L g10178 ( 
.A(n_9770),
.Y(n_10178)
);

INVx1_ASAP7_75t_L g10179 ( 
.A(n_9792),
.Y(n_10179)
);

NAND2x1_ASAP7_75t_L g10180 ( 
.A(n_9793),
.B(n_6524),
.Y(n_10180)
);

INVxp67_ASAP7_75t_SL g10181 ( 
.A(n_9379),
.Y(n_10181)
);

NOR2xp33_ASAP7_75t_L g10182 ( 
.A(n_9536),
.B(n_6470),
.Y(n_10182)
);

INVx2_ASAP7_75t_L g10183 ( 
.A(n_9796),
.Y(n_10183)
);

AOI22xp33_ASAP7_75t_L g10184 ( 
.A1(n_9660),
.A2(n_9802),
.B1(n_9473),
.B2(n_9805),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_SL g10185 ( 
.A(n_9651),
.B(n_6472),
.Y(n_10185)
);

NAND2xp5_ASAP7_75t_SL g10186 ( 
.A(n_9658),
.B(n_6473),
.Y(n_10186)
);

INVx1_ASAP7_75t_L g10187 ( 
.A(n_9798),
.Y(n_10187)
);

BUFx6f_ASAP7_75t_L g10188 ( 
.A(n_9636),
.Y(n_10188)
);

NOR2xp33_ASAP7_75t_L g10189 ( 
.A(n_9543),
.B(n_6474),
.Y(n_10189)
);

INVx1_ASAP7_75t_L g10190 ( 
.A(n_9799),
.Y(n_10190)
);

NOR3xp33_ASAP7_75t_L g10191 ( 
.A(n_9663),
.B(n_6544),
.C(n_6542),
.Y(n_10191)
);

NOR2xp33_ASAP7_75t_L g10192 ( 
.A(n_9550),
.B(n_6475),
.Y(n_10192)
);

BUFx5_ASAP7_75t_L g10193 ( 
.A(n_9823),
.Y(n_10193)
);

INVx2_ASAP7_75t_L g10194 ( 
.A(n_9800),
.Y(n_10194)
);

CKINVDCx11_ASAP7_75t_R g10195 ( 
.A(n_9468),
.Y(n_10195)
);

INVx2_ASAP7_75t_L g10196 ( 
.A(n_9807),
.Y(n_10196)
);

INVx2_ASAP7_75t_SL g10197 ( 
.A(n_9442),
.Y(n_10197)
);

NAND2xp5_ASAP7_75t_L g10198 ( 
.A(n_9748),
.B(n_6570),
.Y(n_10198)
);

AOI22xp5_ASAP7_75t_SL g10199 ( 
.A1(n_9814),
.A2(n_6477),
.B1(n_6481),
.B2(n_6476),
.Y(n_10199)
);

AND2x2_ASAP7_75t_L g10200 ( 
.A(n_9529),
.B(n_6485),
.Y(n_10200)
);

INVx1_ASAP7_75t_L g10201 ( 
.A(n_9808),
.Y(n_10201)
);

AOI221xp5_ASAP7_75t_L g10202 ( 
.A1(n_9821),
.A2(n_6590),
.B1(n_6592),
.B2(n_6581),
.C(n_6576),
.Y(n_10202)
);

INVx2_ASAP7_75t_SL g10203 ( 
.A(n_9464),
.Y(n_10203)
);

NOR2xp33_ASAP7_75t_L g10204 ( 
.A(n_9695),
.B(n_6486),
.Y(n_10204)
);

NAND2xp5_ASAP7_75t_L g10205 ( 
.A(n_9751),
.B(n_9752),
.Y(n_10205)
);

NAND2xp33_ASAP7_75t_L g10206 ( 
.A(n_9649),
.B(n_6487),
.Y(n_10206)
);

INVx1_ASAP7_75t_L g10207 ( 
.A(n_9697),
.Y(n_10207)
);

NOR2xp33_ASAP7_75t_L g10208 ( 
.A(n_9431),
.B(n_6488),
.Y(n_10208)
);

NAND2xp5_ASAP7_75t_SL g10209 ( 
.A(n_9636),
.B(n_6492),
.Y(n_10209)
);

INVx2_ASAP7_75t_L g10210 ( 
.A(n_9801),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_9478),
.Y(n_10211)
);

NAND2xp5_ASAP7_75t_SL g10212 ( 
.A(n_9757),
.B(n_6499),
.Y(n_10212)
);

NOR2xp33_ASAP7_75t_L g10213 ( 
.A(n_9461),
.B(n_6500),
.Y(n_10213)
);

BUFx6f_ASAP7_75t_SL g10214 ( 
.A(n_9372),
.Y(n_10214)
);

NOR3xp33_ASAP7_75t_L g10215 ( 
.A(n_9670),
.B(n_6595),
.C(n_6593),
.Y(n_10215)
);

INVx2_ASAP7_75t_L g10216 ( 
.A(n_9662),
.Y(n_10216)
);

NAND2xp5_ASAP7_75t_L g10217 ( 
.A(n_9753),
.B(n_6598),
.Y(n_10217)
);

INVx1_ASAP7_75t_L g10218 ( 
.A(n_9677),
.Y(n_10218)
);

OAI22xp33_ASAP7_75t_L g10219 ( 
.A1(n_9704),
.A2(n_6502),
.B1(n_6504),
.B2(n_6501),
.Y(n_10219)
);

INVx1_ASAP7_75t_L g10220 ( 
.A(n_9678),
.Y(n_10220)
);

AND2x4_ASAP7_75t_L g10221 ( 
.A(n_9702),
.B(n_6609),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_9746),
.Y(n_10222)
);

NOR2xp33_ASAP7_75t_L g10223 ( 
.A(n_9446),
.B(n_6507),
.Y(n_10223)
);

INVx2_ASAP7_75t_L g10224 ( 
.A(n_9698),
.Y(n_10224)
);

NAND2xp5_ASAP7_75t_L g10225 ( 
.A(n_9754),
.B(n_6620),
.Y(n_10225)
);

NAND2xp5_ASAP7_75t_SL g10226 ( 
.A(n_9673),
.B(n_6510),
.Y(n_10226)
);

NAND2xp5_ASAP7_75t_L g10227 ( 
.A(n_9782),
.B(n_9649),
.Y(n_10227)
);

NOR2xp33_ASAP7_75t_L g10228 ( 
.A(n_9448),
.B(n_9424),
.Y(n_10228)
);

INVx2_ASAP7_75t_SL g10229 ( 
.A(n_9327),
.Y(n_10229)
);

INVx2_ASAP7_75t_L g10230 ( 
.A(n_9726),
.Y(n_10230)
);

INVx2_ASAP7_75t_L g10231 ( 
.A(n_9729),
.Y(n_10231)
);

OAI22xp5_ASAP7_75t_SL g10232 ( 
.A1(n_9684),
.A2(n_6512),
.B1(n_6514),
.B2(n_6511),
.Y(n_10232)
);

INVx1_ASAP7_75t_L g10233 ( 
.A(n_9763),
.Y(n_10233)
);

INVxp67_ASAP7_75t_L g10234 ( 
.A(n_9533),
.Y(n_10234)
);

NAND2xp5_ASAP7_75t_L g10235 ( 
.A(n_9745),
.B(n_6516),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9760),
.Y(n_10236)
);

INVx2_ASAP7_75t_L g10237 ( 
.A(n_9767),
.Y(n_10237)
);

OAI22xp5_ASAP7_75t_L g10238 ( 
.A1(n_9700),
.A2(n_6518),
.B1(n_6519),
.B2(n_6517),
.Y(n_10238)
);

AOI22xp5_ASAP7_75t_L g10239 ( 
.A1(n_9387),
.A2(n_6530),
.B1(n_6531),
.B2(n_6523),
.Y(n_10239)
);

NAND3xp33_ASAP7_75t_L g10240 ( 
.A(n_9653),
.B(n_6541),
.C(n_6538),
.Y(n_10240)
);

NAND2xp5_ASAP7_75t_L g10241 ( 
.A(n_9789),
.B(n_6543),
.Y(n_10241)
);

INVx2_ASAP7_75t_L g10242 ( 
.A(n_9773),
.Y(n_10242)
);

BUFx8_ASAP7_75t_L g10243 ( 
.A(n_9778),
.Y(n_10243)
);

INVx2_ASAP7_75t_L g10244 ( 
.A(n_9738),
.Y(n_10244)
);

INVx1_ASAP7_75t_L g10245 ( 
.A(n_9471),
.Y(n_10245)
);

INVx1_ASAP7_75t_L g10246 ( 
.A(n_9539),
.Y(n_10246)
);

NOR2xp33_ASAP7_75t_L g10247 ( 
.A(n_9642),
.B(n_9750),
.Y(n_10247)
);

AOI22xp5_ASAP7_75t_L g10248 ( 
.A1(n_9427),
.A2(n_9588),
.B1(n_9558),
.B2(n_9449),
.Y(n_10248)
);

INVx1_ASAP7_75t_L g10249 ( 
.A(n_9578),
.Y(n_10249)
);

NOR2xp67_ASAP7_75t_L g10250 ( 
.A(n_9438),
.B(n_4588),
.Y(n_10250)
);

INVx2_ASAP7_75t_L g10251 ( 
.A(n_9605),
.Y(n_10251)
);

NAND2xp5_ASAP7_75t_L g10252 ( 
.A(n_9668),
.B(n_9669),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_9806),
.Y(n_10253)
);

NAND2xp5_ASAP7_75t_SL g10254 ( 
.A(n_9764),
.B(n_6545),
.Y(n_10254)
);

INVx1_ASAP7_75t_L g10255 ( 
.A(n_9812),
.Y(n_10255)
);

INVx2_ASAP7_75t_L g10256 ( 
.A(n_9512),
.Y(n_10256)
);

XOR2xp5_ASAP7_75t_L g10257 ( 
.A(n_9701),
.B(n_4590),
.Y(n_10257)
);

NOR2xp33_ASAP7_75t_L g10258 ( 
.A(n_9758),
.B(n_6546),
.Y(n_10258)
);

BUFx3_ASAP7_75t_L g10259 ( 
.A(n_9445),
.Y(n_10259)
);

AND2x2_ASAP7_75t_L g10260 ( 
.A(n_9675),
.B(n_6550),
.Y(n_10260)
);

INVx3_ASAP7_75t_L g10261 ( 
.A(n_9572),
.Y(n_10261)
);

NAND2xp5_ASAP7_75t_L g10262 ( 
.A(n_9699),
.B(n_6554),
.Y(n_10262)
);

AOI22xp5_ASAP7_75t_L g10263 ( 
.A1(n_9558),
.A2(n_9588),
.B1(n_9455),
.B2(n_9691),
.Y(n_10263)
);

NAND3xp33_ASAP7_75t_L g10264 ( 
.A(n_9657),
.B(n_6562),
.C(n_6558),
.Y(n_10264)
);

NOR2xp33_ASAP7_75t_L g10265 ( 
.A(n_9579),
.B(n_6564),
.Y(n_10265)
);

NAND2xp5_ASAP7_75t_SL g10266 ( 
.A(n_9538),
.B(n_6565),
.Y(n_10266)
);

NAND2xp5_ASAP7_75t_L g10267 ( 
.A(n_9428),
.B(n_6567),
.Y(n_10267)
);

NAND2xp5_ASAP7_75t_SL g10268 ( 
.A(n_9593),
.B(n_6568),
.Y(n_10268)
);

INVx8_ASAP7_75t_L g10269 ( 
.A(n_9607),
.Y(n_10269)
);

OR2x2_ASAP7_75t_L g10270 ( 
.A(n_9516),
.B(n_6569),
.Y(n_10270)
);

INVx1_ASAP7_75t_L g10271 ( 
.A(n_9524),
.Y(n_10271)
);

INVx2_ASAP7_75t_SL g10272 ( 
.A(n_9547),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9411),
.Y(n_10273)
);

INVx1_ASAP7_75t_L g10274 ( 
.A(n_9415),
.Y(n_10274)
);

O2A1O1Ixp5_ASAP7_75t_L g10275 ( 
.A1(n_9714),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_10275)
);

INVxp67_ASAP7_75t_L g10276 ( 
.A(n_9604),
.Y(n_10276)
);

INVx1_ASAP7_75t_L g10277 ( 
.A(n_9795),
.Y(n_10277)
);

NOR2xp33_ASAP7_75t_L g10278 ( 
.A(n_9619),
.B(n_6571),
.Y(n_10278)
);

NAND2xp33_ASAP7_75t_L g10279 ( 
.A(n_9428),
.B(n_6572),
.Y(n_10279)
);

NAND2xp5_ASAP7_75t_L g10280 ( 
.A(n_9406),
.B(n_6575),
.Y(n_10280)
);

INVx2_ASAP7_75t_L g10281 ( 
.A(n_9526),
.Y(n_10281)
);

NOR2xp33_ASAP7_75t_L g10282 ( 
.A(n_9630),
.B(n_6578),
.Y(n_10282)
);

NAND2xp5_ASAP7_75t_L g10283 ( 
.A(n_9406),
.B(n_6580),
.Y(n_10283)
);

AOI22xp5_ASAP7_75t_L g10284 ( 
.A1(n_9465),
.A2(n_6584),
.B1(n_6585),
.B2(n_6583),
.Y(n_10284)
);

NAND2xp5_ASAP7_75t_L g10285 ( 
.A(n_9666),
.B(n_6586),
.Y(n_10285)
);

INVx3_ASAP7_75t_L g10286 ( 
.A(n_9532),
.Y(n_10286)
);

NAND2xp5_ASAP7_75t_L g10287 ( 
.A(n_9546),
.B(n_6587),
.Y(n_10287)
);

NAND2x1_ASAP7_75t_L g10288 ( 
.A(n_9570),
.B(n_4591),
.Y(n_10288)
);

INVxp33_ASAP7_75t_L g10289 ( 
.A(n_9620),
.Y(n_10289)
);

NAND2xp5_ASAP7_75t_L g10290 ( 
.A(n_9581),
.B(n_6588),
.Y(n_10290)
);

OAI21xp5_ASAP7_75t_L g10291 ( 
.A1(n_9690),
.A2(n_6589),
.B(n_4593),
.Y(n_10291)
);

AOI21xp5_ASAP7_75t_L g10292 ( 
.A1(n_9407),
.A2(n_4594),
.B(n_4592),
.Y(n_10292)
);

BUFx5_ASAP7_75t_L g10293 ( 
.A(n_9541),
.Y(n_10293)
);

INVx1_ASAP7_75t_L g10294 ( 
.A(n_9586),
.Y(n_10294)
);

NOR2xp33_ASAP7_75t_L g10295 ( 
.A(n_9723),
.B(n_8),
.Y(n_10295)
);

INVx3_ASAP7_75t_L g10296 ( 
.A(n_9514),
.Y(n_10296)
);

INVx2_ASAP7_75t_L g10297 ( 
.A(n_9822),
.Y(n_10297)
);

INVx2_ASAP7_75t_L g10298 ( 
.A(n_9779),
.Y(n_10298)
);

NAND2xp5_ASAP7_75t_L g10299 ( 
.A(n_9597),
.B(n_9),
.Y(n_10299)
);

NAND2xp5_ASAP7_75t_L g10300 ( 
.A(n_9686),
.B(n_10),
.Y(n_10300)
);

NAND2xp5_ASAP7_75t_L g10301 ( 
.A(n_9465),
.B(n_10),
.Y(n_10301)
);

INVx2_ASAP7_75t_SL g10302 ( 
.A(n_9384),
.Y(n_10302)
);

NAND2xp5_ASAP7_75t_L g10303 ( 
.A(n_9525),
.B(n_9537),
.Y(n_10303)
);

NAND2xp5_ASAP7_75t_L g10304 ( 
.A(n_9525),
.B(n_11),
.Y(n_10304)
);

NAND2xp5_ASAP7_75t_L g10305 ( 
.A(n_9537),
.B(n_11),
.Y(n_10305)
);

AND2x6_ASAP7_75t_L g10306 ( 
.A(n_9778),
.B(n_4596),
.Y(n_10306)
);

NAND2xp5_ASAP7_75t_L g10307 ( 
.A(n_9541),
.B(n_9540),
.Y(n_10307)
);

INVx1_ASAP7_75t_L g10308 ( 
.A(n_9501),
.Y(n_10308)
);

INVx3_ASAP7_75t_L g10309 ( 
.A(n_9429),
.Y(n_10309)
);

AND2x2_ASAP7_75t_L g10310 ( 
.A(n_9475),
.B(n_12),
.Y(n_10310)
);

NOR2xp33_ASAP7_75t_L g10311 ( 
.A(n_9815),
.B(n_12),
.Y(n_10311)
);

NAND2xp5_ASAP7_75t_L g10312 ( 
.A(n_9540),
.B(n_13),
.Y(n_10312)
);

OR2x6_ASAP7_75t_L g10313 ( 
.A(n_9603),
.B(n_4597),
.Y(n_10313)
);

NAND2xp5_ASAP7_75t_SL g10314 ( 
.A(n_9811),
.B(n_13),
.Y(n_10314)
);

NAND2xp5_ASAP7_75t_SL g10315 ( 
.A(n_9463),
.B(n_14),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_9429),
.Y(n_10316)
);

NOR2xp33_ASAP7_75t_L g10317 ( 
.A(n_9814),
.B(n_14),
.Y(n_10317)
);

NAND2xp5_ASAP7_75t_SL g10318 ( 
.A(n_9820),
.B(n_15),
.Y(n_10318)
);

INVx1_ASAP7_75t_SL g10319 ( 
.A(n_9435),
.Y(n_10319)
);

INVx1_ASAP7_75t_L g10320 ( 
.A(n_9435),
.Y(n_10320)
);

A2O1A1Ixp33_ASAP7_75t_L g10321 ( 
.A1(n_9626),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_10321)
);

INVx1_ASAP7_75t_L g10322 ( 
.A(n_9444),
.Y(n_10322)
);

NOR2xp33_ASAP7_75t_L g10323 ( 
.A(n_9820),
.B(n_16),
.Y(n_10323)
);

NAND2xp5_ASAP7_75t_L g10324 ( 
.A(n_9444),
.B(n_17),
.Y(n_10324)
);

NAND2xp5_ASAP7_75t_SL g10325 ( 
.A(n_9454),
.B(n_18),
.Y(n_10325)
);

INVx2_ASAP7_75t_L g10326 ( 
.A(n_9641),
.Y(n_10326)
);

NOR2xp33_ASAP7_75t_L g10327 ( 
.A(n_9454),
.B(n_19),
.Y(n_10327)
);

INVx2_ASAP7_75t_SL g10328 ( 
.A(n_9400),
.Y(n_10328)
);

NOR2xp33_ASAP7_75t_L g10329 ( 
.A(n_9343),
.B(n_19),
.Y(n_10329)
);

INVx2_ASAP7_75t_L g10330 ( 
.A(n_9317),
.Y(n_10330)
);

AOI21xp5_ASAP7_75t_L g10331 ( 
.A1(n_9388),
.A2(n_4600),
.B(n_4598),
.Y(n_10331)
);

NAND2xp5_ASAP7_75t_L g10332 ( 
.A(n_9343),
.B(n_20),
.Y(n_10332)
);

OAI21xp5_ASAP7_75t_L g10333 ( 
.A1(n_9316),
.A2(n_4603),
.B(n_4601),
.Y(n_10333)
);

A2O1A1Ixp33_ASAP7_75t_L g10334 ( 
.A1(n_9343),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_10334)
);

NAND2xp5_ASAP7_75t_SL g10335 ( 
.A(n_9343),
.B(n_22),
.Y(n_10335)
);

AND2x2_ASAP7_75t_L g10336 ( 
.A(n_9343),
.B(n_23),
.Y(n_10336)
);

NOR2xp33_ASAP7_75t_L g10337 ( 
.A(n_9343),
.B(n_23),
.Y(n_10337)
);

INVxp67_ASAP7_75t_L g10338 ( 
.A(n_9332),
.Y(n_10338)
);

INVx3_ASAP7_75t_L g10339 ( 
.A(n_9318),
.Y(n_10339)
);

NAND2xp5_ASAP7_75t_L g10340 ( 
.A(n_9343),
.B(n_24),
.Y(n_10340)
);

AND2x4_ASAP7_75t_L g10341 ( 
.A(n_9318),
.B(n_4604),
.Y(n_10341)
);

NAND2xp5_ASAP7_75t_SL g10342 ( 
.A(n_9343),
.B(n_24),
.Y(n_10342)
);

NOR2xp33_ASAP7_75t_L g10343 ( 
.A(n_9343),
.B(n_25),
.Y(n_10343)
);

AND2x4_ASAP7_75t_L g10344 ( 
.A(n_9873),
.B(n_9884),
.Y(n_10344)
);

INVx2_ASAP7_75t_L g10345 ( 
.A(n_9830),
.Y(n_10345)
);

OAI21xp5_ASAP7_75t_L g10346 ( 
.A1(n_9868),
.A2(n_25),
.B(n_26),
.Y(n_10346)
);

NOR2xp33_ASAP7_75t_L g10347 ( 
.A(n_9861),
.B(n_4607),
.Y(n_10347)
);

INVx2_ASAP7_75t_SL g10348 ( 
.A(n_10054),
.Y(n_10348)
);

NOR2xp33_ASAP7_75t_L g10349 ( 
.A(n_9827),
.B(n_4609),
.Y(n_10349)
);

INVx1_ASAP7_75t_L g10350 ( 
.A(n_9835),
.Y(n_10350)
);

INVx1_ASAP7_75t_L g10351 ( 
.A(n_9856),
.Y(n_10351)
);

BUFx3_ASAP7_75t_L g10352 ( 
.A(n_9886),
.Y(n_10352)
);

AND2x2_ASAP7_75t_L g10353 ( 
.A(n_10005),
.B(n_26),
.Y(n_10353)
);

INVx2_ASAP7_75t_L g10354 ( 
.A(n_9897),
.Y(n_10354)
);

INVxp67_ASAP7_75t_L g10355 ( 
.A(n_9870),
.Y(n_10355)
);

INVx2_ASAP7_75t_L g10356 ( 
.A(n_9899),
.Y(n_10356)
);

INVx2_ASAP7_75t_L g10357 ( 
.A(n_9909),
.Y(n_10357)
);

AND2x2_ASAP7_75t_L g10358 ( 
.A(n_10072),
.B(n_27),
.Y(n_10358)
);

INVx6_ASAP7_75t_L g10359 ( 
.A(n_10112),
.Y(n_10359)
);

NAND2xp5_ASAP7_75t_L g10360 ( 
.A(n_9834),
.B(n_9829),
.Y(n_10360)
);

NAND2x1p5_ASAP7_75t_L g10361 ( 
.A(n_10000),
.B(n_4610),
.Y(n_10361)
);

INVx1_ASAP7_75t_L g10362 ( 
.A(n_9913),
.Y(n_10362)
);

AND2x2_ASAP7_75t_L g10363 ( 
.A(n_10336),
.B(n_28),
.Y(n_10363)
);

AOI22xp5_ASAP7_75t_L g10364 ( 
.A1(n_9857),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_10364)
);

INVx1_ASAP7_75t_L g10365 ( 
.A(n_9928),
.Y(n_10365)
);

INVx2_ASAP7_75t_L g10366 ( 
.A(n_9956),
.Y(n_10366)
);

INVx1_ASAP7_75t_L g10367 ( 
.A(n_9960),
.Y(n_10367)
);

AND2x2_ASAP7_75t_L g10368 ( 
.A(n_10128),
.B(n_29),
.Y(n_10368)
);

BUFx3_ASAP7_75t_L g10369 ( 
.A(n_9886),
.Y(n_10369)
);

NAND2xp5_ASAP7_75t_L g10370 ( 
.A(n_9846),
.B(n_31),
.Y(n_10370)
);

AND2x2_ASAP7_75t_L g10371 ( 
.A(n_9952),
.B(n_32),
.Y(n_10371)
);

NOR2xp33_ASAP7_75t_L g10372 ( 
.A(n_9878),
.B(n_4611),
.Y(n_10372)
);

AND2x2_ASAP7_75t_L g10373 ( 
.A(n_9996),
.B(n_32),
.Y(n_10373)
);

NAND2xp5_ASAP7_75t_L g10374 ( 
.A(n_9894),
.B(n_33),
.Y(n_10374)
);

BUFx3_ASAP7_75t_L g10375 ( 
.A(n_9934),
.Y(n_10375)
);

INVx1_ASAP7_75t_SL g10376 ( 
.A(n_9935),
.Y(n_10376)
);

INVx2_ASAP7_75t_L g10377 ( 
.A(n_9962),
.Y(n_10377)
);

HB1xp67_ASAP7_75t_L g10378 ( 
.A(n_9940),
.Y(n_10378)
);

BUFx3_ASAP7_75t_L g10379 ( 
.A(n_9934),
.Y(n_10379)
);

INVx2_ASAP7_75t_L g10380 ( 
.A(n_9966),
.Y(n_10380)
);

AND2x2_ASAP7_75t_SL g10381 ( 
.A(n_10329),
.B(n_33),
.Y(n_10381)
);

AND2x2_ASAP7_75t_L g10382 ( 
.A(n_9923),
.B(n_34),
.Y(n_10382)
);

AND2x4_ASAP7_75t_L g10383 ( 
.A(n_9949),
.B(n_4613),
.Y(n_10383)
);

INVxp67_ASAP7_75t_SL g10384 ( 
.A(n_9986),
.Y(n_10384)
);

INVx3_ASAP7_75t_L g10385 ( 
.A(n_9848),
.Y(n_10385)
);

INVx2_ASAP7_75t_L g10386 ( 
.A(n_9982),
.Y(n_10386)
);

AND2x2_ASAP7_75t_L g10387 ( 
.A(n_10260),
.B(n_35),
.Y(n_10387)
);

BUFx3_ASAP7_75t_L g10388 ( 
.A(n_10002),
.Y(n_10388)
);

AND2x2_ASAP7_75t_L g10389 ( 
.A(n_10228),
.B(n_10108),
.Y(n_10389)
);

HB1xp67_ASAP7_75t_L g10390 ( 
.A(n_9826),
.Y(n_10390)
);

AND2x2_ASAP7_75t_L g10391 ( 
.A(n_10256),
.B(n_35),
.Y(n_10391)
);

NAND2xp5_ASAP7_75t_L g10392 ( 
.A(n_9847),
.B(n_37),
.Y(n_10392)
);

BUFx6f_ASAP7_75t_L g10393 ( 
.A(n_9858),
.Y(n_10393)
);

INVx2_ASAP7_75t_L g10394 ( 
.A(n_9983),
.Y(n_10394)
);

INVx2_ASAP7_75t_SL g10395 ( 
.A(n_10002),
.Y(n_10395)
);

HB1xp67_ASAP7_75t_L g10396 ( 
.A(n_10338),
.Y(n_10396)
);

INVxp67_ASAP7_75t_L g10397 ( 
.A(n_10133),
.Y(n_10397)
);

NAND2xp5_ASAP7_75t_SL g10398 ( 
.A(n_9854),
.B(n_37),
.Y(n_10398)
);

INVx2_ASAP7_75t_SL g10399 ( 
.A(n_10000),
.Y(n_10399)
);

NAND2xp5_ASAP7_75t_L g10400 ( 
.A(n_10205),
.B(n_38),
.Y(n_10400)
);

NAND2xp5_ASAP7_75t_L g10401 ( 
.A(n_9825),
.B(n_38),
.Y(n_10401)
);

AND2x2_ASAP7_75t_L g10402 ( 
.A(n_10200),
.B(n_39),
.Y(n_10402)
);

OAI21xp5_ASAP7_75t_L g10403 ( 
.A1(n_9887),
.A2(n_39),
.B(n_40),
.Y(n_10403)
);

OAI21xp5_ASAP7_75t_L g10404 ( 
.A1(n_9892),
.A2(n_40),
.B(n_41),
.Y(n_10404)
);

INVx2_ASAP7_75t_L g10405 ( 
.A(n_9992),
.Y(n_10405)
);

AND2x2_ASAP7_75t_L g10406 ( 
.A(n_10335),
.B(n_42),
.Y(n_10406)
);

AND2x6_ASAP7_75t_L g10407 ( 
.A(n_10207),
.B(n_4615),
.Y(n_10407)
);

AND2x2_ASAP7_75t_L g10408 ( 
.A(n_10342),
.B(n_42),
.Y(n_10408)
);

NOR2xp33_ASAP7_75t_L g10409 ( 
.A(n_9839),
.B(n_4616),
.Y(n_10409)
);

BUFx3_ASAP7_75t_L g10410 ( 
.A(n_9858),
.Y(n_10410)
);

OR2x2_ASAP7_75t_L g10411 ( 
.A(n_10100),
.B(n_43),
.Y(n_10411)
);

AND2x4_ASAP7_75t_L g10412 ( 
.A(n_10061),
.B(n_4617),
.Y(n_10412)
);

INVx2_ASAP7_75t_L g10413 ( 
.A(n_10027),
.Y(n_10413)
);

HB1xp67_ASAP7_75t_L g10414 ( 
.A(n_10080),
.Y(n_10414)
);

BUFx5_ASAP7_75t_L g10415 ( 
.A(n_9833),
.Y(n_10415)
);

INVx1_ASAP7_75t_L g10416 ( 
.A(n_10028),
.Y(n_10416)
);

NAND2xp5_ASAP7_75t_L g10417 ( 
.A(n_9866),
.B(n_43),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_10330),
.Y(n_10418)
);

INVx2_ASAP7_75t_L g10419 ( 
.A(n_10063),
.Y(n_10419)
);

INVx2_ASAP7_75t_L g10420 ( 
.A(n_10064),
.Y(n_10420)
);

AND2x2_ASAP7_75t_L g10421 ( 
.A(n_10271),
.B(n_10273),
.Y(n_10421)
);

AND2x2_ASAP7_75t_L g10422 ( 
.A(n_10274),
.B(n_44),
.Y(n_10422)
);

BUFx3_ASAP7_75t_L g10423 ( 
.A(n_9871),
.Y(n_10423)
);

BUFx6f_ASAP7_75t_L g10424 ( 
.A(n_10112),
.Y(n_10424)
);

NAND2xp5_ASAP7_75t_L g10425 ( 
.A(n_9961),
.B(n_45),
.Y(n_10425)
);

AND2x2_ASAP7_75t_L g10426 ( 
.A(n_10343),
.B(n_45),
.Y(n_10426)
);

INVx2_ASAP7_75t_L g10427 ( 
.A(n_10073),
.Y(n_10427)
);

NAND2xp5_ASAP7_75t_L g10428 ( 
.A(n_9844),
.B(n_46),
.Y(n_10428)
);

INVx1_ASAP7_75t_L g10429 ( 
.A(n_9841),
.Y(n_10429)
);

INVx2_ASAP7_75t_L g10430 ( 
.A(n_10183),
.Y(n_10430)
);

AND2x2_ASAP7_75t_L g10431 ( 
.A(n_10337),
.B(n_46),
.Y(n_10431)
);

BUFx2_ASAP7_75t_L g10432 ( 
.A(n_10000),
.Y(n_10432)
);

NAND2xp5_ASAP7_75t_L g10433 ( 
.A(n_9860),
.B(n_47),
.Y(n_10433)
);

INVx1_ASAP7_75t_L g10434 ( 
.A(n_9842),
.Y(n_10434)
);

AND2x2_ASAP7_75t_L g10435 ( 
.A(n_9922),
.B(n_47),
.Y(n_10435)
);

AND2x2_ASAP7_75t_L g10436 ( 
.A(n_10218),
.B(n_10220),
.Y(n_10436)
);

INVx2_ASAP7_75t_L g10437 ( 
.A(n_10194),
.Y(n_10437)
);

CKINVDCx20_ASAP7_75t_R g10438 ( 
.A(n_10195),
.Y(n_10438)
);

NAND2xp5_ASAP7_75t_L g10439 ( 
.A(n_9853),
.B(n_48),
.Y(n_10439)
);

CKINVDCx20_ASAP7_75t_R g10440 ( 
.A(n_9907),
.Y(n_10440)
);

AND2x4_ASAP7_75t_L g10441 ( 
.A(n_9840),
.B(n_4618),
.Y(n_10441)
);

INVx2_ASAP7_75t_SL g10442 ( 
.A(n_10269),
.Y(n_10442)
);

AND2x2_ASAP7_75t_L g10443 ( 
.A(n_10222),
.B(n_10233),
.Y(n_10443)
);

AND2x2_ASAP7_75t_L g10444 ( 
.A(n_10016),
.B(n_48),
.Y(n_10444)
);

INVx2_ASAP7_75t_L g10445 ( 
.A(n_10196),
.Y(n_10445)
);

INVx2_ASAP7_75t_L g10446 ( 
.A(n_10046),
.Y(n_10446)
);

AND2x2_ASAP7_75t_L g10447 ( 
.A(n_10332),
.B(n_49),
.Y(n_10447)
);

AND2x4_ASAP7_75t_L g10448 ( 
.A(n_10127),
.B(n_10339),
.Y(n_10448)
);

NAND2xp5_ASAP7_75t_L g10449 ( 
.A(n_10031),
.B(n_49),
.Y(n_10449)
);

INVx2_ASAP7_75t_L g10450 ( 
.A(n_10078),
.Y(n_10450)
);

HB1xp67_ASAP7_75t_L g10451 ( 
.A(n_10178),
.Y(n_10451)
);

AND2x2_ASAP7_75t_L g10452 ( 
.A(n_10340),
.B(n_50),
.Y(n_10452)
);

HB1xp67_ASAP7_75t_L g10453 ( 
.A(n_10272),
.Y(n_10453)
);

AND2x4_ASAP7_75t_SL g10454 ( 
.A(n_10296),
.B(n_4619),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_9850),
.Y(n_10455)
);

AND2x2_ASAP7_75t_L g10456 ( 
.A(n_10082),
.B(n_50),
.Y(n_10456)
);

OR2x2_ASAP7_75t_L g10457 ( 
.A(n_9893),
.B(n_51),
.Y(n_10457)
);

INVx2_ASAP7_75t_SL g10458 ( 
.A(n_10269),
.Y(n_10458)
);

BUFx3_ASAP7_75t_L g10459 ( 
.A(n_10160),
.Y(n_10459)
);

OR2x2_ASAP7_75t_L g10460 ( 
.A(n_9979),
.B(n_51),
.Y(n_10460)
);

AND2x4_ASAP7_75t_L g10461 ( 
.A(n_10302),
.B(n_10259),
.Y(n_10461)
);

INVx1_ASAP7_75t_SL g10462 ( 
.A(n_9837),
.Y(n_10462)
);

AND2x2_ASAP7_75t_L g10463 ( 
.A(n_10113),
.B(n_52),
.Y(n_10463)
);

INVx2_ASAP7_75t_L g10464 ( 
.A(n_10120),
.Y(n_10464)
);

INVx3_ASAP7_75t_L g10465 ( 
.A(n_10160),
.Y(n_10465)
);

AND2x2_ASAP7_75t_L g10466 ( 
.A(n_10129),
.B(n_52),
.Y(n_10466)
);

INVx2_ASAP7_75t_L g10467 ( 
.A(n_10135),
.Y(n_10467)
);

AND2x2_ASAP7_75t_L g10468 ( 
.A(n_10145),
.B(n_53),
.Y(n_10468)
);

NAND2xp5_ASAP7_75t_L g10469 ( 
.A(n_10115),
.B(n_53),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_9852),
.Y(n_10470)
);

NAND2x1p5_ASAP7_75t_L g10471 ( 
.A(n_10188),
.B(n_4620),
.Y(n_10471)
);

OAI21xp5_ASAP7_75t_L g10472 ( 
.A1(n_9938),
.A2(n_9948),
.B(n_9828),
.Y(n_10472)
);

INVx2_ASAP7_75t_L g10473 ( 
.A(n_10159),
.Y(n_10473)
);

BUFx3_ASAP7_75t_L g10474 ( 
.A(n_10188),
.Y(n_10474)
);

INVx3_ASAP7_75t_L g10475 ( 
.A(n_10136),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_9863),
.Y(n_10476)
);

AND2x2_ASAP7_75t_L g10477 ( 
.A(n_10165),
.B(n_10168),
.Y(n_10477)
);

INVx2_ASAP7_75t_L g10478 ( 
.A(n_10171),
.Y(n_10478)
);

CKINVDCx5p33_ASAP7_75t_R g10479 ( 
.A(n_9919),
.Y(n_10479)
);

HB1xp67_ASAP7_75t_L g10480 ( 
.A(n_10052),
.Y(n_10480)
);

INVx3_ASAP7_75t_L g10481 ( 
.A(n_10143),
.Y(n_10481)
);

NOR2xp67_ASAP7_75t_L g10482 ( 
.A(n_10261),
.B(n_4621),
.Y(n_10482)
);

NAND2xp5_ASAP7_75t_L g10483 ( 
.A(n_9864),
.B(n_54),
.Y(n_10483)
);

INVx2_ASAP7_75t_L g10484 ( 
.A(n_10172),
.Y(n_10484)
);

INVx1_ASAP7_75t_L g10485 ( 
.A(n_9867),
.Y(n_10485)
);

INVx2_ASAP7_75t_SL g10486 ( 
.A(n_10093),
.Y(n_10486)
);

INVx3_ASAP7_75t_SL g10487 ( 
.A(n_10109),
.Y(n_10487)
);

INVx2_ASAP7_75t_L g10488 ( 
.A(n_10175),
.Y(n_10488)
);

AND2x4_ASAP7_75t_L g10489 ( 
.A(n_10151),
.B(n_4622),
.Y(n_10489)
);

AND2x2_ASAP7_75t_L g10490 ( 
.A(n_9950),
.B(n_55),
.Y(n_10490)
);

INVxp67_ASAP7_75t_L g10491 ( 
.A(n_10041),
.Y(n_10491)
);

OR2x2_ASAP7_75t_L g10492 ( 
.A(n_9971),
.B(n_55),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_9874),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_9882),
.Y(n_10494)
);

BUFx6f_ASAP7_75t_L g10495 ( 
.A(n_9831),
.Y(n_10495)
);

INVx1_ASAP7_75t_SL g10496 ( 
.A(n_10277),
.Y(n_10496)
);

AND2x2_ASAP7_75t_L g10497 ( 
.A(n_9968),
.B(n_56),
.Y(n_10497)
);

INVx1_ASAP7_75t_L g10498 ( 
.A(n_9888),
.Y(n_10498)
);

BUFx6f_ASAP7_75t_L g10499 ( 
.A(n_10328),
.Y(n_10499)
);

AND2x2_ASAP7_75t_L g10500 ( 
.A(n_9900),
.B(n_56),
.Y(n_10500)
);

HB1xp67_ASAP7_75t_L g10501 ( 
.A(n_10076),
.Y(n_10501)
);

BUFx3_ASAP7_75t_L g10502 ( 
.A(n_10146),
.Y(n_10502)
);

INVx2_ASAP7_75t_L g10503 ( 
.A(n_9896),
.Y(n_10503)
);

BUFx6f_ASAP7_75t_L g10504 ( 
.A(n_10173),
.Y(n_10504)
);

AND2x2_ASAP7_75t_L g10505 ( 
.A(n_9939),
.B(n_58),
.Y(n_10505)
);

HB1xp67_ASAP7_75t_L g10506 ( 
.A(n_10079),
.Y(n_10506)
);

AND2x2_ASAP7_75t_L g10507 ( 
.A(n_10003),
.B(n_58),
.Y(n_10507)
);

AND2x2_ASAP7_75t_L g10508 ( 
.A(n_10092),
.B(n_59),
.Y(n_10508)
);

BUFx3_ASAP7_75t_L g10509 ( 
.A(n_9843),
.Y(n_10509)
);

AND2x2_ASAP7_75t_L g10510 ( 
.A(n_10244),
.B(n_10253),
.Y(n_10510)
);

AND2x6_ASAP7_75t_L g10511 ( 
.A(n_9845),
.B(n_4623),
.Y(n_10511)
);

AND2x2_ASAP7_75t_L g10512 ( 
.A(n_10255),
.B(n_59),
.Y(n_10512)
);

AND2x2_ASAP7_75t_L g10513 ( 
.A(n_10051),
.B(n_60),
.Y(n_10513)
);

HB1xp67_ASAP7_75t_L g10514 ( 
.A(n_10251),
.Y(n_10514)
);

AND2x2_ASAP7_75t_L g10515 ( 
.A(n_10055),
.B(n_61),
.Y(n_10515)
);

NAND2xp5_ASAP7_75t_L g10516 ( 
.A(n_9838),
.B(n_10067),
.Y(n_10516)
);

AND2x6_ASAP7_75t_L g10517 ( 
.A(n_10124),
.B(n_4624),
.Y(n_10517)
);

CKINVDCx5p33_ASAP7_75t_R g10518 ( 
.A(n_10109),
.Y(n_10518)
);

INVx4_ASAP7_75t_L g10519 ( 
.A(n_10109),
.Y(n_10519)
);

INVx4_ASAP7_75t_L g10520 ( 
.A(n_10065),
.Y(n_10520)
);

AND2x2_ASAP7_75t_L g10521 ( 
.A(n_10020),
.B(n_61),
.Y(n_10521)
);

INVx2_ASAP7_75t_L g10522 ( 
.A(n_9912),
.Y(n_10522)
);

INVx3_ASAP7_75t_L g10523 ( 
.A(n_10163),
.Y(n_10523)
);

BUFx6f_ASAP7_75t_L g10524 ( 
.A(n_10065),
.Y(n_10524)
);

INVx2_ASAP7_75t_L g10525 ( 
.A(n_9914),
.Y(n_10525)
);

INVx2_ASAP7_75t_SL g10526 ( 
.A(n_10162),
.Y(n_10526)
);

NAND2xp5_ASAP7_75t_L g10527 ( 
.A(n_9865),
.B(n_62),
.Y(n_10527)
);

NOR2xp33_ASAP7_75t_L g10528 ( 
.A(n_9836),
.B(n_4625),
.Y(n_10528)
);

AND2x4_ASAP7_75t_L g10529 ( 
.A(n_10298),
.B(n_10297),
.Y(n_10529)
);

INVxp67_ASAP7_75t_SL g10530 ( 
.A(n_10049),
.Y(n_10530)
);

INVx1_ASAP7_75t_L g10531 ( 
.A(n_9920),
.Y(n_10531)
);

OR2x6_ASAP7_75t_L g10532 ( 
.A(n_10114),
.B(n_4626),
.Y(n_10532)
);

NAND2xp5_ASAP7_75t_L g10533 ( 
.A(n_9890),
.B(n_62),
.Y(n_10533)
);

BUFx2_ASAP7_75t_L g10534 ( 
.A(n_10181),
.Y(n_10534)
);

OAI21xp5_ASAP7_75t_L g10535 ( 
.A1(n_10291),
.A2(n_63),
.B(n_64),
.Y(n_10535)
);

INVx2_ASAP7_75t_L g10536 ( 
.A(n_9927),
.Y(n_10536)
);

NAND2xp5_ASAP7_75t_L g10537 ( 
.A(n_9898),
.B(n_63),
.Y(n_10537)
);

NAND2xp5_ASAP7_75t_L g10538 ( 
.A(n_9901),
.B(n_65),
.Y(n_10538)
);

INVx3_ASAP7_75t_L g10539 ( 
.A(n_9869),
.Y(n_10539)
);

AND2x2_ASAP7_75t_L g10540 ( 
.A(n_10038),
.B(n_65),
.Y(n_10540)
);

INVx2_ASAP7_75t_L g10541 ( 
.A(n_9929),
.Y(n_10541)
);

INVx1_ASAP7_75t_L g10542 ( 
.A(n_9930),
.Y(n_10542)
);

OR2x6_ASAP7_75t_L g10543 ( 
.A(n_10114),
.B(n_4627),
.Y(n_10543)
);

INVx3_ASAP7_75t_L g10544 ( 
.A(n_9973),
.Y(n_10544)
);

BUFx6f_ASAP7_75t_L g10545 ( 
.A(n_10197),
.Y(n_10545)
);

INVx2_ASAP7_75t_SL g10546 ( 
.A(n_10229),
.Y(n_10546)
);

INVx2_ASAP7_75t_L g10547 ( 
.A(n_9933),
.Y(n_10547)
);

INVx1_ASAP7_75t_SL g10548 ( 
.A(n_10270),
.Y(n_10548)
);

AND2x2_ASAP7_75t_L g10549 ( 
.A(n_10050),
.B(n_66),
.Y(n_10549)
);

HB1xp67_ASAP7_75t_L g10550 ( 
.A(n_10245),
.Y(n_10550)
);

HB1xp67_ASAP7_75t_L g10551 ( 
.A(n_10246),
.Y(n_10551)
);

AND2x2_ASAP7_75t_L g10552 ( 
.A(n_10071),
.B(n_66),
.Y(n_10552)
);

INVx2_ASAP7_75t_L g10553 ( 
.A(n_9941),
.Y(n_10553)
);

INVx1_ASAP7_75t_SL g10554 ( 
.A(n_10174),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_10074),
.B(n_67),
.Y(n_10555)
);

NAND2xp5_ASAP7_75t_L g10556 ( 
.A(n_9904),
.B(n_68),
.Y(n_10556)
);

BUFx6f_ASAP7_75t_L g10557 ( 
.A(n_10203),
.Y(n_10557)
);

AND2x2_ASAP7_75t_L g10558 ( 
.A(n_9975),
.B(n_68),
.Y(n_10558)
);

AND2x2_ASAP7_75t_L g10559 ( 
.A(n_10208),
.B(n_69),
.Y(n_10559)
);

INVx2_ASAP7_75t_SL g10560 ( 
.A(n_9946),
.Y(n_10560)
);

NAND2xp5_ASAP7_75t_L g10561 ( 
.A(n_9905),
.B(n_69),
.Y(n_10561)
);

INVx1_ASAP7_75t_SL g10562 ( 
.A(n_9862),
.Y(n_10562)
);

AND2x2_ASAP7_75t_L g10563 ( 
.A(n_10213),
.B(n_70),
.Y(n_10563)
);

INVx1_ASAP7_75t_L g10564 ( 
.A(n_9943),
.Y(n_10564)
);

AND2x2_ASAP7_75t_L g10565 ( 
.A(n_10341),
.B(n_10029),
.Y(n_10565)
);

BUFx6f_ASAP7_75t_L g10566 ( 
.A(n_9954),
.Y(n_10566)
);

AND2x2_ASAP7_75t_L g10567 ( 
.A(n_10216),
.B(n_70),
.Y(n_10567)
);

AND2x2_ASAP7_75t_L g10568 ( 
.A(n_10224),
.B(n_71),
.Y(n_10568)
);

BUFx8_ASAP7_75t_SL g10569 ( 
.A(n_9945),
.Y(n_10569)
);

NOR2xp33_ASAP7_75t_L g10570 ( 
.A(n_10004),
.B(n_4628),
.Y(n_10570)
);

HB1xp67_ASAP7_75t_L g10571 ( 
.A(n_10249),
.Y(n_10571)
);

NAND2xp5_ASAP7_75t_L g10572 ( 
.A(n_9911),
.B(n_71),
.Y(n_10572)
);

BUFx3_ASAP7_75t_L g10573 ( 
.A(n_10243),
.Y(n_10573)
);

OR2x6_ASAP7_75t_L g10574 ( 
.A(n_10313),
.B(n_4630),
.Y(n_10574)
);

NOR2xp33_ASAP7_75t_L g10575 ( 
.A(n_9849),
.B(n_4631),
.Y(n_10575)
);

NAND2xp5_ASAP7_75t_L g10576 ( 
.A(n_9918),
.B(n_72),
.Y(n_10576)
);

INVx2_ASAP7_75t_L g10577 ( 
.A(n_9963),
.Y(n_10577)
);

INVx1_ASAP7_75t_SL g10578 ( 
.A(n_10286),
.Y(n_10578)
);

AND2x2_ASAP7_75t_L g10579 ( 
.A(n_10230),
.B(n_73),
.Y(n_10579)
);

AOI22xp5_ASAP7_75t_L g10580 ( 
.A1(n_10032),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_10580)
);

INVx1_ASAP7_75t_L g10581 ( 
.A(n_9978),
.Y(n_10581)
);

INVx2_ASAP7_75t_L g10582 ( 
.A(n_9997),
.Y(n_10582)
);

AND2x2_ASAP7_75t_L g10583 ( 
.A(n_10231),
.B(n_74),
.Y(n_10583)
);

INVx1_ASAP7_75t_SL g10584 ( 
.A(n_10281),
.Y(n_10584)
);

INVx2_ASAP7_75t_L g10585 ( 
.A(n_9998),
.Y(n_10585)
);

INVx1_ASAP7_75t_L g10586 ( 
.A(n_10007),
.Y(n_10586)
);

BUFx3_ASAP7_75t_L g10587 ( 
.A(n_10326),
.Y(n_10587)
);

AND2x2_ASAP7_75t_L g10588 ( 
.A(n_10237),
.B(n_10242),
.Y(n_10588)
);

BUFx3_ASAP7_75t_L g10589 ( 
.A(n_10308),
.Y(n_10589)
);

OAI21xp5_ASAP7_75t_L g10590 ( 
.A1(n_9883),
.A2(n_10333),
.B(n_9921),
.Y(n_10590)
);

HB1xp67_ASAP7_75t_L g10591 ( 
.A(n_10234),
.Y(n_10591)
);

INVxp33_ASAP7_75t_L g10592 ( 
.A(n_10247),
.Y(n_10592)
);

INVxp67_ASAP7_75t_L g10593 ( 
.A(n_10148),
.Y(n_10593)
);

INVx2_ASAP7_75t_SL g10594 ( 
.A(n_9964),
.Y(n_10594)
);

NAND2xp5_ASAP7_75t_L g10595 ( 
.A(n_9924),
.B(n_75),
.Y(n_10595)
);

AND2x2_ASAP7_75t_L g10596 ( 
.A(n_10040),
.B(n_77),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_10013),
.Y(n_10597)
);

INVx2_ASAP7_75t_L g10598 ( 
.A(n_10015),
.Y(n_10598)
);

INVx1_ASAP7_75t_L g10599 ( 
.A(n_10019),
.Y(n_10599)
);

INVx1_ASAP7_75t_L g10600 ( 
.A(n_10034),
.Y(n_10600)
);

INVx3_ASAP7_75t_L g10601 ( 
.A(n_10214),
.Y(n_10601)
);

INVxp33_ASAP7_75t_L g10602 ( 
.A(n_10149),
.Y(n_10602)
);

INVx3_ASAP7_75t_L g10603 ( 
.A(n_10221),
.Y(n_10603)
);

NAND2xp5_ASAP7_75t_L g10604 ( 
.A(n_9936),
.B(n_78),
.Y(n_10604)
);

NAND2xp5_ASAP7_75t_L g10605 ( 
.A(n_9937),
.B(n_78),
.Y(n_10605)
);

INVx1_ASAP7_75t_SL g10606 ( 
.A(n_10287),
.Y(n_10606)
);

AND2x2_ASAP7_75t_L g10607 ( 
.A(n_10042),
.B(n_10043),
.Y(n_10607)
);

INVx2_ASAP7_75t_L g10608 ( 
.A(n_10139),
.Y(n_10608)
);

AND2x2_ASAP7_75t_L g10609 ( 
.A(n_10169),
.B(n_79),
.Y(n_10609)
);

AND2x2_ASAP7_75t_L g10610 ( 
.A(n_10170),
.B(n_79),
.Y(n_10610)
);

CKINVDCx20_ASAP7_75t_R g10611 ( 
.A(n_10257),
.Y(n_10611)
);

INVx3_ASAP7_75t_L g10612 ( 
.A(n_10294),
.Y(n_10612)
);

INVx3_ASAP7_75t_L g10613 ( 
.A(n_10236),
.Y(n_10613)
);

AND2x2_ASAP7_75t_L g10614 ( 
.A(n_10154),
.B(n_80),
.Y(n_10614)
);

INVx1_ASAP7_75t_SL g10615 ( 
.A(n_10290),
.Y(n_10615)
);

NOR2xp33_ASAP7_75t_L g10616 ( 
.A(n_10227),
.B(n_4632),
.Y(n_10616)
);

AND2x2_ASAP7_75t_L g10617 ( 
.A(n_10156),
.B(n_80),
.Y(n_10617)
);

INVx2_ASAP7_75t_L g10618 ( 
.A(n_10077),
.Y(n_10618)
);

HB1xp67_ASAP7_75t_L g10619 ( 
.A(n_10276),
.Y(n_10619)
);

AND2x2_ASAP7_75t_L g10620 ( 
.A(n_10161),
.B(n_81),
.Y(n_10620)
);

INVx2_ASAP7_75t_L g10621 ( 
.A(n_10087),
.Y(n_10621)
);

AND2x2_ASAP7_75t_L g10622 ( 
.A(n_10166),
.B(n_81),
.Y(n_10622)
);

OAI21xp5_ASAP7_75t_L g10623 ( 
.A1(n_9917),
.A2(n_82),
.B(n_83),
.Y(n_10623)
);

INVxp67_ASAP7_75t_L g10624 ( 
.A(n_10204),
.Y(n_10624)
);

INVx3_ASAP7_75t_L g10625 ( 
.A(n_9965),
.Y(n_10625)
);

OR2x2_ASAP7_75t_L g10626 ( 
.A(n_9942),
.B(n_82),
.Y(n_10626)
);

INVx1_ASAP7_75t_L g10627 ( 
.A(n_10101),
.Y(n_10627)
);

NAND2xp5_ASAP7_75t_L g10628 ( 
.A(n_10176),
.B(n_83),
.Y(n_10628)
);

AND2x2_ASAP7_75t_L g10629 ( 
.A(n_10182),
.B(n_84),
.Y(n_10629)
);

INVx1_ASAP7_75t_L g10630 ( 
.A(n_10111),
.Y(n_10630)
);

INVx1_ASAP7_75t_L g10631 ( 
.A(n_10118),
.Y(n_10631)
);

INVx2_ASAP7_75t_L g10632 ( 
.A(n_10119),
.Y(n_10632)
);

AND2x2_ASAP7_75t_L g10633 ( 
.A(n_10189),
.B(n_84),
.Y(n_10633)
);

NAND2xp5_ASAP7_75t_L g10634 ( 
.A(n_9879),
.B(n_85),
.Y(n_10634)
);

INVx2_ASAP7_75t_SL g10635 ( 
.A(n_10090),
.Y(n_10635)
);

OAI21xp5_ASAP7_75t_L g10636 ( 
.A1(n_10085),
.A2(n_85),
.B(n_87),
.Y(n_10636)
);

INVx1_ASAP7_75t_SL g10637 ( 
.A(n_10018),
.Y(n_10637)
);

NAND2xp5_ASAP7_75t_SL g10638 ( 
.A(n_10069),
.B(n_87),
.Y(n_10638)
);

AND2x2_ASAP7_75t_L g10639 ( 
.A(n_10192),
.B(n_10075),
.Y(n_10639)
);

NAND2xp5_ASAP7_75t_L g10640 ( 
.A(n_10177),
.B(n_88),
.Y(n_10640)
);

HB1xp67_ASAP7_75t_L g10641 ( 
.A(n_10132),
.Y(n_10641)
);

INVx4_ASAP7_75t_L g10642 ( 
.A(n_10309),
.Y(n_10642)
);

AND2x2_ASAP7_75t_L g10643 ( 
.A(n_9931),
.B(n_89),
.Y(n_10643)
);

OR2x2_ASAP7_75t_L g10644 ( 
.A(n_9974),
.B(n_89),
.Y(n_10644)
);

BUFx3_ASAP7_75t_L g10645 ( 
.A(n_10316),
.Y(n_10645)
);

NAND2xp5_ASAP7_75t_SL g10646 ( 
.A(n_9859),
.B(n_90),
.Y(n_10646)
);

NAND2xp5_ASAP7_75t_L g10647 ( 
.A(n_10198),
.B(n_90),
.Y(n_10647)
);

AND2x2_ASAP7_75t_L g10648 ( 
.A(n_9889),
.B(n_91),
.Y(n_10648)
);

BUFx3_ASAP7_75t_L g10649 ( 
.A(n_10320),
.Y(n_10649)
);

INVx3_ASAP7_75t_L g10650 ( 
.A(n_10138),
.Y(n_10650)
);

INVx2_ASAP7_75t_L g10651 ( 
.A(n_10179),
.Y(n_10651)
);

INVx3_ASAP7_75t_L g10652 ( 
.A(n_10187),
.Y(n_10652)
);

BUFx6f_ASAP7_75t_L g10653 ( 
.A(n_10322),
.Y(n_10653)
);

HB1xp67_ASAP7_75t_L g10654 ( 
.A(n_10190),
.Y(n_10654)
);

INVx2_ASAP7_75t_L g10655 ( 
.A(n_10201),
.Y(n_10655)
);

INVx2_ASAP7_75t_SL g10656 ( 
.A(n_10068),
.Y(n_10656)
);

INVx2_ASAP7_75t_L g10657 ( 
.A(n_10210),
.Y(n_10657)
);

INVx2_ASAP7_75t_L g10658 ( 
.A(n_10057),
.Y(n_10658)
);

INVx1_ASAP7_75t_L g10659 ( 
.A(n_10116),
.Y(n_10659)
);

OAI21xp5_ASAP7_75t_L g10660 ( 
.A1(n_10103),
.A2(n_91),
.B(n_92),
.Y(n_10660)
);

NAND2xp5_ASAP7_75t_L g10661 ( 
.A(n_10217),
.B(n_92),
.Y(n_10661)
);

NOR2xp33_ASAP7_75t_SL g10662 ( 
.A(n_10319),
.B(n_4633),
.Y(n_10662)
);

INVx1_ASAP7_75t_L g10663 ( 
.A(n_10117),
.Y(n_10663)
);

BUFx6f_ASAP7_75t_L g10664 ( 
.A(n_10180),
.Y(n_10664)
);

INVx1_ASAP7_75t_L g10665 ( 
.A(n_10121),
.Y(n_10665)
);

INVx1_ASAP7_75t_L g10666 ( 
.A(n_10123),
.Y(n_10666)
);

OAI21xp5_ASAP7_75t_L g10667 ( 
.A1(n_10104),
.A2(n_93),
.B(n_94),
.Y(n_10667)
);

INVx2_ASAP7_75t_L g10668 ( 
.A(n_9908),
.Y(n_10668)
);

INVx1_ASAP7_75t_SL g10669 ( 
.A(n_9932),
.Y(n_10669)
);

INVx2_ASAP7_75t_L g10670 ( 
.A(n_9908),
.Y(n_10670)
);

INVx1_ASAP7_75t_L g10671 ( 
.A(n_10125),
.Y(n_10671)
);

INVx2_ASAP7_75t_L g10672 ( 
.A(n_9908),
.Y(n_10672)
);

BUFx12f_ASAP7_75t_L g10673 ( 
.A(n_10035),
.Y(n_10673)
);

INVx1_ASAP7_75t_L g10674 ( 
.A(n_10130),
.Y(n_10674)
);

NAND2xp5_ASAP7_75t_L g10675 ( 
.A(n_10225),
.B(n_94),
.Y(n_10675)
);

NAND2xp5_ASAP7_75t_L g10676 ( 
.A(n_10184),
.B(n_95),
.Y(n_10676)
);

OAI21xp5_ASAP7_75t_L g10677 ( 
.A1(n_10086),
.A2(n_95),
.B(n_96),
.Y(n_10677)
);

HB1xp67_ASAP7_75t_L g10678 ( 
.A(n_10289),
.Y(n_10678)
);

INVxp33_ASAP7_75t_L g10679 ( 
.A(n_10265),
.Y(n_10679)
);

BUFx3_ASAP7_75t_L g10680 ( 
.A(n_10293),
.Y(n_10680)
);

NAND2xp5_ASAP7_75t_L g10681 ( 
.A(n_9855),
.B(n_96),
.Y(n_10681)
);

INVx3_ASAP7_75t_L g10682 ( 
.A(n_10288),
.Y(n_10682)
);

AND2x2_ASAP7_75t_L g10683 ( 
.A(n_10258),
.B(n_97),
.Y(n_10683)
);

AND2x2_ASAP7_75t_L g10684 ( 
.A(n_9910),
.B(n_98),
.Y(n_10684)
);

OAI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_9955),
.A2(n_98),
.B(n_99),
.Y(n_10685)
);

AND2x2_ASAP7_75t_L g10686 ( 
.A(n_9959),
.B(n_99),
.Y(n_10686)
);

INVxp33_ASAP7_75t_L g10687 ( 
.A(n_10278),
.Y(n_10687)
);

INVx2_ASAP7_75t_L g10688 ( 
.A(n_9908),
.Y(n_10688)
);

NAND2xp5_ASAP7_75t_L g10689 ( 
.A(n_10223),
.B(n_100),
.Y(n_10689)
);

OAI21xp5_ASAP7_75t_L g10690 ( 
.A1(n_10023),
.A2(n_100),
.B(n_101),
.Y(n_10690)
);

BUFx4f_ASAP7_75t_L g10691 ( 
.A(n_10306),
.Y(n_10691)
);

NOR2xp33_ASAP7_75t_L g10692 ( 
.A(n_9872),
.B(n_4634),
.Y(n_10692)
);

AND2x4_ASAP7_75t_SL g10693 ( 
.A(n_10313),
.B(n_10248),
.Y(n_10693)
);

INVx1_ASAP7_75t_L g10694 ( 
.A(n_10134),
.Y(n_10694)
);

INVx2_ASAP7_75t_SL g10695 ( 
.A(n_10089),
.Y(n_10695)
);

INVx1_ASAP7_75t_L g10696 ( 
.A(n_10137),
.Y(n_10696)
);

INVx1_ASAP7_75t_L g10697 ( 
.A(n_10140),
.Y(n_10697)
);

AND2x2_ASAP7_75t_L g10698 ( 
.A(n_9993),
.B(n_102),
.Y(n_10698)
);

INVx2_ASAP7_75t_L g10699 ( 
.A(n_10193),
.Y(n_10699)
);

NAND2xp5_ASAP7_75t_L g10700 ( 
.A(n_9851),
.B(n_102),
.Y(n_10700)
);

AND2x2_ASAP7_75t_L g10701 ( 
.A(n_10024),
.B(n_103),
.Y(n_10701)
);

INVx3_ASAP7_75t_L g10702 ( 
.A(n_10306),
.Y(n_10702)
);

NAND2xp5_ASAP7_75t_SL g10703 ( 
.A(n_9880),
.B(n_103),
.Y(n_10703)
);

AND2x2_ASAP7_75t_L g10704 ( 
.A(n_10009),
.B(n_104),
.Y(n_10704)
);

NAND2xp5_ASAP7_75t_SL g10705 ( 
.A(n_10263),
.B(n_104),
.Y(n_10705)
);

AND2x2_ASAP7_75t_L g10706 ( 
.A(n_10215),
.B(n_105),
.Y(n_10706)
);

HB1xp67_ASAP7_75t_L g10707 ( 
.A(n_10106),
.Y(n_10707)
);

OAI21xp33_ASAP7_75t_L g10708 ( 
.A1(n_9976),
.A2(n_106),
.B(n_107),
.Y(n_10708)
);

BUFx3_ASAP7_75t_L g10709 ( 
.A(n_10293),
.Y(n_10709)
);

INVx1_ASAP7_75t_SL g10710 ( 
.A(n_9985),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_SL g10711 ( 
.A(n_9824),
.B(n_106),
.Y(n_10711)
);

INVx2_ASAP7_75t_L g10712 ( 
.A(n_10193),
.Y(n_10712)
);

BUFx6f_ASAP7_75t_L g10713 ( 
.A(n_10303),
.Y(n_10713)
);

NAND2x1p5_ASAP7_75t_L g10714 ( 
.A(n_10048),
.B(n_4635),
.Y(n_10714)
);

NAND2xp5_ASAP7_75t_L g10715 ( 
.A(n_9991),
.B(n_107),
.Y(n_10715)
);

BUFx3_ASAP7_75t_L g10716 ( 
.A(n_10293),
.Y(n_10716)
);

AND2x2_ASAP7_75t_L g10717 ( 
.A(n_10095),
.B(n_108),
.Y(n_10717)
);

NOR2xp33_ASAP7_75t_L g10718 ( 
.A(n_9925),
.B(n_4636),
.Y(n_10718)
);

INVx2_ASAP7_75t_L g10719 ( 
.A(n_10193),
.Y(n_10719)
);

AND2x2_ASAP7_75t_SL g10720 ( 
.A(n_10299),
.B(n_108),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_10081),
.B(n_109),
.Y(n_10721)
);

INVx3_ASAP7_75t_SL g10722 ( 
.A(n_10212),
.Y(n_10722)
);

NAND2xp5_ASAP7_75t_L g10723 ( 
.A(n_10282),
.B(n_109),
.Y(n_10723)
);

NAND2xp5_ASAP7_75t_L g10724 ( 
.A(n_9875),
.B(n_9999),
.Y(n_10724)
);

INVx1_ASAP7_75t_L g10725 ( 
.A(n_10141),
.Y(n_10725)
);

AND2x2_ASAP7_75t_L g10726 ( 
.A(n_10083),
.B(n_110),
.Y(n_10726)
);

INVx1_ASAP7_75t_SL g10727 ( 
.A(n_9915),
.Y(n_10727)
);

BUFx4f_ASAP7_75t_L g10728 ( 
.A(n_10306),
.Y(n_10728)
);

NAND2xp5_ASAP7_75t_L g10729 ( 
.A(n_10001),
.B(n_110),
.Y(n_10729)
);

INVx2_ASAP7_75t_SL g10730 ( 
.A(n_10209),
.Y(n_10730)
);

NAND2xp5_ASAP7_75t_L g10731 ( 
.A(n_10097),
.B(n_111),
.Y(n_10731)
);

BUFx3_ASAP7_75t_L g10732 ( 
.A(n_10293),
.Y(n_10732)
);

INVx1_ASAP7_75t_L g10733 ( 
.A(n_10150),
.Y(n_10733)
);

AND2x2_ASAP7_75t_L g10734 ( 
.A(n_10084),
.B(n_111),
.Y(n_10734)
);

NAND2xp5_ASAP7_75t_L g10735 ( 
.A(n_9895),
.B(n_9916),
.Y(n_10735)
);

INVx3_ASAP7_75t_L g10736 ( 
.A(n_10310),
.Y(n_10736)
);

NOR2xp33_ASAP7_75t_L g10737 ( 
.A(n_9926),
.B(n_9944),
.Y(n_10737)
);

AND2x2_ASAP7_75t_L g10738 ( 
.A(n_10191),
.B(n_112),
.Y(n_10738)
);

AND2x2_ASAP7_75t_L g10739 ( 
.A(n_10199),
.B(n_112),
.Y(n_10739)
);

INVx1_ASAP7_75t_L g10740 ( 
.A(n_10153),
.Y(n_10740)
);

NAND2xp5_ASAP7_75t_L g10741 ( 
.A(n_9951),
.B(n_114),
.Y(n_10741)
);

INVx2_ASAP7_75t_L g10742 ( 
.A(n_10193),
.Y(n_10742)
);

BUFx4_ASAP7_75t_SL g10743 ( 
.A(n_10240),
.Y(n_10743)
);

AND2x2_ASAP7_75t_L g10744 ( 
.A(n_10157),
.B(n_114),
.Y(n_10744)
);

OAI21xp5_ASAP7_75t_L g10745 ( 
.A1(n_10235),
.A2(n_115),
.B(n_116),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_10164),
.Y(n_10746)
);

INVxp67_ASAP7_75t_SL g10747 ( 
.A(n_9876),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_10167),
.Y(n_10748)
);

INVxp67_ASAP7_75t_L g10749 ( 
.A(n_9969),
.Y(n_10749)
);

AND2x2_ASAP7_75t_L g10750 ( 
.A(n_10267),
.B(n_115),
.Y(n_10750)
);

CKINVDCx5p33_ASAP7_75t_R g10751 ( 
.A(n_10025),
.Y(n_10751)
);

AND2x4_ASAP7_75t_L g10752 ( 
.A(n_10147),
.B(n_10152),
.Y(n_10752)
);

AND2x2_ASAP7_75t_L g10753 ( 
.A(n_10241),
.B(n_116),
.Y(n_10753)
);

BUFx3_ASAP7_75t_L g10754 ( 
.A(n_10307),
.Y(n_10754)
);

INVx2_ASAP7_75t_SL g10755 ( 
.A(n_9832),
.Y(n_10755)
);

INVx2_ASAP7_75t_L g10756 ( 
.A(n_10211),
.Y(n_10756)
);

INVx1_ASAP7_75t_L g10757 ( 
.A(n_10036),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_L g10758 ( 
.A(n_10008),
.B(n_117),
.Y(n_10758)
);

NOR2xp33_ASAP7_75t_R g10759 ( 
.A(n_9984),
.B(n_4637),
.Y(n_10759)
);

INVx2_ASAP7_75t_SL g10760 ( 
.A(n_10056),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_10039),
.Y(n_10761)
);

HB1xp67_ASAP7_75t_L g10762 ( 
.A(n_10044),
.Y(n_10762)
);

AND2x2_ASAP7_75t_L g10763 ( 
.A(n_10262),
.B(n_117),
.Y(n_10763)
);

AND2x2_ASAP7_75t_L g10764 ( 
.A(n_10311),
.B(n_118),
.Y(n_10764)
);

AND2x2_ASAP7_75t_L g10765 ( 
.A(n_10321),
.B(n_118),
.Y(n_10765)
);

AND2x2_ASAP7_75t_L g10766 ( 
.A(n_10285),
.B(n_9947),
.Y(n_10766)
);

NAND2x1p5_ASAP7_75t_L g10767 ( 
.A(n_9957),
.B(n_4638),
.Y(n_10767)
);

AND2x2_ASAP7_75t_SL g10768 ( 
.A(n_10300),
.B(n_10317),
.Y(n_10768)
);

NAND2xp5_ASAP7_75t_L g10769 ( 
.A(n_10010),
.B(n_119),
.Y(n_10769)
);

INVx2_ASAP7_75t_L g10770 ( 
.A(n_10047),
.Y(n_10770)
);

HB1xp67_ASAP7_75t_L g10771 ( 
.A(n_10053),
.Y(n_10771)
);

INVx1_ASAP7_75t_L g10772 ( 
.A(n_10058),
.Y(n_10772)
);

INVx1_ASAP7_75t_L g10773 ( 
.A(n_10059),
.Y(n_10773)
);

AND2x2_ASAP7_75t_L g10774 ( 
.A(n_9981),
.B(n_120),
.Y(n_10774)
);

NAND2xp5_ASAP7_75t_L g10775 ( 
.A(n_10011),
.B(n_121),
.Y(n_10775)
);

NAND2x1p5_ASAP7_75t_L g10776 ( 
.A(n_9953),
.B(n_4640),
.Y(n_10776)
);

INVx1_ASAP7_75t_L g10777 ( 
.A(n_10060),
.Y(n_10777)
);

INVx1_ASAP7_75t_L g10778 ( 
.A(n_10062),
.Y(n_10778)
);

INVx2_ASAP7_75t_L g10779 ( 
.A(n_10070),
.Y(n_10779)
);

INVxp67_ASAP7_75t_L g10780 ( 
.A(n_10142),
.Y(n_10780)
);

AND2x2_ASAP7_75t_L g10781 ( 
.A(n_10323),
.B(n_121),
.Y(n_10781)
);

AND2x2_ASAP7_75t_L g10782 ( 
.A(n_10334),
.B(n_122),
.Y(n_10782)
);

NAND2xp5_ASAP7_75t_L g10783 ( 
.A(n_10012),
.B(n_122),
.Y(n_10783)
);

INVx1_ASAP7_75t_L g10784 ( 
.A(n_9977),
.Y(n_10784)
);

INVx2_ASAP7_75t_L g10785 ( 
.A(n_9988),
.Y(n_10785)
);

BUFx3_ASAP7_75t_L g10786 ( 
.A(n_10280),
.Y(n_10786)
);

NAND2xp5_ASAP7_75t_L g10787 ( 
.A(n_10017),
.B(n_123),
.Y(n_10787)
);

AND2x2_ASAP7_75t_L g10788 ( 
.A(n_10126),
.B(n_123),
.Y(n_10788)
);

HB1xp67_ASAP7_75t_L g10789 ( 
.A(n_10155),
.Y(n_10789)
);

BUFx6f_ASAP7_75t_L g10790 ( 
.A(n_10158),
.Y(n_10790)
);

BUFx6f_ASAP7_75t_L g10791 ( 
.A(n_10096),
.Y(n_10791)
);

NAND2xp5_ASAP7_75t_L g10792 ( 
.A(n_10022),
.B(n_124),
.Y(n_10792)
);

INVx1_ASAP7_75t_L g10793 ( 
.A(n_9990),
.Y(n_10793)
);

AND2x4_ASAP7_75t_L g10794 ( 
.A(n_10099),
.B(n_4641),
.Y(n_10794)
);

INVxp67_ASAP7_75t_L g10795 ( 
.A(n_10105),
.Y(n_10795)
);

AND2x6_ASAP7_75t_L g10796 ( 
.A(n_10301),
.B(n_4642),
.Y(n_10796)
);

INVx2_ASAP7_75t_L g10797 ( 
.A(n_9994),
.Y(n_10797)
);

NAND2xp5_ASAP7_75t_L g10798 ( 
.A(n_10026),
.B(n_9995),
.Y(n_10798)
);

BUFx6f_ASAP7_75t_L g10799 ( 
.A(n_10254),
.Y(n_10799)
);

INVxp33_ASAP7_75t_L g10800 ( 
.A(n_10226),
.Y(n_10800)
);

AND2x2_ASAP7_75t_L g10801 ( 
.A(n_10327),
.B(n_124),
.Y(n_10801)
);

AND2x2_ASAP7_75t_L g10802 ( 
.A(n_10304),
.B(n_125),
.Y(n_10802)
);

NAND2xp5_ASAP7_75t_L g10803 ( 
.A(n_10006),
.B(n_125),
.Y(n_10803)
);

INVx1_ASAP7_75t_L g10804 ( 
.A(n_10122),
.Y(n_10804)
);

BUFx3_ASAP7_75t_L g10805 ( 
.A(n_10283),
.Y(n_10805)
);

NOR2xp33_ASAP7_75t_L g10806 ( 
.A(n_10232),
.B(n_4643),
.Y(n_10806)
);

HB1xp67_ASAP7_75t_L g10807 ( 
.A(n_10268),
.Y(n_10807)
);

AND2x2_ASAP7_75t_SL g10808 ( 
.A(n_10279),
.B(n_126),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_9906),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_10066),
.Y(n_10810)
);

INVx2_ASAP7_75t_L g10811 ( 
.A(n_10275),
.Y(n_10811)
);

AND2x2_ASAP7_75t_SL g10812 ( 
.A(n_10206),
.B(n_127),
.Y(n_10812)
);

NAND2xp5_ASAP7_75t_L g10813 ( 
.A(n_10033),
.B(n_127),
.Y(n_10813)
);

HB1xp67_ASAP7_75t_L g10814 ( 
.A(n_10144),
.Y(n_10814)
);

AND2x2_ASAP7_75t_L g10815 ( 
.A(n_10305),
.B(n_10312),
.Y(n_10815)
);

AND2x2_ASAP7_75t_L g10816 ( 
.A(n_10324),
.B(n_10295),
.Y(n_10816)
);

INVx2_ASAP7_75t_SL g10817 ( 
.A(n_9958),
.Y(n_10817)
);

INVx3_ASAP7_75t_L g10818 ( 
.A(n_10252),
.Y(n_10818)
);

INVx3_ASAP7_75t_L g10819 ( 
.A(n_10250),
.Y(n_10819)
);

BUFx6f_ASAP7_75t_L g10820 ( 
.A(n_10185),
.Y(n_10820)
);

INVx1_ASAP7_75t_SL g10821 ( 
.A(n_10186),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_10030),
.Y(n_10822)
);

BUFx3_ASAP7_75t_L g10823 ( 
.A(n_9877),
.Y(n_10823)
);

INVx1_ASAP7_75t_L g10824 ( 
.A(n_9891),
.Y(n_10824)
);

CKINVDCx5p33_ASAP7_75t_R g10825 ( 
.A(n_9902),
.Y(n_10825)
);

AND2x4_ASAP7_75t_L g10826 ( 
.A(n_9972),
.B(n_4644),
.Y(n_10826)
);

AND2x2_ASAP7_75t_L g10827 ( 
.A(n_10088),
.B(n_129),
.Y(n_10827)
);

INVx2_ASAP7_75t_L g10828 ( 
.A(n_10264),
.Y(n_10828)
);

INVx1_ASAP7_75t_L g10829 ( 
.A(n_9903),
.Y(n_10829)
);

INVx1_ASAP7_75t_L g10830 ( 
.A(n_9987),
.Y(n_10830)
);

BUFx3_ASAP7_75t_L g10831 ( 
.A(n_10239),
.Y(n_10831)
);

INVx2_ASAP7_75t_L g10832 ( 
.A(n_10102),
.Y(n_10832)
);

NAND2xp5_ASAP7_75t_SL g10833 ( 
.A(n_10219),
.B(n_129),
.Y(n_10833)
);

NAND2x1p5_ASAP7_75t_L g10834 ( 
.A(n_10314),
.B(n_4645),
.Y(n_10834)
);

AND2x2_ASAP7_75t_L g10835 ( 
.A(n_10037),
.B(n_10131),
.Y(n_10835)
);

NAND2xp5_ASAP7_75t_L g10836 ( 
.A(n_9970),
.B(n_130),
.Y(n_10836)
);

AND2x4_ASAP7_75t_L g10837 ( 
.A(n_9980),
.B(n_4646),
.Y(n_10837)
);

NAND2xp5_ASAP7_75t_L g10838 ( 
.A(n_9989),
.B(n_10098),
.Y(n_10838)
);

INVx2_ASAP7_75t_L g10839 ( 
.A(n_9885),
.Y(n_10839)
);

INVx2_ASAP7_75t_L g10840 ( 
.A(n_10238),
.Y(n_10840)
);

NAND2xp5_ASAP7_75t_SL g10841 ( 
.A(n_9881),
.B(n_130),
.Y(n_10841)
);

INVxp67_ASAP7_75t_L g10842 ( 
.A(n_9967),
.Y(n_10842)
);

AND2x2_ASAP7_75t_L g10843 ( 
.A(n_10318),
.B(n_131),
.Y(n_10843)
);

INVx5_ASAP7_75t_L g10844 ( 
.A(n_10266),
.Y(n_10844)
);

AND2x2_ASAP7_75t_L g10845 ( 
.A(n_10014),
.B(n_131),
.Y(n_10845)
);

NAND2xp5_ASAP7_75t_L g10846 ( 
.A(n_10091),
.B(n_132),
.Y(n_10846)
);

INVx2_ASAP7_75t_L g10847 ( 
.A(n_10325),
.Y(n_10847)
);

INVx2_ASAP7_75t_L g10848 ( 
.A(n_10021),
.Y(n_10848)
);

HB1xp67_ASAP7_75t_L g10849 ( 
.A(n_10045),
.Y(n_10849)
);

OAI21xp5_ASAP7_75t_L g10850 ( 
.A1(n_10331),
.A2(n_132),
.B(n_133),
.Y(n_10850)
);

INVx1_ASAP7_75t_L g10851 ( 
.A(n_10202),
.Y(n_10851)
);

INVx2_ASAP7_75t_L g10852 ( 
.A(n_10094),
.Y(n_10852)
);

AND2x2_ASAP7_75t_SL g10853 ( 
.A(n_10107),
.B(n_133),
.Y(n_10853)
);

HB1xp67_ASAP7_75t_L g10854 ( 
.A(n_10315),
.Y(n_10854)
);

INVx1_ASAP7_75t_L g10855 ( 
.A(n_10110),
.Y(n_10855)
);

INVx2_ASAP7_75t_L g10856 ( 
.A(n_10284),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_10292),
.Y(n_10857)
);

AND2x2_ASAP7_75t_L g10858 ( 
.A(n_10005),
.B(n_134),
.Y(n_10858)
);

AND2x4_ASAP7_75t_L g10859 ( 
.A(n_9873),
.B(n_4647),
.Y(n_10859)
);

INVx1_ASAP7_75t_L g10860 ( 
.A(n_9830),
.Y(n_10860)
);

NAND2xp5_ASAP7_75t_SL g10861 ( 
.A(n_9868),
.B(n_134),
.Y(n_10861)
);

AND2x2_ASAP7_75t_L g10862 ( 
.A(n_10005),
.B(n_135),
.Y(n_10862)
);

AND2x4_ASAP7_75t_L g10863 ( 
.A(n_9873),
.B(n_4648),
.Y(n_10863)
);

AND2x2_ASAP7_75t_L g10864 ( 
.A(n_10005),
.B(n_135),
.Y(n_10864)
);

AND2x2_ASAP7_75t_L g10865 ( 
.A(n_10005),
.B(n_136),
.Y(n_10865)
);

INVx2_ASAP7_75t_SL g10866 ( 
.A(n_10054),
.Y(n_10866)
);

INVxp67_ASAP7_75t_SL g10867 ( 
.A(n_9870),
.Y(n_10867)
);

INVx3_ASAP7_75t_L g10868 ( 
.A(n_9848),
.Y(n_10868)
);

AND2x2_ASAP7_75t_L g10869 ( 
.A(n_10005),
.B(n_137),
.Y(n_10869)
);

INVx2_ASAP7_75t_L g10870 ( 
.A(n_9830),
.Y(n_10870)
);

AND2x4_ASAP7_75t_L g10871 ( 
.A(n_9873),
.B(n_4650),
.Y(n_10871)
);

AND2x2_ASAP7_75t_L g10872 ( 
.A(n_10005),
.B(n_137),
.Y(n_10872)
);

AND2x2_ASAP7_75t_L g10873 ( 
.A(n_10005),
.B(n_138),
.Y(n_10873)
);

NAND2xp5_ASAP7_75t_L g10874 ( 
.A(n_9868),
.B(n_138),
.Y(n_10874)
);

AND2x2_ASAP7_75t_L g10875 ( 
.A(n_10005),
.B(n_139),
.Y(n_10875)
);

INVx2_ASAP7_75t_SL g10876 ( 
.A(n_10054),
.Y(n_10876)
);

NOR2xp67_ASAP7_75t_L g10877 ( 
.A(n_9919),
.B(n_4651),
.Y(n_10877)
);

AND2x2_ASAP7_75t_L g10878 ( 
.A(n_10005),
.B(n_139),
.Y(n_10878)
);

INVx3_ASAP7_75t_L g10879 ( 
.A(n_9848),
.Y(n_10879)
);

BUFx4f_ASAP7_75t_L g10880 ( 
.A(n_9858),
.Y(n_10880)
);

AND2x2_ASAP7_75t_L g10881 ( 
.A(n_10005),
.B(n_140),
.Y(n_10881)
);

INVx4_ASAP7_75t_L g10882 ( 
.A(n_10112),
.Y(n_10882)
);

AND2x2_ASAP7_75t_L g10883 ( 
.A(n_10005),
.B(n_140),
.Y(n_10883)
);

AND2x6_ASAP7_75t_L g10884 ( 
.A(n_10207),
.B(n_4652),
.Y(n_10884)
);

AND2x2_ASAP7_75t_SL g10885 ( 
.A(n_9868),
.B(n_141),
.Y(n_10885)
);

AND2x2_ASAP7_75t_L g10886 ( 
.A(n_10005),
.B(n_141),
.Y(n_10886)
);

INVx1_ASAP7_75t_L g10887 ( 
.A(n_9830),
.Y(n_10887)
);

AND2x2_ASAP7_75t_L g10888 ( 
.A(n_10005),
.B(n_142),
.Y(n_10888)
);

BUFx2_ASAP7_75t_L g10889 ( 
.A(n_9870),
.Y(n_10889)
);

INVx2_ASAP7_75t_L g10890 ( 
.A(n_9830),
.Y(n_10890)
);

BUFx6f_ASAP7_75t_L g10891 ( 
.A(n_9858),
.Y(n_10891)
);

INVxp67_ASAP7_75t_L g10892 ( 
.A(n_9870),
.Y(n_10892)
);

AND2x2_ASAP7_75t_L g10893 ( 
.A(n_10005),
.B(n_142),
.Y(n_10893)
);

INVx3_ASAP7_75t_L g10894 ( 
.A(n_9848),
.Y(n_10894)
);

NOR2xp33_ASAP7_75t_SL g10895 ( 
.A(n_9919),
.B(n_4653),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_10005),
.B(n_143),
.Y(n_10896)
);

BUFx3_ASAP7_75t_L g10897 ( 
.A(n_10054),
.Y(n_10897)
);

OR2x2_ASAP7_75t_L g10898 ( 
.A(n_9878),
.B(n_143),
.Y(n_10898)
);

AND2x2_ASAP7_75t_L g10899 ( 
.A(n_10005),
.B(n_144),
.Y(n_10899)
);

NAND2xp5_ASAP7_75t_SL g10900 ( 
.A(n_9868),
.B(n_144),
.Y(n_10900)
);

INVx2_ASAP7_75t_L g10901 ( 
.A(n_9830),
.Y(n_10901)
);

NAND2xp5_ASAP7_75t_L g10902 ( 
.A(n_9868),
.B(n_145),
.Y(n_10902)
);

INVx1_ASAP7_75t_SL g10903 ( 
.A(n_9935),
.Y(n_10903)
);

INVx1_ASAP7_75t_L g10904 ( 
.A(n_9830),
.Y(n_10904)
);

NAND2xp5_ASAP7_75t_L g10905 ( 
.A(n_9868),
.B(n_145),
.Y(n_10905)
);

INVx2_ASAP7_75t_L g10906 ( 
.A(n_9830),
.Y(n_10906)
);

INVx2_ASAP7_75t_L g10907 ( 
.A(n_9830),
.Y(n_10907)
);

OAI21x1_ASAP7_75t_L g10908 ( 
.A1(n_9903),
.A2(n_4656),
.B(n_4654),
.Y(n_10908)
);

AND2x2_ASAP7_75t_L g10909 ( 
.A(n_10005),
.B(n_146),
.Y(n_10909)
);

INVx1_ASAP7_75t_L g10910 ( 
.A(n_9830),
.Y(n_10910)
);

AND2x2_ASAP7_75t_L g10911 ( 
.A(n_10005),
.B(n_146),
.Y(n_10911)
);

INVx1_ASAP7_75t_L g10912 ( 
.A(n_9830),
.Y(n_10912)
);

HB1xp67_ASAP7_75t_L g10913 ( 
.A(n_9870),
.Y(n_10913)
);

INVx2_ASAP7_75t_SL g10914 ( 
.A(n_10054),
.Y(n_10914)
);

AND2x2_ASAP7_75t_L g10915 ( 
.A(n_10005),
.B(n_147),
.Y(n_10915)
);

NAND2xp5_ASAP7_75t_L g10916 ( 
.A(n_9868),
.B(n_147),
.Y(n_10916)
);

OAI21xp5_ASAP7_75t_L g10917 ( 
.A1(n_9868),
.A2(n_148),
.B(n_149),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_9830),
.Y(n_10918)
);

AND2x2_ASAP7_75t_L g10919 ( 
.A(n_10005),
.B(n_148),
.Y(n_10919)
);

HB1xp67_ASAP7_75t_L g10920 ( 
.A(n_9870),
.Y(n_10920)
);

AND2x2_ASAP7_75t_SL g10921 ( 
.A(n_9868),
.B(n_149),
.Y(n_10921)
);

NAND2xp5_ASAP7_75t_L g10922 ( 
.A(n_9868),
.B(n_150),
.Y(n_10922)
);

HB1xp67_ASAP7_75t_L g10923 ( 
.A(n_9870),
.Y(n_10923)
);

AND2x2_ASAP7_75t_L g10924 ( 
.A(n_10005),
.B(n_150),
.Y(n_10924)
);

AND2x4_ASAP7_75t_L g10925 ( 
.A(n_9873),
.B(n_4658),
.Y(n_10925)
);

BUFx6f_ASAP7_75t_L g10926 ( 
.A(n_9858),
.Y(n_10926)
);

AND2x2_ASAP7_75t_L g10927 ( 
.A(n_10005),
.B(n_151),
.Y(n_10927)
);

BUFx4f_ASAP7_75t_L g10928 ( 
.A(n_9858),
.Y(n_10928)
);

AND2x2_ASAP7_75t_L g10929 ( 
.A(n_10005),
.B(n_152),
.Y(n_10929)
);

NAND2xp5_ASAP7_75t_L g10930 ( 
.A(n_9868),
.B(n_152),
.Y(n_10930)
);

CKINVDCx5p33_ASAP7_75t_R g10931 ( 
.A(n_9919),
.Y(n_10931)
);

NAND2xp5_ASAP7_75t_SL g10932 ( 
.A(n_9868),
.B(n_153),
.Y(n_10932)
);

NAND2xp5_ASAP7_75t_SL g10933 ( 
.A(n_9868),
.B(n_154),
.Y(n_10933)
);

INVx2_ASAP7_75t_L g10934 ( 
.A(n_9830),
.Y(n_10934)
);

INVx6_ASAP7_75t_L g10935 ( 
.A(n_10112),
.Y(n_10935)
);

NAND2xp5_ASAP7_75t_L g10936 ( 
.A(n_9868),
.B(n_154),
.Y(n_10936)
);

AND2x2_ASAP7_75t_L g10937 ( 
.A(n_10005),
.B(n_155),
.Y(n_10937)
);

AND2x2_ASAP7_75t_L g10938 ( 
.A(n_10005),
.B(n_155),
.Y(n_10938)
);

AND2x2_ASAP7_75t_L g10939 ( 
.A(n_10005),
.B(n_156),
.Y(n_10939)
);

INVx1_ASAP7_75t_SL g10940 ( 
.A(n_9935),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_9830),
.Y(n_10941)
);

AND2x4_ASAP7_75t_L g10942 ( 
.A(n_9873),
.B(n_4660),
.Y(n_10942)
);

INVx1_ASAP7_75t_L g10943 ( 
.A(n_9830),
.Y(n_10943)
);

INVx1_ASAP7_75t_L g10944 ( 
.A(n_9830),
.Y(n_10944)
);

NAND2xp5_ASAP7_75t_L g10945 ( 
.A(n_9868),
.B(n_157),
.Y(n_10945)
);

NAND2xp5_ASAP7_75t_L g10946 ( 
.A(n_9868),
.B(n_157),
.Y(n_10946)
);

INVx1_ASAP7_75t_L g10947 ( 
.A(n_9830),
.Y(n_10947)
);

INVx1_ASAP7_75t_L g10948 ( 
.A(n_9830),
.Y(n_10948)
);

BUFx3_ASAP7_75t_L g10949 ( 
.A(n_10054),
.Y(n_10949)
);

BUFx3_ASAP7_75t_L g10950 ( 
.A(n_10054),
.Y(n_10950)
);

INVx2_ASAP7_75t_L g10951 ( 
.A(n_9830),
.Y(n_10951)
);

NAND2xp5_ASAP7_75t_L g10952 ( 
.A(n_9868),
.B(n_158),
.Y(n_10952)
);

INVx1_ASAP7_75t_L g10953 ( 
.A(n_9830),
.Y(n_10953)
);

OR2x2_ASAP7_75t_L g10954 ( 
.A(n_9878),
.B(n_158),
.Y(n_10954)
);

AND2x2_ASAP7_75t_SL g10955 ( 
.A(n_9868),
.B(n_159),
.Y(n_10955)
);

AND2x2_ASAP7_75t_L g10956 ( 
.A(n_10005),
.B(n_159),
.Y(n_10956)
);

AND2x2_ASAP7_75t_L g10957 ( 
.A(n_10005),
.B(n_160),
.Y(n_10957)
);

NAND2xp5_ASAP7_75t_L g10958 ( 
.A(n_9868),
.B(n_160),
.Y(n_10958)
);

AND2x2_ASAP7_75t_L g10959 ( 
.A(n_10005),
.B(n_161),
.Y(n_10959)
);

BUFx3_ASAP7_75t_L g10960 ( 
.A(n_10054),
.Y(n_10960)
);

NAND2xp5_ASAP7_75t_L g10961 ( 
.A(n_9868),
.B(n_161),
.Y(n_10961)
);

INVx1_ASAP7_75t_L g10962 ( 
.A(n_9830),
.Y(n_10962)
);

NOR2xp33_ASAP7_75t_L g10963 ( 
.A(n_9868),
.B(n_4661),
.Y(n_10963)
);

AND2x2_ASAP7_75t_L g10964 ( 
.A(n_10005),
.B(n_162),
.Y(n_10964)
);

AND2x2_ASAP7_75t_L g10965 ( 
.A(n_10005),
.B(n_163),
.Y(n_10965)
);

INVx2_ASAP7_75t_L g10966 ( 
.A(n_9830),
.Y(n_10966)
);

AOI21xp5_ASAP7_75t_L g10967 ( 
.A1(n_10590),
.A2(n_4663),
.B(n_4662),
.Y(n_10967)
);

OR2x6_ASAP7_75t_L g10968 ( 
.A(n_10574),
.B(n_4666),
.Y(n_10968)
);

BUFx4f_ASAP7_75t_L g10969 ( 
.A(n_10393),
.Y(n_10969)
);

AOI21xp5_ASAP7_75t_L g10970 ( 
.A1(n_10472),
.A2(n_4669),
.B(n_4667),
.Y(n_10970)
);

NOR2xp33_ASAP7_75t_L g10971 ( 
.A(n_10592),
.B(n_10516),
.Y(n_10971)
);

NAND2xp5_ASAP7_75t_SL g10972 ( 
.A(n_10768),
.B(n_4670),
.Y(n_10972)
);

O2A1O1Ixp33_ASAP7_75t_L g10973 ( 
.A1(n_10535),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_10973)
);

AOI21xp5_ASAP7_75t_L g10974 ( 
.A1(n_10857),
.A2(n_4672),
.B(n_4671),
.Y(n_10974)
);

NOR2xp67_ASAP7_75t_L g10975 ( 
.A(n_10593),
.B(n_4673),
.Y(n_10975)
);

NAND2xp5_ASAP7_75t_L g10976 ( 
.A(n_10360),
.B(n_164),
.Y(n_10976)
);

AOI21xp5_ASAP7_75t_L g10977 ( 
.A1(n_10850),
.A2(n_4675),
.B(n_4674),
.Y(n_10977)
);

AOI21xp5_ASAP7_75t_L g10978 ( 
.A1(n_10829),
.A2(n_10798),
.B(n_10530),
.Y(n_10978)
);

OAI21xp5_ASAP7_75t_L g10979 ( 
.A1(n_10677),
.A2(n_165),
.B(n_167),
.Y(n_10979)
);

NAND2xp5_ASAP7_75t_L g10980 ( 
.A(n_10818),
.B(n_167),
.Y(n_10980)
);

INVx4_ASAP7_75t_L g10981 ( 
.A(n_10880),
.Y(n_10981)
);

OAI21xp5_ASAP7_75t_L g10982 ( 
.A1(n_10349),
.A2(n_168),
.B(n_169),
.Y(n_10982)
);

NOR2xp33_ASAP7_75t_L g10983 ( 
.A(n_10679),
.B(n_4677),
.Y(n_10983)
);

OAI21xp5_ASAP7_75t_L g10984 ( 
.A1(n_10469),
.A2(n_169),
.B(n_170),
.Y(n_10984)
);

AOI21xp5_ASAP7_75t_L g10985 ( 
.A1(n_10747),
.A2(n_4679),
.B(n_4678),
.Y(n_10985)
);

O2A1O1Ixp5_ASAP7_75t_L g10986 ( 
.A1(n_10660),
.A2(n_10667),
.B(n_10623),
.C(n_10646),
.Y(n_10986)
);

INVx2_ASAP7_75t_L g10987 ( 
.A(n_10345),
.Y(n_10987)
);

AOI21xp5_ASAP7_75t_L g10988 ( 
.A1(n_10347),
.A2(n_4682),
.B(n_4681),
.Y(n_10988)
);

INVx2_ASAP7_75t_L g10989 ( 
.A(n_10354),
.Y(n_10989)
);

NAND2xp5_ASAP7_75t_L g10990 ( 
.A(n_10659),
.B(n_10663),
.Y(n_10990)
);

NAND3xp33_ASAP7_75t_L g10991 ( 
.A(n_10745),
.B(n_170),
.C(n_171),
.Y(n_10991)
);

AOI21xp5_ASAP7_75t_L g10992 ( 
.A1(n_10838),
.A2(n_4684),
.B(n_4683),
.Y(n_10992)
);

NAND2xp5_ASAP7_75t_L g10993 ( 
.A(n_10665),
.B(n_171),
.Y(n_10993)
);

AOI21xp5_ASAP7_75t_L g10994 ( 
.A1(n_10690),
.A2(n_4686),
.B(n_4685),
.Y(n_10994)
);

AOI21xp5_ASAP7_75t_L g10995 ( 
.A1(n_10685),
.A2(n_4688),
.B(n_4687),
.Y(n_10995)
);

INVx1_ASAP7_75t_L g10996 ( 
.A(n_10641),
.Y(n_10996)
);

OAI22xp5_ASAP7_75t_L g10997 ( 
.A1(n_10724),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_10997)
);

INVx1_ASAP7_75t_L g10998 ( 
.A(n_10654),
.Y(n_10998)
);

INVx1_ASAP7_75t_L g10999 ( 
.A(n_10429),
.Y(n_10999)
);

NOR3xp33_ASAP7_75t_L g11000 ( 
.A(n_10703),
.B(n_10708),
.C(n_10689),
.Y(n_11000)
);

AOI21xp5_ASAP7_75t_L g11001 ( 
.A1(n_10691),
.A2(n_4690),
.B(n_4689),
.Y(n_11001)
);

OAI22xp5_ASAP7_75t_L g11002 ( 
.A1(n_10397),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_11002)
);

NAND2xp5_ASAP7_75t_L g11003 ( 
.A(n_10666),
.B(n_176),
.Y(n_11003)
);

INVxp67_ASAP7_75t_L g11004 ( 
.A(n_10913),
.Y(n_11004)
);

AOI21xp5_ASAP7_75t_L g11005 ( 
.A1(n_10728),
.A2(n_10409),
.B(n_10404),
.Y(n_11005)
);

AOI21xp5_ASAP7_75t_L g11006 ( 
.A1(n_10403),
.A2(n_4694),
.B(n_4691),
.Y(n_11006)
);

INVx1_ASAP7_75t_L g11007 ( 
.A(n_10434),
.Y(n_11007)
);

AOI21xp5_ASAP7_75t_L g11008 ( 
.A1(n_10963),
.A2(n_4697),
.B(n_4695),
.Y(n_11008)
);

AO22x1_ASAP7_75t_L g11009 ( 
.A1(n_10511),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_11009)
);

AOI21xp5_ASAP7_75t_L g11010 ( 
.A1(n_10735),
.A2(n_4703),
.B(n_4699),
.Y(n_11010)
);

AOI21xp5_ASAP7_75t_L g11011 ( 
.A1(n_10855),
.A2(n_4705),
.B(n_4704),
.Y(n_11011)
);

BUFx6f_ASAP7_75t_L g11012 ( 
.A(n_10928),
.Y(n_11012)
);

NAND2xp5_ASAP7_75t_L g11013 ( 
.A(n_10671),
.B(n_177),
.Y(n_11013)
);

AND2x2_ASAP7_75t_L g11014 ( 
.A(n_10815),
.B(n_4706),
.Y(n_11014)
);

AND2x2_ASAP7_75t_L g11015 ( 
.A(n_10447),
.B(n_4707),
.Y(n_11015)
);

NAND2xp5_ASAP7_75t_L g11016 ( 
.A(n_10674),
.B(n_178),
.Y(n_11016)
);

INVx2_ASAP7_75t_L g11017 ( 
.A(n_10356),
.Y(n_11017)
);

BUFx12f_ASAP7_75t_L g11018 ( 
.A(n_10518),
.Y(n_11018)
);

OAI321xp33_ASAP7_75t_L g11019 ( 
.A1(n_10346),
.A2(n_181),
.A3(n_183),
.B1(n_179),
.B2(n_180),
.C(n_182),
.Y(n_11019)
);

OAI22xp5_ASAP7_75t_L g11020 ( 
.A1(n_10823),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_11020)
);

OAI21xp5_ASAP7_75t_L g11021 ( 
.A1(n_10830),
.A2(n_183),
.B(n_184),
.Y(n_11021)
);

OR2x2_ASAP7_75t_L g11022 ( 
.A(n_10462),
.B(n_184),
.Y(n_11022)
);

OAI21xp5_ASAP7_75t_L g11023 ( 
.A1(n_10449),
.A2(n_185),
.B(n_186),
.Y(n_11023)
);

INVx1_ASAP7_75t_L g11024 ( 
.A(n_10455),
.Y(n_11024)
);

BUFx6f_ASAP7_75t_L g11025 ( 
.A(n_10897),
.Y(n_11025)
);

NOR2xp33_ASAP7_75t_L g11026 ( 
.A(n_10687),
.B(n_4711),
.Y(n_11026)
);

AOI21xp5_ASAP7_75t_L g11027 ( 
.A1(n_10636),
.A2(n_4715),
.B(n_4714),
.Y(n_11027)
);

AOI21xp5_ASAP7_75t_L g11028 ( 
.A1(n_10917),
.A2(n_4718),
.B(n_4717),
.Y(n_11028)
);

OAI21xp5_ASAP7_75t_L g11029 ( 
.A1(n_10624),
.A2(n_185),
.B(n_186),
.Y(n_11029)
);

AOI21xp5_ASAP7_75t_L g11030 ( 
.A1(n_10766),
.A2(n_4720),
.B(n_4719),
.Y(n_11030)
);

OR2x6_ASAP7_75t_L g11031 ( 
.A(n_10574),
.B(n_4721),
.Y(n_11031)
);

HB1xp67_ASAP7_75t_L g11032 ( 
.A(n_10920),
.Y(n_11032)
);

NAND2xp5_ASAP7_75t_L g11033 ( 
.A(n_10694),
.B(n_187),
.Y(n_11033)
);

NAND2xp5_ASAP7_75t_L g11034 ( 
.A(n_10696),
.B(n_187),
.Y(n_11034)
);

INVx1_ASAP7_75t_L g11035 ( 
.A(n_10470),
.Y(n_11035)
);

BUFx6f_ASAP7_75t_L g11036 ( 
.A(n_10949),
.Y(n_11036)
);

HB1xp67_ASAP7_75t_L g11037 ( 
.A(n_10923),
.Y(n_11037)
);

NOR2xp33_ASAP7_75t_L g11038 ( 
.A(n_10389),
.B(n_4722),
.Y(n_11038)
);

O2A1O1Ixp33_ASAP7_75t_L g11039 ( 
.A1(n_10833),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_11039)
);

NAND2xp5_ASAP7_75t_L g11040 ( 
.A(n_10784),
.B(n_188),
.Y(n_11040)
);

INVx1_ASAP7_75t_L g11041 ( 
.A(n_10476),
.Y(n_11041)
);

NAND3xp33_ASAP7_75t_L g11042 ( 
.A(n_10580),
.B(n_189),
.C(n_190),
.Y(n_11042)
);

A2O1A1Ixp33_ASAP7_75t_L g11043 ( 
.A1(n_10570),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_11043)
);

A2O1A1Ixp33_ASAP7_75t_L g11044 ( 
.A1(n_10835),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_11044)
);

NAND2xp5_ASAP7_75t_L g11045 ( 
.A(n_10793),
.B(n_194),
.Y(n_11045)
);

NOR3xp33_ASAP7_75t_L g11046 ( 
.A(n_10715),
.B(n_195),
.C(n_196),
.Y(n_11046)
);

OAI21xp5_ASAP7_75t_L g11047 ( 
.A1(n_10762),
.A2(n_196),
.B(n_197),
.Y(n_11047)
);

AOI21xp5_ASAP7_75t_L g11048 ( 
.A1(n_10785),
.A2(n_4724),
.B(n_4723),
.Y(n_11048)
);

NAND2xp5_ASAP7_75t_L g11049 ( 
.A(n_10797),
.B(n_197),
.Y(n_11049)
);

O2A1O1Ixp33_ASAP7_75t_L g11050 ( 
.A1(n_10700),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_11050)
);

NAND2xp5_ASAP7_75t_SL g11051 ( 
.A(n_10755),
.B(n_10761),
.Y(n_11051)
);

INVx1_ASAP7_75t_L g11052 ( 
.A(n_10485),
.Y(n_11052)
);

INVx3_ASAP7_75t_L g11053 ( 
.A(n_10502),
.Y(n_11053)
);

AND2x2_ASAP7_75t_L g11054 ( 
.A(n_10452),
.B(n_4728),
.Y(n_11054)
);

INVx3_ASAP7_75t_L g11055 ( 
.A(n_10344),
.Y(n_11055)
);

NOR2xp33_ASAP7_75t_L g11056 ( 
.A(n_10562),
.B(n_4729),
.Y(n_11056)
);

INVx2_ASAP7_75t_L g11057 ( 
.A(n_10357),
.Y(n_11057)
);

NAND2xp5_ASAP7_75t_L g11058 ( 
.A(n_10771),
.B(n_198),
.Y(n_11058)
);

OAI21xp33_ASAP7_75t_L g11059 ( 
.A1(n_10417),
.A2(n_200),
.B(n_201),
.Y(n_11059)
);

AOI21xp5_ASAP7_75t_L g11060 ( 
.A1(n_10770),
.A2(n_10779),
.B(n_10528),
.Y(n_11060)
);

NAND2xp5_ASAP7_75t_L g11061 ( 
.A(n_10697),
.B(n_201),
.Y(n_11061)
);

AOI21x1_ASAP7_75t_L g11062 ( 
.A1(n_10811),
.A2(n_10824),
.B(n_10804),
.Y(n_11062)
);

AOI21xp5_ASAP7_75t_L g11063 ( 
.A1(n_10725),
.A2(n_4731),
.B(n_4730),
.Y(n_11063)
);

NOR2x1_ASAP7_75t_L g11064 ( 
.A(n_10819),
.B(n_202),
.Y(n_11064)
);

AOI21xp5_ASAP7_75t_L g11065 ( 
.A1(n_10733),
.A2(n_4733),
.B(n_4732),
.Y(n_11065)
);

NOR2xp33_ASAP7_75t_L g11066 ( 
.A(n_10639),
.B(n_10602),
.Y(n_11066)
);

AOI21x1_ASAP7_75t_L g11067 ( 
.A1(n_10809),
.A2(n_4736),
.B(n_4735),
.Y(n_11067)
);

AOI21xp5_ASAP7_75t_L g11068 ( 
.A1(n_10740),
.A2(n_4738),
.B(n_4737),
.Y(n_11068)
);

OAI22xp5_ASAP7_75t_L g11069 ( 
.A1(n_10381),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_11069)
);

AO22x1_ASAP7_75t_L g11070 ( 
.A1(n_10511),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_11070)
);

NAND2xp5_ASAP7_75t_L g11071 ( 
.A(n_10746),
.B(n_10748),
.Y(n_11071)
);

A2O1A1Ixp33_ASAP7_75t_L g11072 ( 
.A1(n_10575),
.A2(n_208),
.B(n_205),
.C(n_207),
.Y(n_11072)
);

O2A1O1Ixp33_ASAP7_75t_L g11073 ( 
.A1(n_10705),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_11073)
);

INVx2_ASAP7_75t_L g11074 ( 
.A(n_10366),
.Y(n_11074)
);

OAI22xp5_ASAP7_75t_L g11075 ( 
.A1(n_10370),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_11075)
);

OAI22xp5_ASAP7_75t_L g11076 ( 
.A1(n_10831),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_11076)
);

NAND2xp5_ASAP7_75t_L g11077 ( 
.A(n_10757),
.B(n_213),
.Y(n_11077)
);

AOI22xp5_ASAP7_75t_L g11078 ( 
.A1(n_10511),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_11078)
);

NOR2xp33_ASAP7_75t_SL g11079 ( 
.A(n_10479),
.B(n_4741),
.Y(n_11079)
);

AND2x6_ASAP7_75t_SL g11080 ( 
.A(n_10816),
.B(n_214),
.Y(n_11080)
);

AOI22xp5_ASAP7_75t_L g11081 ( 
.A1(n_10669),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_11081)
);

AOI21xp5_ASAP7_75t_L g11082 ( 
.A1(n_10772),
.A2(n_4743),
.B(n_4742),
.Y(n_11082)
);

NAND2xp5_ASAP7_75t_L g11083 ( 
.A(n_10773),
.B(n_217),
.Y(n_11083)
);

AOI21xp5_ASAP7_75t_L g11084 ( 
.A1(n_10777),
.A2(n_4745),
.B(n_4744),
.Y(n_11084)
);

NAND2xp5_ASAP7_75t_SL g11085 ( 
.A(n_10606),
.B(n_4746),
.Y(n_11085)
);

NOR2x1_ASAP7_75t_L g11086 ( 
.A(n_10702),
.B(n_218),
.Y(n_11086)
);

AOI21xp5_ASAP7_75t_L g11087 ( 
.A1(n_10778),
.A2(n_4748),
.B(n_4747),
.Y(n_11087)
);

NOR2x1_ASAP7_75t_L g11088 ( 
.A(n_10680),
.B(n_218),
.Y(n_11088)
);

O2A1O1Ixp5_ASAP7_75t_L g11089 ( 
.A1(n_10398),
.A2(n_10711),
.B(n_10900),
.C(n_10861),
.Y(n_11089)
);

AOI21x1_ASAP7_75t_L g11090 ( 
.A1(n_10822),
.A2(n_4750),
.B(n_4749),
.Y(n_11090)
);

NAND2xp5_ASAP7_75t_L g11091 ( 
.A(n_10707),
.B(n_10658),
.Y(n_11091)
);

AOI21xp5_ASAP7_75t_L g11092 ( 
.A1(n_10372),
.A2(n_4753),
.B(n_4752),
.Y(n_11092)
);

A2O1A1Ixp33_ASAP7_75t_L g11093 ( 
.A1(n_10718),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_11093)
);

NOR2xp33_ASAP7_75t_L g11094 ( 
.A(n_10615),
.B(n_4754),
.Y(n_11094)
);

O2A1O1Ixp33_ASAP7_75t_L g11095 ( 
.A1(n_10527),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_10493),
.Y(n_11096)
);

NAND2xp5_ASAP7_75t_L g11097 ( 
.A(n_10392),
.B(n_222),
.Y(n_11097)
);

AOI21xp5_ASAP7_75t_L g11098 ( 
.A1(n_10682),
.A2(n_4757),
.B(n_4755),
.Y(n_11098)
);

AOI21xp5_ASAP7_75t_L g11099 ( 
.A1(n_10841),
.A2(n_4760),
.B(n_4759),
.Y(n_11099)
);

OR2x2_ASAP7_75t_L g11100 ( 
.A(n_10867),
.B(n_222),
.Y(n_11100)
);

AOI21xp5_ASAP7_75t_L g11101 ( 
.A1(n_10810),
.A2(n_4764),
.B(n_4763),
.Y(n_11101)
);

NOR2xp33_ASAP7_75t_L g11102 ( 
.A(n_10565),
.B(n_4765),
.Y(n_11102)
);

NAND2xp5_ASAP7_75t_L g11103 ( 
.A(n_10889),
.B(n_223),
.Y(n_11103)
);

AOI22xp5_ASAP7_75t_L g11104 ( 
.A1(n_10614),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_11104)
);

NAND2xp5_ASAP7_75t_L g11105 ( 
.A(n_10433),
.B(n_224),
.Y(n_11105)
);

AOI21xp5_ASAP7_75t_L g11106 ( 
.A1(n_10668),
.A2(n_4767),
.B(n_4766),
.Y(n_11106)
);

OR2x2_ASAP7_75t_L g11107 ( 
.A(n_10503),
.B(n_225),
.Y(n_11107)
);

NAND2xp5_ASAP7_75t_L g11108 ( 
.A(n_10628),
.B(n_226),
.Y(n_11108)
);

OAI21xp33_ASAP7_75t_SL g11109 ( 
.A1(n_10853),
.A2(n_227),
.B(n_228),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_10377),
.Y(n_11110)
);

AOI21xp5_ASAP7_75t_L g11111 ( 
.A1(n_10670),
.A2(n_4771),
.B(n_4769),
.Y(n_11111)
);

INVx1_ASAP7_75t_L g11112 ( 
.A(n_10494),
.Y(n_11112)
);

A2O1A1Ixp33_ASAP7_75t_L g11113 ( 
.A1(n_10851),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_11113)
);

NAND2xp5_ASAP7_75t_L g11114 ( 
.A(n_10400),
.B(n_230),
.Y(n_11114)
);

INVx4_ASAP7_75t_L g11115 ( 
.A(n_10950),
.Y(n_11115)
);

AO21x1_ASAP7_75t_L g11116 ( 
.A1(n_10932),
.A2(n_230),
.B(n_231),
.Y(n_11116)
);

NAND2xp5_ASAP7_75t_L g11117 ( 
.A(n_10634),
.B(n_231),
.Y(n_11117)
);

INVx3_ASAP7_75t_L g11118 ( 
.A(n_10448),
.Y(n_11118)
);

NAND3xp33_ASAP7_75t_L g11119 ( 
.A(n_10364),
.B(n_232),
.C(n_233),
.Y(n_11119)
);

AOI21x1_ASAP7_75t_L g11120 ( 
.A1(n_10908),
.A2(n_4773),
.B(n_4772),
.Y(n_11120)
);

O2A1O1Ixp33_ASAP7_75t_L g11121 ( 
.A1(n_10933),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_11121)
);

INVx11_ASAP7_75t_L g11122 ( 
.A(n_10673),
.Y(n_11122)
);

INVx1_ASAP7_75t_L g11123 ( 
.A(n_10498),
.Y(n_11123)
);

OAI22xp5_ASAP7_75t_L g11124 ( 
.A1(n_10780),
.A2(n_10491),
.B1(n_10749),
.B2(n_10847),
.Y(n_11124)
);

AOI21x1_ASAP7_75t_L g11125 ( 
.A1(n_10756),
.A2(n_4777),
.B(n_4775),
.Y(n_11125)
);

OAI21xp5_ASAP7_75t_L g11126 ( 
.A1(n_10723),
.A2(n_234),
.B(n_235),
.Y(n_11126)
);

AOI21xp5_ASAP7_75t_L g11127 ( 
.A1(n_10672),
.A2(n_4779),
.B(n_4778),
.Y(n_11127)
);

NOR3xp33_ASAP7_75t_L g11128 ( 
.A(n_10681),
.B(n_236),
.C(n_237),
.Y(n_11128)
);

INVx3_ASAP7_75t_L g11129 ( 
.A(n_10960),
.Y(n_11129)
);

BUFx6f_ASAP7_75t_L g11130 ( 
.A(n_10393),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_SL g11131 ( 
.A(n_10786),
.B(n_4780),
.Y(n_11131)
);

INVx1_ASAP7_75t_L g11132 ( 
.A(n_10531),
.Y(n_11132)
);

AOI21xp5_ASAP7_75t_L g11133 ( 
.A1(n_10688),
.A2(n_4782),
.B(n_4781),
.Y(n_11133)
);

INVx1_ASAP7_75t_L g11134 ( 
.A(n_10542),
.Y(n_11134)
);

AOI21xp5_ASAP7_75t_L g11135 ( 
.A1(n_10699),
.A2(n_4785),
.B(n_4783),
.Y(n_11135)
);

A2O1A1Ixp33_ASAP7_75t_L g11136 ( 
.A1(n_10806),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_11136)
);

AOI21xp5_ASAP7_75t_L g11137 ( 
.A1(n_10712),
.A2(n_4788),
.B(n_4786),
.Y(n_11137)
);

AOI21xp5_ASAP7_75t_L g11138 ( 
.A1(n_10719),
.A2(n_4790),
.B(n_4789),
.Y(n_11138)
);

NAND2xp5_ASAP7_75t_L g11139 ( 
.A(n_10425),
.B(n_10477),
.Y(n_11139)
);

NAND2xp5_ASAP7_75t_SL g11140 ( 
.A(n_10805),
.B(n_4792),
.Y(n_11140)
);

NAND2xp5_ASAP7_75t_SL g11141 ( 
.A(n_10844),
.B(n_4795),
.Y(n_11141)
);

AOI21xp5_ASAP7_75t_L g11142 ( 
.A1(n_10742),
.A2(n_4799),
.B(n_4797),
.Y(n_11142)
);

INVx2_ASAP7_75t_L g11143 ( 
.A(n_10380),
.Y(n_11143)
);

AND2x2_ASAP7_75t_L g11144 ( 
.A(n_10507),
.B(n_4800),
.Y(n_11144)
);

AOI21xp5_ASAP7_75t_L g11145 ( 
.A1(n_10828),
.A2(n_4802),
.B(n_4801),
.Y(n_11145)
);

BUFx4f_ASAP7_75t_L g11146 ( 
.A(n_10424),
.Y(n_11146)
);

NAND2x1p5_ASAP7_75t_L g11147 ( 
.A(n_10520),
.B(n_4803),
.Y(n_11147)
);

NAND2xp33_ASAP7_75t_L g11148 ( 
.A(n_10759),
.B(n_239),
.Y(n_11148)
);

NOR2xp33_ASAP7_75t_L g11149 ( 
.A(n_10376),
.B(n_4804),
.Y(n_11149)
);

NAND2xp5_ASAP7_75t_L g11150 ( 
.A(n_10355),
.B(n_239),
.Y(n_11150)
);

AOI21xp5_ASAP7_75t_L g11151 ( 
.A1(n_10832),
.A2(n_4808),
.B(n_4805),
.Y(n_11151)
);

NAND3xp33_ASAP7_75t_L g11152 ( 
.A(n_10729),
.B(n_240),
.C(n_241),
.Y(n_11152)
);

AOI21xp5_ASAP7_75t_L g11153 ( 
.A1(n_10895),
.A2(n_4810),
.B(n_4809),
.Y(n_11153)
);

INVx2_ASAP7_75t_L g11154 ( 
.A(n_10386),
.Y(n_11154)
);

AOI21xp5_ASAP7_75t_L g11155 ( 
.A1(n_10776),
.A2(n_4812),
.B(n_4811),
.Y(n_11155)
);

INVx3_ASAP7_75t_L g11156 ( 
.A(n_10423),
.Y(n_11156)
);

NAND2xp5_ASAP7_75t_L g11157 ( 
.A(n_10892),
.B(n_240),
.Y(n_11157)
);

NAND2xp5_ASAP7_75t_L g11158 ( 
.A(n_10428),
.B(n_241),
.Y(n_11158)
);

AOI21xp5_ASAP7_75t_L g11159 ( 
.A1(n_10788),
.A2(n_4814),
.B(n_4813),
.Y(n_11159)
);

NAND3xp33_ASAP7_75t_L g11160 ( 
.A(n_10846),
.B(n_242),
.C(n_243),
.Y(n_11160)
);

OAI22xp5_ASAP7_75t_L g11161 ( 
.A1(n_10795),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_11161)
);

OAI21xp5_ASAP7_75t_L g11162 ( 
.A1(n_10533),
.A2(n_244),
.B(n_245),
.Y(n_11162)
);

AOI21xp5_ASAP7_75t_L g11163 ( 
.A1(n_10767),
.A2(n_4817),
.B(n_4815),
.Y(n_11163)
);

INVx1_ASAP7_75t_L g11164 ( 
.A(n_10564),
.Y(n_11164)
);

AOI21xp5_ASAP7_75t_L g11165 ( 
.A1(n_10616),
.A2(n_4819),
.B(n_4818),
.Y(n_11165)
);

AOI21xp5_ASAP7_75t_L g11166 ( 
.A1(n_10714),
.A2(n_4821),
.B(n_4820),
.Y(n_11166)
);

OAI21xp5_ASAP7_75t_L g11167 ( 
.A1(n_10537),
.A2(n_246),
.B(n_247),
.Y(n_11167)
);

NOR2xp33_ASAP7_75t_L g11168 ( 
.A(n_10903),
.B(n_4822),
.Y(n_11168)
);

BUFx4f_ASAP7_75t_L g11169 ( 
.A(n_10424),
.Y(n_11169)
);

INVx1_ASAP7_75t_L g11170 ( 
.A(n_10581),
.Y(n_11170)
);

INVx4_ASAP7_75t_L g11171 ( 
.A(n_10891),
.Y(n_11171)
);

AOI21xp5_ASAP7_75t_L g11172 ( 
.A1(n_10840),
.A2(n_4824),
.B(n_4823),
.Y(n_11172)
);

BUFx6f_ASAP7_75t_L g11173 ( 
.A(n_10891),
.Y(n_11173)
);

NAND2xp5_ASAP7_75t_L g11174 ( 
.A(n_10394),
.B(n_246),
.Y(n_11174)
);

AOI21xp5_ASAP7_75t_L g11175 ( 
.A1(n_10856),
.A2(n_4827),
.B(n_4826),
.Y(n_11175)
);

AOI21xp5_ASAP7_75t_L g11176 ( 
.A1(n_10852),
.A2(n_4831),
.B(n_4828),
.Y(n_11176)
);

INVx1_ASAP7_75t_L g11177 ( 
.A(n_10586),
.Y(n_11177)
);

BUFx2_ASAP7_75t_L g11178 ( 
.A(n_10534),
.Y(n_11178)
);

OAI21xp33_ASAP7_75t_L g11179 ( 
.A1(n_10836),
.A2(n_247),
.B(n_248),
.Y(n_11179)
);

HB1xp67_ASAP7_75t_L g11180 ( 
.A(n_10550),
.Y(n_11180)
);

AOI21xp5_ASAP7_75t_L g11181 ( 
.A1(n_10657),
.A2(n_4834),
.B(n_4832),
.Y(n_11181)
);

INVx1_ASAP7_75t_L g11182 ( 
.A(n_10597),
.Y(n_11182)
);

INVx5_ASAP7_75t_L g11183 ( 
.A(n_10407),
.Y(n_11183)
);

INVx2_ASAP7_75t_L g11184 ( 
.A(n_10405),
.Y(n_11184)
);

INVx2_ASAP7_75t_L g11185 ( 
.A(n_10413),
.Y(n_11185)
);

A2O1A1Ixp33_ASAP7_75t_L g11186 ( 
.A1(n_10538),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_11186)
);

INVx3_ASAP7_75t_L g11187 ( 
.A(n_10545),
.Y(n_11187)
);

AOI21xp5_ASAP7_75t_L g11188 ( 
.A1(n_10808),
.A2(n_4836),
.B(n_4835),
.Y(n_11188)
);

NAND2x1p5_ASAP7_75t_L g11189 ( 
.A(n_10432),
.B(n_4837),
.Y(n_11189)
);

INVx2_ASAP7_75t_L g11190 ( 
.A(n_10870),
.Y(n_11190)
);

NOR2xp33_ASAP7_75t_L g11191 ( 
.A(n_10940),
.B(n_4838),
.Y(n_11191)
);

AOI21xp5_ASAP7_75t_L g11192 ( 
.A1(n_10812),
.A2(n_4840),
.B(n_4839),
.Y(n_11192)
);

OAI21xp5_ASAP7_75t_L g11193 ( 
.A1(n_10556),
.A2(n_249),
.B(n_250),
.Y(n_11193)
);

AND2x2_ASAP7_75t_SL g11194 ( 
.A(n_10885),
.B(n_251),
.Y(n_11194)
);

INVx2_ASAP7_75t_L g11195 ( 
.A(n_10890),
.Y(n_11195)
);

OAI21xp5_ASAP7_75t_L g11196 ( 
.A1(n_10561),
.A2(n_252),
.B(n_253),
.Y(n_11196)
);

CKINVDCx10_ASAP7_75t_R g11197 ( 
.A(n_10532),
.Y(n_11197)
);

BUFx6f_ASAP7_75t_L g11198 ( 
.A(n_10926),
.Y(n_11198)
);

AOI21xp5_ASAP7_75t_L g11199 ( 
.A1(n_10650),
.A2(n_4842),
.B(n_4841),
.Y(n_11199)
);

O2A1O1Ixp33_ASAP7_75t_SL g11200 ( 
.A1(n_10813),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_11200)
);

BUFx3_ASAP7_75t_L g11201 ( 
.A(n_10474),
.Y(n_11201)
);

HB1xp67_ASAP7_75t_L g11202 ( 
.A(n_10551),
.Y(n_11202)
);

NAND2xp5_ASAP7_75t_L g11203 ( 
.A(n_10901),
.B(n_254),
.Y(n_11203)
);

AOI21xp5_ASAP7_75t_L g11204 ( 
.A1(n_10652),
.A2(n_4844),
.B(n_4843),
.Y(n_11204)
);

INVx1_ASAP7_75t_L g11205 ( 
.A(n_10599),
.Y(n_11205)
);

HB1xp67_ASAP7_75t_L g11206 ( 
.A(n_10571),
.Y(n_11206)
);

AND2x4_ASAP7_75t_L g11207 ( 
.A(n_10601),
.B(n_4845),
.Y(n_11207)
);

NAND2xp5_ASAP7_75t_L g11208 ( 
.A(n_10906),
.B(n_255),
.Y(n_11208)
);

OAI22xp5_ASAP7_75t_L g11209 ( 
.A1(n_10548),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_11209)
);

NAND2xp5_ASAP7_75t_L g11210 ( 
.A(n_10907),
.B(n_256),
.Y(n_11210)
);

BUFx4f_ASAP7_75t_L g11211 ( 
.A(n_10926),
.Y(n_11211)
);

INVx1_ASAP7_75t_SL g11212 ( 
.A(n_10578),
.Y(n_11212)
);

AOI21xp5_ASAP7_75t_L g11213 ( 
.A1(n_10430),
.A2(n_4849),
.B(n_4846),
.Y(n_11213)
);

NAND2xp5_ASAP7_75t_L g11214 ( 
.A(n_10934),
.B(n_10951),
.Y(n_11214)
);

AO21x1_ASAP7_75t_L g11215 ( 
.A1(n_10439),
.A2(n_257),
.B(n_258),
.Y(n_11215)
);

NOR2xp33_ASAP7_75t_L g11216 ( 
.A(n_10727),
.B(n_10710),
.Y(n_11216)
);

INVx2_ASAP7_75t_L g11217 ( 
.A(n_10966),
.Y(n_11217)
);

BUFx12f_ASAP7_75t_L g11218 ( 
.A(n_10931),
.Y(n_11218)
);

AOI21xp5_ASAP7_75t_L g11219 ( 
.A1(n_10437),
.A2(n_4851),
.B(n_4850),
.Y(n_11219)
);

AO22x1_ASAP7_75t_L g11220 ( 
.A1(n_10517),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_11220)
);

INVx1_ASAP7_75t_L g11221 ( 
.A(n_10600),
.Y(n_11221)
);

INVx1_ASAP7_75t_L g11222 ( 
.A(n_10627),
.Y(n_11222)
);

O2A1O1Ixp33_ASAP7_75t_L g11223 ( 
.A1(n_10638),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_11223)
);

INVx5_ASAP7_75t_L g11224 ( 
.A(n_10407),
.Y(n_11224)
);

OAI21xp5_ASAP7_75t_L g11225 ( 
.A1(n_10572),
.A2(n_261),
.B(n_263),
.Y(n_11225)
);

NAND2xp5_ASAP7_75t_L g11226 ( 
.A(n_10607),
.B(n_263),
.Y(n_11226)
);

AOI21x1_ASAP7_75t_L g11227 ( 
.A1(n_10483),
.A2(n_4853),
.B(n_4852),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_10630),
.Y(n_11228)
);

NAND2xp5_ASAP7_75t_L g11229 ( 
.A(n_10401),
.B(n_264),
.Y(n_11229)
);

AOI21xp5_ASAP7_75t_L g11230 ( 
.A1(n_10445),
.A2(n_4855),
.B(n_4854),
.Y(n_11230)
);

INVx1_ASAP7_75t_L g11231 ( 
.A(n_10631),
.Y(n_11231)
);

AOI21x1_ASAP7_75t_L g11232 ( 
.A1(n_10350),
.A2(n_4857),
.B(n_4856),
.Y(n_11232)
);

AOI21xp5_ASAP7_75t_L g11233 ( 
.A1(n_10632),
.A2(n_4859),
.B(n_4858),
.Y(n_11233)
);

AOI21xp5_ASAP7_75t_L g11234 ( 
.A1(n_10651),
.A2(n_4862),
.B(n_4861),
.Y(n_11234)
);

BUFx3_ASAP7_75t_L g11235 ( 
.A(n_10459),
.Y(n_11235)
);

NAND2xp5_ASAP7_75t_L g11236 ( 
.A(n_10384),
.B(n_264),
.Y(n_11236)
);

OAI22xp5_ASAP7_75t_L g11237 ( 
.A1(n_10921),
.A2(n_10955),
.B1(n_10554),
.B2(n_10854),
.Y(n_11237)
);

AOI21xp5_ASAP7_75t_L g11238 ( 
.A1(n_10655),
.A2(n_4864),
.B(n_4863),
.Y(n_11238)
);

OAI21xp5_ASAP7_75t_L g11239 ( 
.A1(n_10576),
.A2(n_10604),
.B(n_10595),
.Y(n_11239)
);

O2A1O1Ixp33_ASAP7_75t_L g11240 ( 
.A1(n_10874),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_11240)
);

AOI21xp5_ASAP7_75t_L g11241 ( 
.A1(n_10361),
.A2(n_4866),
.B(n_4865),
.Y(n_11241)
);

NAND2xp5_ASAP7_75t_L g11242 ( 
.A(n_10390),
.B(n_265),
.Y(n_11242)
);

BUFx6f_ASAP7_75t_L g11243 ( 
.A(n_10352),
.Y(n_11243)
);

OAI21xp5_ASAP7_75t_L g11244 ( 
.A1(n_10605),
.A2(n_266),
.B(n_267),
.Y(n_11244)
);

NAND2xp5_ASAP7_75t_L g11245 ( 
.A(n_10396),
.B(n_268),
.Y(n_11245)
);

AND2x2_ASAP7_75t_L g11246 ( 
.A(n_10802),
.B(n_4867),
.Y(n_11246)
);

NAND2xp5_ASAP7_75t_L g11247 ( 
.A(n_10378),
.B(n_269),
.Y(n_11247)
);

OAI22xp5_ASAP7_75t_L g11248 ( 
.A1(n_10842),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_11248)
);

NAND2xp5_ASAP7_75t_L g11249 ( 
.A(n_10451),
.B(n_270),
.Y(n_11249)
);

INVx3_ASAP7_75t_L g11250 ( 
.A(n_10545),
.Y(n_11250)
);

NOR2xp33_ASAP7_75t_SL g11251 ( 
.A(n_10438),
.B(n_4868),
.Y(n_11251)
);

INVx1_ASAP7_75t_L g11252 ( 
.A(n_10522),
.Y(n_11252)
);

NOR2xp33_ASAP7_75t_L g11253 ( 
.A(n_10800),
.B(n_4869),
.Y(n_11253)
);

NOR3xp33_ASAP7_75t_L g11254 ( 
.A(n_10617),
.B(n_271),
.C(n_272),
.Y(n_11254)
);

INVx1_ASAP7_75t_SL g11255 ( 
.A(n_10453),
.Y(n_11255)
);

NOR3xp33_ASAP7_75t_L g11256 ( 
.A(n_10620),
.B(n_272),
.C(n_273),
.Y(n_11256)
);

AO32x1_ASAP7_75t_L g11257 ( 
.A1(n_10521),
.A2(n_276),
.A3(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_11257)
);

NAND2xp5_ASAP7_75t_SL g11258 ( 
.A(n_10844),
.B(n_4870),
.Y(n_11258)
);

AOI21xp5_ASAP7_75t_L g11259 ( 
.A1(n_10482),
.A2(n_4872),
.B(n_4871),
.Y(n_11259)
);

AOI21xp5_ASAP7_75t_L g11260 ( 
.A1(n_10532),
.A2(n_4874),
.B(n_4873),
.Y(n_11260)
);

OA22x2_ASAP7_75t_L g11261 ( 
.A1(n_10543),
.A2(n_277),
.B1(n_274),
.B2(n_275),
.Y(n_11261)
);

BUFx8_ASAP7_75t_L g11262 ( 
.A(n_10573),
.Y(n_11262)
);

BUFx6f_ASAP7_75t_L g11263 ( 
.A(n_10369),
.Y(n_11263)
);

AOI21xp5_ASAP7_75t_L g11264 ( 
.A1(n_10543),
.A2(n_4876),
.B(n_4875),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_10525),
.Y(n_11265)
);

AOI21xp5_ASAP7_75t_L g11266 ( 
.A1(n_10536),
.A2(n_4878),
.B(n_4877),
.Y(n_11266)
);

INVx2_ASAP7_75t_L g11267 ( 
.A(n_10541),
.Y(n_11267)
);

NOR2xp33_ASAP7_75t_L g11268 ( 
.A(n_10736),
.B(n_4879),
.Y(n_11268)
);

AND2x2_ASAP7_75t_SL g11269 ( 
.A(n_10693),
.B(n_278),
.Y(n_11269)
);

OAI21xp5_ASAP7_75t_L g11270 ( 
.A1(n_10640),
.A2(n_278),
.B(n_279),
.Y(n_11270)
);

AOI21x1_ASAP7_75t_L g11271 ( 
.A1(n_10351),
.A2(n_4881),
.B(n_4880),
.Y(n_11271)
);

AOI21xp5_ASAP7_75t_L g11272 ( 
.A1(n_10547),
.A2(n_4884),
.B(n_4882),
.Y(n_11272)
);

OAI21xp5_ASAP7_75t_L g11273 ( 
.A1(n_10647),
.A2(n_279),
.B(n_280),
.Y(n_11273)
);

OAI22xp5_ASAP7_75t_L g11274 ( 
.A1(n_10821),
.A2(n_283),
.B1(n_280),
.B2(n_282),
.Y(n_11274)
);

NAND3xp33_ASAP7_75t_L g11275 ( 
.A(n_10622),
.B(n_282),
.C(n_283),
.Y(n_11275)
);

NAND2xp5_ASAP7_75t_L g11276 ( 
.A(n_10414),
.B(n_284),
.Y(n_11276)
);

O2A1O1Ixp33_ASAP7_75t_L g11277 ( 
.A1(n_10902),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_11277)
);

HB1xp67_ASAP7_75t_L g11278 ( 
.A(n_10553),
.Y(n_11278)
);

INVxp67_ASAP7_75t_L g11279 ( 
.A(n_10514),
.Y(n_11279)
);

NOR3xp33_ASAP7_75t_L g11280 ( 
.A(n_10629),
.B(n_285),
.C(n_286),
.Y(n_11280)
);

OAI21xp5_ASAP7_75t_L g11281 ( 
.A1(n_10661),
.A2(n_287),
.B(n_288),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_L g11282 ( 
.A(n_10362),
.B(n_287),
.Y(n_11282)
);

AOI21xp5_ASAP7_75t_L g11283 ( 
.A1(n_10577),
.A2(n_4886),
.B(n_4885),
.Y(n_11283)
);

O2A1O1Ixp33_ASAP7_75t_L g11284 ( 
.A1(n_10905),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_11284)
);

O2A1O1Ixp33_ASAP7_75t_L g11285 ( 
.A1(n_10916),
.A2(n_293),
.B(n_290),
.C(n_292),
.Y(n_11285)
);

NAND2xp5_ASAP7_75t_L g11286 ( 
.A(n_10365),
.B(n_292),
.Y(n_11286)
);

AOI22xp33_ASAP7_75t_L g11287 ( 
.A1(n_10559),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_11287)
);

NOR2xp33_ASAP7_75t_SL g11288 ( 
.A(n_10882),
.B(n_4887),
.Y(n_11288)
);

AOI21xp5_ASAP7_75t_L g11289 ( 
.A1(n_10582),
.A2(n_4889),
.B(n_4888),
.Y(n_11289)
);

INVx2_ASAP7_75t_L g11290 ( 
.A(n_10585),
.Y(n_11290)
);

NAND2xp5_ASAP7_75t_SL g11291 ( 
.A(n_10790),
.B(n_4890),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_10598),
.Y(n_11292)
);

NOR2x1_ASAP7_75t_L g11293 ( 
.A(n_10709),
.B(n_295),
.Y(n_11293)
);

BUFx12f_ASAP7_75t_L g11294 ( 
.A(n_10519),
.Y(n_11294)
);

AOI21xp5_ASAP7_75t_L g11295 ( 
.A1(n_10618),
.A2(n_4892),
.B(n_4891),
.Y(n_11295)
);

AOI21xp5_ASAP7_75t_L g11296 ( 
.A1(n_10621),
.A2(n_4894),
.B(n_4893),
.Y(n_11296)
);

NAND3xp33_ASAP7_75t_L g11297 ( 
.A(n_10633),
.B(n_10683),
.C(n_10563),
.Y(n_11297)
);

OAI22xp5_ASAP7_75t_L g11298 ( 
.A1(n_10676),
.A2(n_10922),
.B1(n_10936),
.B2(n_10930),
.Y(n_11298)
);

NOR2xp33_ASAP7_75t_SL g11299 ( 
.A(n_10569),
.B(n_10440),
.Y(n_11299)
);

A2O1A1Ixp33_ASAP7_75t_L g11300 ( 
.A1(n_10675),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_11300)
);

A2O1A1Ixp33_ASAP7_75t_L g11301 ( 
.A1(n_10945),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_11301)
);

INVx2_ASAP7_75t_L g11302 ( 
.A(n_10419),
.Y(n_11302)
);

NAND2xp5_ASAP7_75t_L g11303 ( 
.A(n_10367),
.B(n_299),
.Y(n_11303)
);

OAI22x1_ASAP7_75t_L g11304 ( 
.A1(n_10497),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_11304)
);

NAND2xp5_ASAP7_75t_L g11305 ( 
.A(n_10416),
.B(n_300),
.Y(n_11305)
);

NOR2xp33_ASAP7_75t_L g11306 ( 
.A(n_10692),
.B(n_4896),
.Y(n_11306)
);

AOI21xp5_ASAP7_75t_L g11307 ( 
.A1(n_10608),
.A2(n_4899),
.B(n_4898),
.Y(n_11307)
);

AOI21xp5_ASAP7_75t_L g11308 ( 
.A1(n_10418),
.A2(n_10887),
.B(n_10860),
.Y(n_11308)
);

AOI22xp5_ASAP7_75t_L g11309 ( 
.A1(n_10517),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_11309)
);

O2A1O1Ixp33_ASAP7_75t_L g11310 ( 
.A1(n_10946),
.A2(n_10952),
.B(n_10961),
.C(n_10958),
.Y(n_11310)
);

NAND2xp5_ASAP7_75t_L g11311 ( 
.A(n_10904),
.B(n_303),
.Y(n_11311)
);

AOI21xp5_ASAP7_75t_L g11312 ( 
.A1(n_10910),
.A2(n_4901),
.B(n_4900),
.Y(n_11312)
);

AOI21xp5_ASAP7_75t_L g11313 ( 
.A1(n_10912),
.A2(n_10941),
.B(n_10918),
.Y(n_11313)
);

A2O1A1Ixp33_ASAP7_75t_L g11314 ( 
.A1(n_10508),
.A2(n_10515),
.B(n_10513),
.C(n_10737),
.Y(n_11314)
);

HB1xp67_ASAP7_75t_L g11315 ( 
.A(n_10496),
.Y(n_11315)
);

BUFx12f_ASAP7_75t_L g11316 ( 
.A(n_10359),
.Y(n_11316)
);

INVx2_ASAP7_75t_L g11317 ( 
.A(n_10420),
.Y(n_11317)
);

NAND2xp5_ASAP7_75t_SL g11318 ( 
.A(n_10790),
.B(n_4903),
.Y(n_11318)
);

A2O1A1Ixp33_ASAP7_75t_L g11319 ( 
.A1(n_10741),
.A2(n_306),
.B(n_304),
.C(n_305),
.Y(n_11319)
);

NAND2xp5_ASAP7_75t_L g11320 ( 
.A(n_10943),
.B(n_306),
.Y(n_11320)
);

NAND2xp5_ASAP7_75t_L g11321 ( 
.A(n_10944),
.B(n_307),
.Y(n_11321)
);

BUFx8_ASAP7_75t_L g11322 ( 
.A(n_10348),
.Y(n_11322)
);

CKINVDCx8_ASAP7_75t_R g11323 ( 
.A(n_10461),
.Y(n_11323)
);

OAI21xp5_ASAP7_75t_L g11324 ( 
.A1(n_10803),
.A2(n_307),
.B(n_308),
.Y(n_11324)
);

NAND2xp5_ASAP7_75t_SL g11325 ( 
.A(n_10754),
.B(n_4904),
.Y(n_11325)
);

AND2x4_ASAP7_75t_L g11326 ( 
.A(n_10587),
.B(n_4905),
.Y(n_11326)
);

NAND2xp5_ASAP7_75t_L g11327 ( 
.A(n_10947),
.B(n_308),
.Y(n_11327)
);

INVx1_ASAP7_75t_L g11328 ( 
.A(n_10948),
.Y(n_11328)
);

AOI21xp5_ASAP7_75t_L g11329 ( 
.A1(n_10953),
.A2(n_4908),
.B(n_4907),
.Y(n_11329)
);

AOI21xp5_ASAP7_75t_L g11330 ( 
.A1(n_10962),
.A2(n_4911),
.B(n_4910),
.Y(n_11330)
);

O2A1O1Ixp33_ASAP7_75t_L g11331 ( 
.A1(n_10435),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_11331)
);

NAND2xp5_ASAP7_75t_SL g11332 ( 
.A(n_10791),
.B(n_4915),
.Y(n_11332)
);

AOI21xp5_ASAP7_75t_L g11333 ( 
.A1(n_10662),
.A2(n_4917),
.B(n_4916),
.Y(n_11333)
);

NAND2xp5_ASAP7_75t_L g11334 ( 
.A(n_10427),
.B(n_310),
.Y(n_11334)
);

INVx2_ASAP7_75t_L g11335 ( 
.A(n_10446),
.Y(n_11335)
);

INVx1_ASAP7_75t_L g11336 ( 
.A(n_10450),
.Y(n_11336)
);

OR2x2_ASAP7_75t_L g11337 ( 
.A(n_10898),
.B(n_312),
.Y(n_11337)
);

AOI21xp5_ASAP7_75t_L g11338 ( 
.A1(n_10782),
.A2(n_4919),
.B(n_4918),
.Y(n_11338)
);

INVx4_ASAP7_75t_L g11339 ( 
.A(n_10935),
.Y(n_11339)
);

NAND2xp5_ASAP7_75t_L g11340 ( 
.A(n_10464),
.B(n_312),
.Y(n_11340)
);

AOI21x1_ASAP7_75t_L g11341 ( 
.A1(n_10807),
.A2(n_4921),
.B(n_4920),
.Y(n_11341)
);

AOI21xp5_ASAP7_75t_L g11342 ( 
.A1(n_10374),
.A2(n_4923),
.B(n_4922),
.Y(n_11342)
);

OAI21xp5_ASAP7_75t_L g11343 ( 
.A1(n_10731),
.A2(n_313),
.B(n_314),
.Y(n_11343)
);

NAND2xp5_ASAP7_75t_L g11344 ( 
.A(n_10467),
.B(n_313),
.Y(n_11344)
);

NAND3xp33_ASAP7_75t_L g11345 ( 
.A(n_10765),
.B(n_316),
.C(n_317),
.Y(n_11345)
);

AOI21xp5_ASAP7_75t_L g11346 ( 
.A1(n_10758),
.A2(n_4926),
.B(n_4925),
.Y(n_11346)
);

O2A1O1Ixp33_ASAP7_75t_L g11347 ( 
.A1(n_10426),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_11347)
);

NAND2xp5_ASAP7_75t_L g11348 ( 
.A(n_10473),
.B(n_319),
.Y(n_11348)
);

NAND2xp5_ASAP7_75t_SL g11349 ( 
.A(n_10791),
.B(n_4928),
.Y(n_11349)
);

AOI21xp5_ASAP7_75t_L g11350 ( 
.A1(n_10769),
.A2(n_4930),
.B(n_4929),
.Y(n_11350)
);

NOR3xp33_ASAP7_75t_L g11351 ( 
.A(n_10817),
.B(n_10845),
.C(n_10431),
.Y(n_11351)
);

NOR2xp33_ASAP7_75t_L g11352 ( 
.A(n_10637),
.B(n_4931),
.Y(n_11352)
);

OAI21xp5_ASAP7_75t_L g11353 ( 
.A1(n_10775),
.A2(n_319),
.B(n_320),
.Y(n_11353)
);

NAND2xp5_ASAP7_75t_L g11354 ( 
.A(n_10478),
.B(n_320),
.Y(n_11354)
);

OAI22xp33_ASAP7_75t_L g11355 ( 
.A1(n_10492),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_11355)
);

NAND2xp5_ASAP7_75t_L g11356 ( 
.A(n_10484),
.B(n_321),
.Y(n_11356)
);

OAI22xp5_ASAP7_75t_L g11357 ( 
.A1(n_10789),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_11357)
);

NAND2xp5_ASAP7_75t_L g11358 ( 
.A(n_10488),
.B(n_325),
.Y(n_11358)
);

OAI21xp5_ASAP7_75t_L g11359 ( 
.A1(n_10783),
.A2(n_325),
.B(n_326),
.Y(n_11359)
);

AOI21xp5_ASAP7_75t_L g11360 ( 
.A1(n_10787),
.A2(n_4934),
.B(n_4933),
.Y(n_11360)
);

AOI21xp5_ASAP7_75t_L g11361 ( 
.A1(n_10792),
.A2(n_4936),
.B(n_4935),
.Y(n_11361)
);

AOI21xp5_ASAP7_75t_L g11362 ( 
.A1(n_10471),
.A2(n_4939),
.B(n_4937),
.Y(n_11362)
);

NAND2xp5_ASAP7_75t_SL g11363 ( 
.A(n_10799),
.B(n_4940),
.Y(n_11363)
);

AOI21xp5_ASAP7_75t_L g11364 ( 
.A1(n_10839),
.A2(n_4944),
.B(n_4943),
.Y(n_11364)
);

NAND2xp5_ASAP7_75t_SL g11365 ( 
.A(n_10799),
.B(n_4945),
.Y(n_11365)
);

CKINVDCx5p33_ASAP7_75t_R g11366 ( 
.A(n_10487),
.Y(n_11366)
);

A2O1A1Ixp33_ASAP7_75t_L g11367 ( 
.A1(n_10753),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_11367)
);

NAND2xp5_ASAP7_75t_L g11368 ( 
.A(n_10720),
.B(n_327),
.Y(n_11368)
);

NOR2xp33_ASAP7_75t_L g11369 ( 
.A(n_10722),
.B(n_4949),
.Y(n_11369)
);

NOR2xp33_ASAP7_75t_L g11370 ( 
.A(n_10678),
.B(n_4950),
.Y(n_11370)
);

NOR3xp33_ASAP7_75t_L g11371 ( 
.A(n_10603),
.B(n_328),
.C(n_329),
.Y(n_11371)
);

NAND2xp5_ASAP7_75t_SL g11372 ( 
.A(n_10566),
.B(n_4952),
.Y(n_11372)
);

NAND2x1_ASAP7_75t_L g11373 ( 
.A(n_10407),
.B(n_4954),
.Y(n_11373)
);

NAND2xp5_ASAP7_75t_L g11374 ( 
.A(n_10406),
.B(n_330),
.Y(n_11374)
);

AOI21xp5_ASAP7_75t_L g11375 ( 
.A1(n_10826),
.A2(n_4956),
.B(n_4955),
.Y(n_11375)
);

BUFx8_ASAP7_75t_L g11376 ( 
.A(n_10866),
.Y(n_11376)
);

CKINVDCx10_ASAP7_75t_R g11377 ( 
.A(n_10751),
.Y(n_11377)
);

AOI21xp5_ASAP7_75t_L g11378 ( 
.A1(n_10794),
.A2(n_4959),
.B(n_4958),
.Y(n_11378)
);

AOI21xp5_ASAP7_75t_L g11379 ( 
.A1(n_10716),
.A2(n_4961),
.B(n_4960),
.Y(n_11379)
);

INVx1_ASAP7_75t_L g11380 ( 
.A(n_10415),
.Y(n_11380)
);

BUFx6f_ASAP7_75t_L g11381 ( 
.A(n_10375),
.Y(n_11381)
);

NOR3xp33_ASAP7_75t_L g11382 ( 
.A(n_10656),
.B(n_330),
.C(n_331),
.Y(n_11382)
);

AOI21xp5_ASAP7_75t_L g11383 ( 
.A1(n_10732),
.A2(n_4963),
.B(n_4962),
.Y(n_11383)
);

INVx1_ASAP7_75t_SL g11384 ( 
.A(n_10501),
.Y(n_11384)
);

AOI22xp5_ASAP7_75t_L g11385 ( 
.A1(n_10517),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_11385)
);

AOI21xp5_ASAP7_75t_L g11386 ( 
.A1(n_10877),
.A2(n_4965),
.B(n_4964),
.Y(n_11386)
);

NAND2xp5_ASAP7_75t_L g11387 ( 
.A(n_10408),
.B(n_332),
.Y(n_11387)
);

AO22x1_ASAP7_75t_L g11388 ( 
.A1(n_10796),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_11388)
);

A2O1A1Ixp33_ASAP7_75t_L g11389 ( 
.A1(n_10763),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_11389)
);

OAI21x1_ASAP7_75t_L g11390 ( 
.A1(n_10613),
.A2(n_4967),
.B(n_4966),
.Y(n_11390)
);

INVx2_ASAP7_75t_SL g11391 ( 
.A(n_10410),
.Y(n_11391)
);

NAND2xp5_ASAP7_75t_SL g11392 ( 
.A(n_10566),
.B(n_4969),
.Y(n_11392)
);

OAI21xp5_ASAP7_75t_L g11393 ( 
.A1(n_10684),
.A2(n_336),
.B(n_337),
.Y(n_11393)
);

AOI21x1_ASAP7_75t_L g11394 ( 
.A1(n_10849),
.A2(n_4972),
.B(n_4970),
.Y(n_11394)
);

O2A1O1Ixp33_ASAP7_75t_L g11395 ( 
.A1(n_10744),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_11395)
);

NAND2xp5_ASAP7_75t_SL g11396 ( 
.A(n_10695),
.B(n_4973),
.Y(n_11396)
);

NAND2xp5_ASAP7_75t_SL g11397 ( 
.A(n_10730),
.B(n_4974),
.Y(n_11397)
);

NAND2xp5_ASAP7_75t_L g11398 ( 
.A(n_10460),
.B(n_338),
.Y(n_11398)
);

NOR2xp33_ASAP7_75t_L g11399 ( 
.A(n_10825),
.B(n_4976),
.Y(n_11399)
);

INVx2_ASAP7_75t_L g11400 ( 
.A(n_10588),
.Y(n_11400)
);

NAND2xp5_ASAP7_75t_L g11401 ( 
.A(n_10954),
.B(n_339),
.Y(n_11401)
);

HB1xp67_ASAP7_75t_L g11402 ( 
.A(n_10635),
.Y(n_11402)
);

NOR2xp33_ASAP7_75t_L g11403 ( 
.A(n_10611),
.B(n_4978),
.Y(n_11403)
);

NAND2xp5_ASAP7_75t_L g11404 ( 
.A(n_10648),
.B(n_340),
.Y(n_11404)
);

AOI21x1_ASAP7_75t_L g11405 ( 
.A1(n_10814),
.A2(n_10848),
.B(n_10752),
.Y(n_11405)
);

AOI22xp5_ASAP7_75t_L g11406 ( 
.A1(n_10837),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_11406)
);

NOR3xp33_ASAP7_75t_L g11407 ( 
.A(n_10625),
.B(n_341),
.C(n_343),
.Y(n_11407)
);

AOI21xp5_ASAP7_75t_L g11408 ( 
.A1(n_10834),
.A2(n_4980),
.B(n_4979),
.Y(n_11408)
);

AOI21xp5_ASAP7_75t_L g11409 ( 
.A1(n_10664),
.A2(n_4983),
.B(n_4981),
.Y(n_11409)
);

AOI21xp5_ASAP7_75t_L g11410 ( 
.A1(n_10664),
.A2(n_4986),
.B(n_4984),
.Y(n_11410)
);

AOI22xp33_ASAP7_75t_L g11411 ( 
.A1(n_10774),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_11411)
);

OAI21xp5_ASAP7_75t_L g11412 ( 
.A1(n_10686),
.A2(n_344),
.B(n_345),
.Y(n_11412)
);

NAND2xp5_ASAP7_75t_L g11413 ( 
.A(n_10698),
.B(n_346),
.Y(n_11413)
);

AOI21xp5_ASAP7_75t_L g11414 ( 
.A1(n_10415),
.A2(n_4988),
.B(n_4987),
.Y(n_11414)
);

AOI21xp5_ASAP7_75t_L g11415 ( 
.A1(n_10415),
.A2(n_4990),
.B(n_4989),
.Y(n_11415)
);

AND2x6_ASAP7_75t_L g11416 ( 
.A(n_10524),
.B(n_4991),
.Y(n_11416)
);

NAND2xp5_ASAP7_75t_L g11417 ( 
.A(n_10510),
.B(n_346),
.Y(n_11417)
);

AOI21x1_ASAP7_75t_L g11418 ( 
.A1(n_10706),
.A2(n_4993),
.B(n_4992),
.Y(n_11418)
);

OR2x2_ASAP7_75t_L g11419 ( 
.A(n_10626),
.B(n_347),
.Y(n_11419)
);

NOR2xp67_ASAP7_75t_L g11420 ( 
.A(n_10539),
.B(n_4994),
.Y(n_11420)
);

AOI21x1_ASAP7_75t_L g11421 ( 
.A1(n_10560),
.A2(n_4996),
.B(n_4995),
.Y(n_11421)
);

AOI21xp5_ASAP7_75t_L g11422 ( 
.A1(n_10454),
.A2(n_4999),
.B(n_4998),
.Y(n_11422)
);

AND2x4_ASAP7_75t_L g11423 ( 
.A(n_10589),
.B(n_5000),
.Y(n_11423)
);

NAND3xp33_ASAP7_75t_L g11424 ( 
.A(n_10500),
.B(n_348),
.C(n_349),
.Y(n_11424)
);

INVx1_ASAP7_75t_L g11425 ( 
.A(n_10612),
.Y(n_11425)
);

AOI21xp5_ASAP7_75t_L g11426 ( 
.A1(n_10644),
.A2(n_5002),
.B(n_5001),
.Y(n_11426)
);

AND2x2_ASAP7_75t_L g11427 ( 
.A(n_10363),
.B(n_5004),
.Y(n_11427)
);

AND2x2_ASAP7_75t_L g11428 ( 
.A(n_10353),
.B(n_5005),
.Y(n_11428)
);

AOI21x1_ASAP7_75t_L g11429 ( 
.A1(n_10717),
.A2(n_5008),
.B(n_5007),
.Y(n_11429)
);

OAI21xp5_ASAP7_75t_L g11430 ( 
.A1(n_10490),
.A2(n_348),
.B(n_349),
.Y(n_11430)
);

AO22x1_ASAP7_75t_L g11431 ( 
.A1(n_10796),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_11431)
);

BUFx4f_ASAP7_75t_L g11432 ( 
.A(n_10524),
.Y(n_11432)
);

AOI21xp5_ASAP7_75t_L g11433 ( 
.A1(n_10383),
.A2(n_5010),
.B(n_5009),
.Y(n_11433)
);

AOI22xp33_ASAP7_75t_L g11434 ( 
.A1(n_10643),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_11434)
);

NAND2xp5_ASAP7_75t_L g11435 ( 
.A(n_10457),
.B(n_354),
.Y(n_11435)
);

INVx1_ASAP7_75t_L g11436 ( 
.A(n_10421),
.Y(n_11436)
);

AOI21xp5_ASAP7_75t_L g11437 ( 
.A1(n_10412),
.A2(n_5012),
.B(n_5011),
.Y(n_11437)
);

NAND3xp33_ASAP7_75t_L g11438 ( 
.A(n_10505),
.B(n_354),
.C(n_355),
.Y(n_11438)
);

OR2x6_ASAP7_75t_SL g11439 ( 
.A(n_10411),
.B(n_355),
.Y(n_11439)
);

HB1xp67_ASAP7_75t_L g11440 ( 
.A(n_10591),
.Y(n_11440)
);

OAI21xp5_ASAP7_75t_L g11441 ( 
.A1(n_10704),
.A2(n_10558),
.B(n_10760),
.Y(n_11441)
);

OAI21xp5_ASAP7_75t_L g11442 ( 
.A1(n_10444),
.A2(n_356),
.B(n_357),
.Y(n_11442)
);

INVx1_ASAP7_75t_L g11443 ( 
.A(n_10436),
.Y(n_11443)
);

AOI21xp5_ASAP7_75t_L g11444 ( 
.A1(n_10859),
.A2(n_5014),
.B(n_5013),
.Y(n_11444)
);

OR2x2_ASAP7_75t_SL g11445 ( 
.A(n_10820),
.B(n_10713),
.Y(n_11445)
);

O2A1O1Ixp33_ASAP7_75t_L g11446 ( 
.A1(n_10738),
.A2(n_10827),
.B(n_10781),
.C(n_10739),
.Y(n_11446)
);

BUFx6f_ASAP7_75t_L g11447 ( 
.A(n_10379),
.Y(n_11447)
);

A2O1A1Ixp33_ASAP7_75t_L g11448 ( 
.A1(n_10701),
.A2(n_359),
.B(n_356),
.C(n_357),
.Y(n_11448)
);

AOI22xp5_ASAP7_75t_L g11449 ( 
.A1(n_10750),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_11449)
);

A2O1A1Ixp33_ASAP7_75t_L g11450 ( 
.A1(n_10555),
.A2(n_10726),
.B(n_10734),
.C(n_10721),
.Y(n_11450)
);

AOI22xp33_ASAP7_75t_L g11451 ( 
.A1(n_10796),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_11451)
);

INVx1_ASAP7_75t_L g11452 ( 
.A(n_10443),
.Y(n_11452)
);

NAND2x1p5_ASAP7_75t_L g11453 ( 
.A(n_10388),
.B(n_5015),
.Y(n_11453)
);

AND2x4_ASAP7_75t_L g11454 ( 
.A(n_10645),
.B(n_10649),
.Y(n_11454)
);

BUFx12f_ASAP7_75t_L g11455 ( 
.A(n_10876),
.Y(n_11455)
);

INVx2_ASAP7_75t_L g11456 ( 
.A(n_10456),
.Y(n_11456)
);

AOI21xp5_ASAP7_75t_L g11457 ( 
.A1(n_10863),
.A2(n_5018),
.B(n_5017),
.Y(n_11457)
);

NAND2xp5_ASAP7_75t_L g11458 ( 
.A(n_10619),
.B(n_363),
.Y(n_11458)
);

OAI21xp5_ASAP7_75t_L g11459 ( 
.A1(n_10526),
.A2(n_363),
.B(n_364),
.Y(n_11459)
);

AOI21xp5_ASAP7_75t_L g11460 ( 
.A1(n_10871),
.A2(n_5020),
.B(n_5019),
.Y(n_11460)
);

O2A1O1Ixp33_ASAP7_75t_L g11461 ( 
.A1(n_10801),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_11461)
);

CKINVDCx5p33_ASAP7_75t_R g11462 ( 
.A(n_10509),
.Y(n_11462)
);

NAND2x1_ASAP7_75t_L g11463 ( 
.A(n_10884),
.B(n_5021),
.Y(n_11463)
);

AOI22xp33_ASAP7_75t_L g11464 ( 
.A1(n_10368),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_11464)
);

OAI22xp5_ASAP7_75t_L g11465 ( 
.A1(n_10506),
.A2(n_10820),
.B1(n_10584),
.B2(n_10653),
.Y(n_11465)
);

INVxp67_ASAP7_75t_SL g11466 ( 
.A(n_10480),
.Y(n_11466)
);

AOI22xp5_ASAP7_75t_L g11467 ( 
.A1(n_10371),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_11467)
);

AOI21x1_ASAP7_75t_L g11468 ( 
.A1(n_10540),
.A2(n_5023),
.B(n_5022),
.Y(n_11468)
);

NAND2xp5_ASAP7_75t_L g11469 ( 
.A(n_10463),
.B(n_369),
.Y(n_11469)
);

NOR2xp67_ASAP7_75t_L g11470 ( 
.A(n_10544),
.B(n_5024),
.Y(n_11470)
);

O2A1O1Ixp33_ASAP7_75t_L g11471 ( 
.A1(n_10843),
.A2(n_372),
.B(n_370),
.C(n_371),
.Y(n_11471)
);

NAND2xp5_ASAP7_75t_L g11472 ( 
.A(n_10466),
.B(n_370),
.Y(n_11472)
);

AOI22xp5_ASAP7_75t_L g11473 ( 
.A1(n_10373),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_11473)
);

AOI21xp5_ASAP7_75t_L g11474 ( 
.A1(n_10925),
.A2(n_5026),
.B(n_5025),
.Y(n_11474)
);

HB1xp67_ASAP7_75t_L g11475 ( 
.A(n_10529),
.Y(n_11475)
);

OAI21xp33_ASAP7_75t_SL g11476 ( 
.A1(n_10549),
.A2(n_373),
.B(n_374),
.Y(n_11476)
);

AND2x2_ASAP7_75t_L g11477 ( 
.A(n_10358),
.B(n_5027),
.Y(n_11477)
);

AND2x2_ASAP7_75t_L g11478 ( 
.A(n_10858),
.B(n_5028),
.Y(n_11478)
);

NAND2xp5_ASAP7_75t_L g11479 ( 
.A(n_10468),
.B(n_374),
.Y(n_11479)
);

OAI21xp5_ASAP7_75t_L g11480 ( 
.A1(n_10382),
.A2(n_375),
.B(n_376),
.Y(n_11480)
);

AOI22xp5_ASAP7_75t_L g11481 ( 
.A1(n_10594),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_11481)
);

INVxp67_ASAP7_75t_L g11482 ( 
.A(n_10486),
.Y(n_11482)
);

NAND2xp5_ASAP7_75t_L g11483 ( 
.A(n_10862),
.B(n_378),
.Y(n_11483)
);

AOI21xp5_ASAP7_75t_L g11484 ( 
.A1(n_10942),
.A2(n_5031),
.B(n_5030),
.Y(n_11484)
);

INVxp33_ASAP7_75t_SL g11485 ( 
.A(n_10743),
.Y(n_11485)
);

NAND2xp5_ASAP7_75t_L g11486 ( 
.A(n_10864),
.B(n_378),
.Y(n_11486)
);

AND2x2_ASAP7_75t_L g11487 ( 
.A(n_10865),
.B(n_10869),
.Y(n_11487)
);

AOI21xp5_ASAP7_75t_L g11488 ( 
.A1(n_10884),
.A2(n_5034),
.B(n_5033),
.Y(n_11488)
);

O2A1O1Ixp33_ASAP7_75t_L g11489 ( 
.A1(n_10764),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_11489)
);

NAND2xp5_ASAP7_75t_L g11490 ( 
.A(n_10872),
.B(n_379),
.Y(n_11490)
);

INVx1_ASAP7_75t_SL g11491 ( 
.A(n_10465),
.Y(n_11491)
);

AOI21xp5_ASAP7_75t_L g11492 ( 
.A1(n_10884),
.A2(n_5037),
.B(n_5036),
.Y(n_11492)
);

OR2x2_ASAP7_75t_L g11493 ( 
.A(n_10873),
.B(n_380),
.Y(n_11493)
);

AOI21xp5_ASAP7_75t_L g11494 ( 
.A1(n_10441),
.A2(n_5039),
.B(n_5038),
.Y(n_11494)
);

NOR3xp33_ASAP7_75t_L g11495 ( 
.A(n_10402),
.B(n_381),
.C(n_382),
.Y(n_11495)
);

NAND2xp5_ASAP7_75t_L g11496 ( 
.A(n_10875),
.B(n_382),
.Y(n_11496)
);

OAI21xp33_ASAP7_75t_L g11497 ( 
.A1(n_10391),
.A2(n_383),
.B(n_384),
.Y(n_11497)
);

INVx2_ASAP7_75t_L g11498 ( 
.A(n_10653),
.Y(n_11498)
);

AOI21xp5_ASAP7_75t_L g11499 ( 
.A1(n_10552),
.A2(n_5042),
.B(n_5041),
.Y(n_11499)
);

OAI321xp33_ASAP7_75t_L g11500 ( 
.A1(n_10387),
.A2(n_385),
.A3(n_387),
.B1(n_383),
.B2(n_384),
.C(n_386),
.Y(n_11500)
);

OAI21xp5_ASAP7_75t_L g11501 ( 
.A1(n_10878),
.A2(n_385),
.B(n_387),
.Y(n_11501)
);

NAND2xp5_ASAP7_75t_L g11502 ( 
.A(n_10881),
.B(n_388),
.Y(n_11502)
);

NAND2xp5_ASAP7_75t_L g11503 ( 
.A(n_10883),
.B(n_388),
.Y(n_11503)
);

NOR2xp33_ASAP7_75t_SL g11504 ( 
.A(n_10642),
.B(n_5043),
.Y(n_11504)
);

NAND2xp5_ASAP7_75t_SL g11505 ( 
.A(n_10713),
.B(n_10475),
.Y(n_11505)
);

A2O1A1Ixp33_ASAP7_75t_L g11506 ( 
.A1(n_10399),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_11506)
);

INVx1_ASAP7_75t_L g11507 ( 
.A(n_10596),
.Y(n_11507)
);

O2A1O1Ixp33_ASAP7_75t_L g11508 ( 
.A1(n_10886),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_11508)
);

INVx1_ASAP7_75t_L g11509 ( 
.A(n_10609),
.Y(n_11509)
);

NAND2xp5_ASAP7_75t_L g11510 ( 
.A(n_10888),
.B(n_392),
.Y(n_11510)
);

NAND2xp5_ASAP7_75t_L g11511 ( 
.A(n_10893),
.B(n_392),
.Y(n_11511)
);

OAI22xp5_ASAP7_75t_L g11512 ( 
.A1(n_10546),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_11512)
);

HB1xp67_ASAP7_75t_L g11513 ( 
.A(n_10481),
.Y(n_11513)
);

INVx2_ASAP7_75t_L g11514 ( 
.A(n_10610),
.Y(n_11514)
);

OR2x6_ASAP7_75t_L g11515 ( 
.A(n_10442),
.B(n_5044),
.Y(n_11515)
);

AOI21xp5_ASAP7_75t_L g11516 ( 
.A1(n_10489),
.A2(n_5046),
.B(n_5045),
.Y(n_11516)
);

INVx1_ASAP7_75t_SL g11517 ( 
.A(n_10504),
.Y(n_11517)
);

AOI21xp5_ASAP7_75t_L g11518 ( 
.A1(n_10458),
.A2(n_5048),
.B(n_5047),
.Y(n_11518)
);

AOI21x1_ASAP7_75t_L g11519 ( 
.A1(n_10567),
.A2(n_5050),
.B(n_5049),
.Y(n_11519)
);

AND2x2_ASAP7_75t_L g11520 ( 
.A(n_10896),
.B(n_5051),
.Y(n_11520)
);

OAI22xp33_ASAP7_75t_L g11521 ( 
.A1(n_10523),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_11521)
);

NAND2xp5_ASAP7_75t_L g11522 ( 
.A(n_10899),
.B(n_396),
.Y(n_11522)
);

AOI21xp5_ASAP7_75t_L g11523 ( 
.A1(n_10909),
.A2(n_5054),
.B(n_5052),
.Y(n_11523)
);

NAND2xp5_ASAP7_75t_L g11524 ( 
.A(n_10911),
.B(n_396),
.Y(n_11524)
);

O2A1O1Ixp33_ASAP7_75t_L g11525 ( 
.A1(n_10915),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_11525)
);

O2A1O1Ixp33_ASAP7_75t_L g11526 ( 
.A1(n_10919),
.A2(n_400),
.B(n_397),
.C(n_398),
.Y(n_11526)
);

INVx2_ASAP7_75t_L g11527 ( 
.A(n_10568),
.Y(n_11527)
);

AOI221xp5_ASAP7_75t_L g11528 ( 
.A1(n_10924),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.C(n_403),
.Y(n_11528)
);

BUFx6f_ASAP7_75t_L g11529 ( 
.A(n_10504),
.Y(n_11529)
);

AOI21xp5_ASAP7_75t_L g11530 ( 
.A1(n_10965),
.A2(n_5057),
.B(n_5055),
.Y(n_11530)
);

CKINVDCx16_ASAP7_75t_R g11531 ( 
.A(n_10927),
.Y(n_11531)
);

NAND2xp5_ASAP7_75t_L g11532 ( 
.A(n_10929),
.B(n_401),
.Y(n_11532)
);

AOI21xp5_ASAP7_75t_L g11533 ( 
.A1(n_10937),
.A2(n_5059),
.B(n_5058),
.Y(n_11533)
);

BUFx8_ASAP7_75t_L g11534 ( 
.A(n_10914),
.Y(n_11534)
);

AND2x2_ASAP7_75t_L g11535 ( 
.A(n_10938),
.B(n_5062),
.Y(n_11535)
);

AOI21x1_ASAP7_75t_L g11536 ( 
.A1(n_10579),
.A2(n_5065),
.B(n_5064),
.Y(n_11536)
);

OAI21x1_ASAP7_75t_L g11537 ( 
.A1(n_10385),
.A2(n_5067),
.B(n_5066),
.Y(n_11537)
);

NAND2xp5_ASAP7_75t_L g11538 ( 
.A(n_10939),
.B(n_402),
.Y(n_11538)
);

AOI22x1_ASAP7_75t_L g11539 ( 
.A1(n_10868),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_11539)
);

OAI21xp5_ASAP7_75t_L g11540 ( 
.A1(n_10964),
.A2(n_406),
.B(n_407),
.Y(n_11540)
);

AO21x1_ASAP7_75t_L g11541 ( 
.A1(n_10583),
.A2(n_10957),
.B(n_10956),
.Y(n_11541)
);

NAND2xp5_ASAP7_75t_L g11542 ( 
.A(n_10959),
.B(n_407),
.Y(n_11542)
);

OAI21xp5_ASAP7_75t_L g11543 ( 
.A1(n_10422),
.A2(n_408),
.B(n_409),
.Y(n_11543)
);

NAND2xp5_ASAP7_75t_L g11544 ( 
.A(n_10512),
.B(n_408),
.Y(n_11544)
);

NOR3xp33_ASAP7_75t_L g11545 ( 
.A(n_10879),
.B(n_409),
.C(n_410),
.Y(n_11545)
);

INVx2_ASAP7_75t_L g11546 ( 
.A(n_10557),
.Y(n_11546)
);

AOI22xp5_ASAP7_75t_L g11547 ( 
.A1(n_10894),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_11547)
);

AND2x4_ASAP7_75t_L g11548 ( 
.A(n_10395),
.B(n_5068),
.Y(n_11548)
);

INVx4_ASAP7_75t_L g11549 ( 
.A(n_10557),
.Y(n_11549)
);

OAI21xp33_ASAP7_75t_L g11550 ( 
.A1(n_10495),
.A2(n_411),
.B(n_412),
.Y(n_11550)
);

NOR2xp33_ASAP7_75t_L g11551 ( 
.A(n_10495),
.B(n_5069),
.Y(n_11551)
);

NAND2xp5_ASAP7_75t_L g11552 ( 
.A(n_10499),
.B(n_413),
.Y(n_11552)
);

AOI21xp5_ASAP7_75t_L g11553 ( 
.A1(n_10499),
.A2(n_5071),
.B(n_5070),
.Y(n_11553)
);

AOI21xp5_ASAP7_75t_L g11554 ( 
.A1(n_10590),
.A2(n_5074),
.B(n_5072),
.Y(n_11554)
);

AOI21xp5_ASAP7_75t_L g11555 ( 
.A1(n_10590),
.A2(n_5077),
.B(n_5075),
.Y(n_11555)
);

BUFx2_ASAP7_75t_L g11556 ( 
.A(n_10889),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_10641),
.Y(n_11557)
);

O2A1O1Ixp33_ASAP7_75t_SL g11558 ( 
.A1(n_10535),
.A2(n_415),
.B(n_413),
.C(n_414),
.Y(n_11558)
);

CKINVDCx16_ASAP7_75t_R g11559 ( 
.A(n_10438),
.Y(n_11559)
);

NAND2xp5_ASAP7_75t_L g11560 ( 
.A(n_10360),
.B(n_414),
.Y(n_11560)
);

OAI21xp5_ASAP7_75t_L g11561 ( 
.A1(n_10590),
.A2(n_415),
.B(n_416),
.Y(n_11561)
);

NOR2x1_ASAP7_75t_L g11562 ( 
.A(n_10818),
.B(n_416),
.Y(n_11562)
);

NOR2xp33_ASAP7_75t_SL g11563 ( 
.A(n_10691),
.B(n_5079),
.Y(n_11563)
);

HB1xp67_ASAP7_75t_L g11564 ( 
.A(n_10913),
.Y(n_11564)
);

AOI22xp33_ASAP7_75t_L g11565 ( 
.A1(n_10823),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_11565)
);

NAND2xp5_ASAP7_75t_L g11566 ( 
.A(n_10360),
.B(n_417),
.Y(n_11566)
);

NAND2xp5_ASAP7_75t_L g11567 ( 
.A(n_10360),
.B(n_418),
.Y(n_11567)
);

AND2x2_ASAP7_75t_L g11568 ( 
.A(n_10815),
.B(n_5080),
.Y(n_11568)
);

A2O1A1Ixp33_ASAP7_75t_L g11569 ( 
.A1(n_10535),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_SL g11570 ( 
.A(n_10516),
.B(n_5081),
.Y(n_11570)
);

INVx1_ASAP7_75t_L g11571 ( 
.A(n_10641),
.Y(n_11571)
);

BUFx6f_ASAP7_75t_L g11572 ( 
.A(n_10880),
.Y(n_11572)
);

AOI21x1_ASAP7_75t_L g11573 ( 
.A1(n_10703),
.A2(n_5083),
.B(n_5082),
.Y(n_11573)
);

NOR2xp33_ASAP7_75t_L g11574 ( 
.A(n_10592),
.B(n_5086),
.Y(n_11574)
);

NOR2xp33_ASAP7_75t_L g11575 ( 
.A(n_10592),
.B(n_5087),
.Y(n_11575)
);

NOR2xp33_ASAP7_75t_L g11576 ( 
.A(n_10592),
.B(n_5088),
.Y(n_11576)
);

AOI21xp5_ASAP7_75t_L g11577 ( 
.A1(n_10590),
.A2(n_5094),
.B(n_5093),
.Y(n_11577)
);

AOI21xp5_ASAP7_75t_L g11578 ( 
.A1(n_10590),
.A2(n_5096),
.B(n_5095),
.Y(n_11578)
);

NAND2xp5_ASAP7_75t_L g11579 ( 
.A(n_10360),
.B(n_421),
.Y(n_11579)
);

BUFx4f_ASAP7_75t_L g11580 ( 
.A(n_10393),
.Y(n_11580)
);

AOI21xp5_ASAP7_75t_L g11581 ( 
.A1(n_10590),
.A2(n_5099),
.B(n_5098),
.Y(n_11581)
);

AOI21xp5_ASAP7_75t_L g11582 ( 
.A1(n_10590),
.A2(n_5101),
.B(n_5100),
.Y(n_11582)
);

AND2x4_ASAP7_75t_L g11583 ( 
.A(n_10502),
.B(n_5102),
.Y(n_11583)
);

AOI21xp5_ASAP7_75t_L g11584 ( 
.A1(n_10590),
.A2(n_5104),
.B(n_5103),
.Y(n_11584)
);

AND2x4_ASAP7_75t_L g11585 ( 
.A(n_10502),
.B(n_5105),
.Y(n_11585)
);

AOI22xp33_ASAP7_75t_SL g11586 ( 
.A1(n_10381),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_11586)
);

AOI21xp5_ASAP7_75t_L g11587 ( 
.A1(n_10590),
.A2(n_5107),
.B(n_5106),
.Y(n_11587)
);

INVx1_ASAP7_75t_L g11588 ( 
.A(n_10641),
.Y(n_11588)
);

AOI21xp5_ASAP7_75t_L g11589 ( 
.A1(n_10590),
.A2(n_5109),
.B(n_5108),
.Y(n_11589)
);

CKINVDCx5p33_ASAP7_75t_R g11590 ( 
.A(n_10479),
.Y(n_11590)
);

NAND2xp5_ASAP7_75t_L g11591 ( 
.A(n_10360),
.B(n_423),
.Y(n_11591)
);

INVx1_ASAP7_75t_L g11592 ( 
.A(n_10641),
.Y(n_11592)
);

NAND2xp5_ASAP7_75t_L g11593 ( 
.A(n_10360),
.B(n_425),
.Y(n_11593)
);

INVxp67_ASAP7_75t_SL g11594 ( 
.A(n_10641),
.Y(n_11594)
);

AOI21xp5_ASAP7_75t_L g11595 ( 
.A1(n_10590),
.A2(n_5111),
.B(n_5110),
.Y(n_11595)
);

BUFx12f_ASAP7_75t_L g11596 ( 
.A(n_10518),
.Y(n_11596)
);

NAND2xp5_ASAP7_75t_L g11597 ( 
.A(n_10360),
.B(n_425),
.Y(n_11597)
);

NAND2xp5_ASAP7_75t_L g11598 ( 
.A(n_10360),
.B(n_426),
.Y(n_11598)
);

NOR2xp67_ASAP7_75t_L g11599 ( 
.A(n_10593),
.B(n_5112),
.Y(n_11599)
);

INVx1_ASAP7_75t_L g11600 ( 
.A(n_10641),
.Y(n_11600)
);

AOI21xp5_ASAP7_75t_L g11601 ( 
.A1(n_10590),
.A2(n_5114),
.B(n_5113),
.Y(n_11601)
);

NAND2xp5_ASAP7_75t_L g11602 ( 
.A(n_10360),
.B(n_427),
.Y(n_11602)
);

INVx2_ASAP7_75t_L g11603 ( 
.A(n_10345),
.Y(n_11603)
);

NAND2xp5_ASAP7_75t_L g11604 ( 
.A(n_10360),
.B(n_427),
.Y(n_11604)
);

NOR2xp33_ASAP7_75t_SL g11605 ( 
.A(n_10691),
.B(n_5115),
.Y(n_11605)
);

OAI21x1_ASAP7_75t_L g11606 ( 
.A1(n_10908),
.A2(n_5117),
.B(n_5116),
.Y(n_11606)
);

NAND2xp5_ASAP7_75t_L g11607 ( 
.A(n_10360),
.B(n_428),
.Y(n_11607)
);

AOI21xp5_ASAP7_75t_L g11608 ( 
.A1(n_10590),
.A2(n_5119),
.B(n_5118),
.Y(n_11608)
);

AOI21xp33_ASAP7_75t_L g11609 ( 
.A1(n_10590),
.A2(n_428),
.B(n_429),
.Y(n_11609)
);

INVx3_ASAP7_75t_L g11610 ( 
.A(n_10502),
.Y(n_11610)
);

NAND2xp5_ASAP7_75t_SL g11611 ( 
.A(n_10516),
.B(n_5120),
.Y(n_11611)
);

NAND2xp5_ASAP7_75t_L g11612 ( 
.A(n_10360),
.B(n_429),
.Y(n_11612)
);

AND2x2_ASAP7_75t_L g11613 ( 
.A(n_10815),
.B(n_5122),
.Y(n_11613)
);

OAI22xp5_ASAP7_75t_L g11614 ( 
.A1(n_10724),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_11614)
);

INVx3_ASAP7_75t_L g11615 ( 
.A(n_10502),
.Y(n_11615)
);

O2A1O1Ixp33_ASAP7_75t_SL g11616 ( 
.A1(n_10535),
.A2(n_433),
.B(n_430),
.C(n_431),
.Y(n_11616)
);

AOI21xp5_ASAP7_75t_L g11617 ( 
.A1(n_10590),
.A2(n_5124),
.B(n_5123),
.Y(n_11617)
);

NAND2xp5_ASAP7_75t_SL g11618 ( 
.A(n_10516),
.B(n_5125),
.Y(n_11618)
);

NAND2xp33_ASAP7_75t_L g11619 ( 
.A(n_10511),
.B(n_433),
.Y(n_11619)
);

INVx2_ASAP7_75t_L g11620 ( 
.A(n_10345),
.Y(n_11620)
);

AOI21xp5_ASAP7_75t_L g11621 ( 
.A1(n_10590),
.A2(n_5128),
.B(n_5126),
.Y(n_11621)
);

OAI21xp5_ASAP7_75t_L g11622 ( 
.A1(n_10590),
.A2(n_434),
.B(n_435),
.Y(n_11622)
);

NAND2xp5_ASAP7_75t_L g11623 ( 
.A(n_10360),
.B(n_434),
.Y(n_11623)
);

INVx1_ASAP7_75t_L g11624 ( 
.A(n_10641),
.Y(n_11624)
);

AOI21x1_ASAP7_75t_L g11625 ( 
.A1(n_10703),
.A2(n_5130),
.B(n_5129),
.Y(n_11625)
);

INVx2_ASAP7_75t_L g11626 ( 
.A(n_10345),
.Y(n_11626)
);

NAND2xp5_ASAP7_75t_L g11627 ( 
.A(n_10360),
.B(n_435),
.Y(n_11627)
);

INVx3_ASAP7_75t_L g11628 ( 
.A(n_10502),
.Y(n_11628)
);

AO21x1_ASAP7_75t_L g11629 ( 
.A1(n_10535),
.A2(n_436),
.B(n_437),
.Y(n_11629)
);

OAI21xp5_ASAP7_75t_L g11630 ( 
.A1(n_10590),
.A2(n_436),
.B(n_437),
.Y(n_11630)
);

NAND2xp5_ASAP7_75t_L g11631 ( 
.A(n_10360),
.B(n_438),
.Y(n_11631)
);

INVx3_ASAP7_75t_L g11632 ( 
.A(n_10502),
.Y(n_11632)
);

AOI21xp5_ASAP7_75t_L g11633 ( 
.A1(n_10590),
.A2(n_5132),
.B(n_5131),
.Y(n_11633)
);

AOI21x1_ASAP7_75t_L g11634 ( 
.A1(n_10703),
.A2(n_5134),
.B(n_5133),
.Y(n_11634)
);

AOI21xp5_ASAP7_75t_L g11635 ( 
.A1(n_10590),
.A2(n_5136),
.B(n_5135),
.Y(n_11635)
);

NAND2xp5_ASAP7_75t_L g11636 ( 
.A(n_10360),
.B(n_438),
.Y(n_11636)
);

A2O1A1Ixp33_ASAP7_75t_L g11637 ( 
.A1(n_10535),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_11637)
);

OAI22xp5_ASAP7_75t_L g11638 ( 
.A1(n_10724),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_11638)
);

INVx1_ASAP7_75t_L g11639 ( 
.A(n_10641),
.Y(n_11639)
);

AOI21xp5_ASAP7_75t_L g11640 ( 
.A1(n_10590),
.A2(n_5139),
.B(n_5138),
.Y(n_11640)
);

INVx2_ASAP7_75t_L g11641 ( 
.A(n_10345),
.Y(n_11641)
);

NAND2xp5_ASAP7_75t_L g11642 ( 
.A(n_10360),
.B(n_442),
.Y(n_11642)
);

INVxp67_ASAP7_75t_L g11643 ( 
.A(n_10913),
.Y(n_11643)
);

O2A1O1Ixp33_ASAP7_75t_L g11644 ( 
.A1(n_10535),
.A2(n_445),
.B(n_443),
.C(n_444),
.Y(n_11644)
);

NAND2xp5_ASAP7_75t_L g11645 ( 
.A(n_10360),
.B(n_443),
.Y(n_11645)
);

AND2x4_ASAP7_75t_SL g11646 ( 
.A(n_10344),
.B(n_5140),
.Y(n_11646)
);

NOR2xp33_ASAP7_75t_L g11647 ( 
.A(n_10592),
.B(n_5142),
.Y(n_11647)
);

AOI21xp5_ASAP7_75t_L g11648 ( 
.A1(n_10590),
.A2(n_5144),
.B(n_5143),
.Y(n_11648)
);

AOI21xp5_ASAP7_75t_L g11649 ( 
.A1(n_10590),
.A2(n_5146),
.B(n_5145),
.Y(n_11649)
);

NAND2xp5_ASAP7_75t_L g11650 ( 
.A(n_10360),
.B(n_444),
.Y(n_11650)
);

OR2x6_ASAP7_75t_L g11651 ( 
.A(n_10574),
.B(n_5147),
.Y(n_11651)
);

INVxp67_ASAP7_75t_L g11652 ( 
.A(n_10913),
.Y(n_11652)
);

NAND2xp5_ASAP7_75t_L g11653 ( 
.A(n_10360),
.B(n_446),
.Y(n_11653)
);

NAND2xp5_ASAP7_75t_L g11654 ( 
.A(n_10360),
.B(n_446),
.Y(n_11654)
);

INVx3_ASAP7_75t_L g11655 ( 
.A(n_10502),
.Y(n_11655)
);

INVx1_ASAP7_75t_L g11656 ( 
.A(n_10641),
.Y(n_11656)
);

AOI22xp5_ASAP7_75t_L g11657 ( 
.A1(n_10823),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_11657)
);

AOI21xp5_ASAP7_75t_L g11658 ( 
.A1(n_10590),
.A2(n_5150),
.B(n_5148),
.Y(n_11658)
);

OAI22xp5_ASAP7_75t_L g11659 ( 
.A1(n_10724),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_11659)
);

AOI21xp5_ASAP7_75t_L g11660 ( 
.A1(n_10590),
.A2(n_5153),
.B(n_5151),
.Y(n_11660)
);

BUFx6f_ASAP7_75t_L g11661 ( 
.A(n_10880),
.Y(n_11661)
);

A2O1A1Ixp33_ASAP7_75t_L g11662 ( 
.A1(n_10535),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_11662)
);

NAND2xp5_ASAP7_75t_L g11663 ( 
.A(n_10360),
.B(n_450),
.Y(n_11663)
);

AOI21xp5_ASAP7_75t_L g11664 ( 
.A1(n_10590),
.A2(n_5156),
.B(n_5155),
.Y(n_11664)
);

AOI21xp5_ASAP7_75t_L g11665 ( 
.A1(n_10590),
.A2(n_5161),
.B(n_5157),
.Y(n_11665)
);

NAND2xp5_ASAP7_75t_L g11666 ( 
.A(n_10360),
.B(n_452),
.Y(n_11666)
);

AOI21xp5_ASAP7_75t_L g11667 ( 
.A1(n_10590),
.A2(n_5164),
.B(n_5163),
.Y(n_11667)
);

INVx2_ASAP7_75t_SL g11668 ( 
.A(n_10880),
.Y(n_11668)
);

AOI21xp5_ASAP7_75t_L g11669 ( 
.A1(n_10590),
.A2(n_5167),
.B(n_5166),
.Y(n_11669)
);

NAND2xp5_ASAP7_75t_L g11670 ( 
.A(n_10360),
.B(n_453),
.Y(n_11670)
);

OAI22xp5_ASAP7_75t_L g11671 ( 
.A1(n_10724),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_11671)
);

INVx2_ASAP7_75t_L g11672 ( 
.A(n_10345),
.Y(n_11672)
);

NAND2xp5_ASAP7_75t_L g11673 ( 
.A(n_10360),
.B(n_454),
.Y(n_11673)
);

O2A1O1Ixp5_ASAP7_75t_L g11674 ( 
.A1(n_10535),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_11674)
);

INVx1_ASAP7_75t_L g11675 ( 
.A(n_10641),
.Y(n_11675)
);

NAND2xp5_ASAP7_75t_L g11676 ( 
.A(n_10360),
.B(n_457),
.Y(n_11676)
);

AOI21xp5_ASAP7_75t_L g11677 ( 
.A1(n_10590),
.A2(n_458),
.B(n_459),
.Y(n_11677)
);

AOI21xp5_ASAP7_75t_L g11678 ( 
.A1(n_10590),
.A2(n_458),
.B(n_459),
.Y(n_11678)
);

INVx1_ASAP7_75t_SL g11679 ( 
.A(n_10376),
.Y(n_11679)
);

A2O1A1Ixp33_ASAP7_75t_L g11680 ( 
.A1(n_10535),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_11680)
);

AOI21xp5_ASAP7_75t_L g11681 ( 
.A1(n_10590),
.A2(n_460),
.B(n_461),
.Y(n_11681)
);

AOI21xp5_ASAP7_75t_L g11682 ( 
.A1(n_10590),
.A2(n_463),
.B(n_464),
.Y(n_11682)
);

OAI22xp5_ASAP7_75t_L g11683 ( 
.A1(n_10724),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_11683)
);

A2O1A1Ixp33_ASAP7_75t_L g11684 ( 
.A1(n_10535),
.A2(n_468),
.B(n_465),
.C(n_466),
.Y(n_11684)
);

INVx2_ASAP7_75t_L g11685 ( 
.A(n_10345),
.Y(n_11685)
);

AOI21xp5_ASAP7_75t_L g11686 ( 
.A1(n_10590),
.A2(n_468),
.B(n_469),
.Y(n_11686)
);

AOI22xp33_ASAP7_75t_L g11687 ( 
.A1(n_10823),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_11687)
);

OAI22xp5_ASAP7_75t_L g11688 ( 
.A1(n_10724),
.A2(n_474),
.B1(n_471),
.B2(n_473),
.Y(n_11688)
);

OAI22xp5_ASAP7_75t_L g11689 ( 
.A1(n_10724),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_11689)
);

A2O1A1Ixp33_ASAP7_75t_L g11690 ( 
.A1(n_10535),
.A2(n_477),
.B(n_475),
.C(n_476),
.Y(n_11690)
);

OAI22xp5_ASAP7_75t_L g11691 ( 
.A1(n_10724),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_11691)
);

NAND2xp5_ASAP7_75t_L g11692 ( 
.A(n_10360),
.B(n_478),
.Y(n_11692)
);

NAND2xp5_ASAP7_75t_L g11693 ( 
.A(n_10360),
.B(n_479),
.Y(n_11693)
);

INVx1_ASAP7_75t_L g11694 ( 
.A(n_10641),
.Y(n_11694)
);

INVx2_ASAP7_75t_L g11695 ( 
.A(n_10345),
.Y(n_11695)
);

AOI21xp5_ASAP7_75t_L g11696 ( 
.A1(n_10590),
.A2(n_480),
.B(n_481),
.Y(n_11696)
);

NAND2xp5_ASAP7_75t_L g11697 ( 
.A(n_10360),
.B(n_481),
.Y(n_11697)
);

NAND2xp5_ASAP7_75t_L g11698 ( 
.A(n_10360),
.B(n_482),
.Y(n_11698)
);

BUFx3_ASAP7_75t_L g11699 ( 
.A(n_10880),
.Y(n_11699)
);

NAND2xp5_ASAP7_75t_L g11700 ( 
.A(n_10360),
.B(n_482),
.Y(n_11700)
);

NAND2xp5_ASAP7_75t_L g11701 ( 
.A(n_10360),
.B(n_483),
.Y(n_11701)
);

OA21x2_ASAP7_75t_L g11702 ( 
.A1(n_10829),
.A2(n_483),
.B(n_485),
.Y(n_11702)
);

INVx1_ASAP7_75t_L g11703 ( 
.A(n_10641),
.Y(n_11703)
);

AND2x2_ASAP7_75t_L g11704 ( 
.A(n_10815),
.B(n_486),
.Y(n_11704)
);

AOI22xp5_ASAP7_75t_L g11705 ( 
.A1(n_10823),
.A2(n_488),
.B1(n_486),
.B2(n_487),
.Y(n_11705)
);

OAI21x1_ASAP7_75t_L g11706 ( 
.A1(n_10908),
.A2(n_488),
.B(n_489),
.Y(n_11706)
);

BUFx4f_ASAP7_75t_L g11707 ( 
.A(n_10393),
.Y(n_11707)
);

AND2x2_ASAP7_75t_L g11708 ( 
.A(n_10815),
.B(n_489),
.Y(n_11708)
);

BUFx3_ASAP7_75t_L g11709 ( 
.A(n_10880),
.Y(n_11709)
);

NAND3xp33_ASAP7_75t_L g11710 ( 
.A(n_10472),
.B(n_490),
.C(n_491),
.Y(n_11710)
);

AOI22xp5_ASAP7_75t_L g11711 ( 
.A1(n_10823),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_11711)
);

INVx2_ASAP7_75t_L g11712 ( 
.A(n_10345),
.Y(n_11712)
);

BUFx6f_ASAP7_75t_L g11713 ( 
.A(n_10880),
.Y(n_11713)
);

AOI21xp5_ASAP7_75t_L g11714 ( 
.A1(n_10590),
.A2(n_492),
.B(n_493),
.Y(n_11714)
);

AOI22xp5_ASAP7_75t_L g11715 ( 
.A1(n_10823),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_11715)
);

AOI21xp5_ASAP7_75t_L g11716 ( 
.A1(n_10590),
.A2(n_495),
.B(n_496),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_10360),
.B(n_496),
.Y(n_11717)
);

AOI21xp5_ASAP7_75t_L g11718 ( 
.A1(n_10590),
.A2(n_497),
.B(n_498),
.Y(n_11718)
);

BUFx2_ASAP7_75t_L g11719 ( 
.A(n_10889),
.Y(n_11719)
);

NOR2xp33_ASAP7_75t_L g11720 ( 
.A(n_10592),
.B(n_497),
.Y(n_11720)
);

INVx1_ASAP7_75t_L g11721 ( 
.A(n_10641),
.Y(n_11721)
);

NAND2xp5_ASAP7_75t_L g11722 ( 
.A(n_10360),
.B(n_499),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_10641),
.Y(n_11723)
);

NOR2xp67_ASAP7_75t_L g11724 ( 
.A(n_10593),
.B(n_499),
.Y(n_11724)
);

INVx2_ASAP7_75t_L g11725 ( 
.A(n_10345),
.Y(n_11725)
);

CKINVDCx10_ASAP7_75t_R g11726 ( 
.A(n_10574),
.Y(n_11726)
);

AOI21xp5_ASAP7_75t_L g11727 ( 
.A1(n_10590),
.A2(n_500),
.B(n_501),
.Y(n_11727)
);

OAI22xp5_ASAP7_75t_L g11728 ( 
.A1(n_10724),
.A2(n_503),
.B1(n_500),
.B2(n_502),
.Y(n_11728)
);

NAND2xp5_ASAP7_75t_L g11729 ( 
.A(n_10360),
.B(n_502),
.Y(n_11729)
);

AO21x1_ASAP7_75t_L g11730 ( 
.A1(n_10535),
.A2(n_503),
.B(n_504),
.Y(n_11730)
);

NAND2xp5_ASAP7_75t_L g11731 ( 
.A(n_10360),
.B(n_504),
.Y(n_11731)
);

AOI21xp5_ASAP7_75t_L g11732 ( 
.A1(n_10590),
.A2(n_505),
.B(n_506),
.Y(n_11732)
);

AOI21xp5_ASAP7_75t_L g11733 ( 
.A1(n_10590),
.A2(n_505),
.B(n_506),
.Y(n_11733)
);

OAI21x1_ASAP7_75t_L g11734 ( 
.A1(n_10908),
.A2(n_507),
.B(n_508),
.Y(n_11734)
);

AOI21xp5_ASAP7_75t_L g11735 ( 
.A1(n_10590),
.A2(n_507),
.B(n_508),
.Y(n_11735)
);

BUFx3_ASAP7_75t_L g11736 ( 
.A(n_10880),
.Y(n_11736)
);

OAI21xp5_ASAP7_75t_L g11737 ( 
.A1(n_10590),
.A2(n_509),
.B(n_510),
.Y(n_11737)
);

AOI22xp5_ASAP7_75t_L g11738 ( 
.A1(n_10823),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_11738)
);

NAND2xp5_ASAP7_75t_L g11739 ( 
.A(n_10360),
.B(n_511),
.Y(n_11739)
);

INVx1_ASAP7_75t_L g11740 ( 
.A(n_10641),
.Y(n_11740)
);

NOR2xp33_ASAP7_75t_R g11741 ( 
.A(n_10438),
.B(n_512),
.Y(n_11741)
);

BUFx6f_ASAP7_75t_L g11742 ( 
.A(n_10880),
.Y(n_11742)
);

AOI21xp5_ASAP7_75t_L g11743 ( 
.A1(n_10590),
.A2(n_512),
.B(n_513),
.Y(n_11743)
);

CKINVDCx10_ASAP7_75t_R g11744 ( 
.A(n_10574),
.Y(n_11744)
);

CKINVDCx5p33_ASAP7_75t_R g11745 ( 
.A(n_10479),
.Y(n_11745)
);

AOI21xp5_ASAP7_75t_L g11746 ( 
.A1(n_10590),
.A2(n_513),
.B(n_514),
.Y(n_11746)
);

INVx3_ASAP7_75t_L g11747 ( 
.A(n_10502),
.Y(n_11747)
);

NAND3xp33_ASAP7_75t_L g11748 ( 
.A(n_10472),
.B(n_515),
.C(n_516),
.Y(n_11748)
);

NOR2xp67_ASAP7_75t_L g11749 ( 
.A(n_10593),
.B(n_515),
.Y(n_11749)
);

NAND2xp5_ASAP7_75t_SL g11750 ( 
.A(n_10516),
.B(n_517),
.Y(n_11750)
);

AOI21xp5_ASAP7_75t_L g11751 ( 
.A1(n_10590),
.A2(n_518),
.B(n_519),
.Y(n_11751)
);

A2O1A1Ixp33_ASAP7_75t_L g11752 ( 
.A1(n_10986),
.A2(n_11619),
.B(n_11148),
.C(n_11005),
.Y(n_11752)
);

NOR2xp33_ASAP7_75t_L g11753 ( 
.A(n_10971),
.B(n_518),
.Y(n_11753)
);

O2A1O1Ixp33_ASAP7_75t_L g11754 ( 
.A1(n_11136),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_11754)
);

OAI22xp33_ASAP7_75t_L g11755 ( 
.A1(n_11309),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_11755)
);

AND2x2_ASAP7_75t_L g11756 ( 
.A(n_11487),
.B(n_523),
.Y(n_11756)
);

INVx2_ASAP7_75t_L g11757 ( 
.A(n_11267),
.Y(n_11757)
);

NAND2xp5_ASAP7_75t_L g11758 ( 
.A(n_11091),
.B(n_523),
.Y(n_11758)
);

NOR2xp33_ASAP7_75t_L g11759 ( 
.A(n_11053),
.B(n_524),
.Y(n_11759)
);

AOI22xp5_ASAP7_75t_L g11760 ( 
.A1(n_11000),
.A2(n_11128),
.B1(n_11046),
.B2(n_10991),
.Y(n_11760)
);

BUFx3_ASAP7_75t_L g11761 ( 
.A(n_11316),
.Y(n_11761)
);

NOR2x1_ASAP7_75t_R g11762 ( 
.A(n_11218),
.B(n_525),
.Y(n_11762)
);

OR2x6_ASAP7_75t_L g11763 ( 
.A(n_10968),
.B(n_525),
.Y(n_11763)
);

INVx3_ASAP7_75t_L g11764 ( 
.A(n_11323),
.Y(n_11764)
);

NOR2xp33_ASAP7_75t_R g11765 ( 
.A(n_11590),
.B(n_526),
.Y(n_11765)
);

INVx2_ASAP7_75t_L g11766 ( 
.A(n_11290),
.Y(n_11766)
);

NAND2xp5_ASAP7_75t_L g11767 ( 
.A(n_11032),
.B(n_526),
.Y(n_11767)
);

AOI21xp5_ASAP7_75t_L g11768 ( 
.A1(n_10978),
.A2(n_527),
.B(n_528),
.Y(n_11768)
);

NAND2xp5_ASAP7_75t_L g11769 ( 
.A(n_11037),
.B(n_527),
.Y(n_11769)
);

INVx2_ASAP7_75t_L g11770 ( 
.A(n_11252),
.Y(n_11770)
);

INVx2_ASAP7_75t_L g11771 ( 
.A(n_11265),
.Y(n_11771)
);

NAND2xp5_ASAP7_75t_L g11772 ( 
.A(n_11564),
.B(n_528),
.Y(n_11772)
);

NAND2xp5_ASAP7_75t_L g11773 ( 
.A(n_11278),
.B(n_529),
.Y(n_11773)
);

AOI21xp5_ASAP7_75t_L g11774 ( 
.A1(n_10977),
.A2(n_529),
.B(n_530),
.Y(n_11774)
);

NAND2xp5_ASAP7_75t_L g11775 ( 
.A(n_11180),
.B(n_530),
.Y(n_11775)
);

NOR2xp33_ASAP7_75t_L g11776 ( 
.A(n_11610),
.B(n_531),
.Y(n_11776)
);

BUFx2_ASAP7_75t_L g11777 ( 
.A(n_11178),
.Y(n_11777)
);

NOR2xp33_ASAP7_75t_R g11778 ( 
.A(n_11745),
.B(n_531),
.Y(n_11778)
);

INVx2_ASAP7_75t_L g11779 ( 
.A(n_11292),
.Y(n_11779)
);

NAND2xp5_ASAP7_75t_L g11780 ( 
.A(n_11202),
.B(n_532),
.Y(n_11780)
);

OAI21x1_ASAP7_75t_SL g11781 ( 
.A1(n_11629),
.A2(n_532),
.B(n_533),
.Y(n_11781)
);

AOI21xp5_ASAP7_75t_L g11782 ( 
.A1(n_10994),
.A2(n_533),
.B(n_534),
.Y(n_11782)
);

HB1xp67_ASAP7_75t_L g11783 ( 
.A(n_11206),
.Y(n_11783)
);

A2O1A1Ixp33_ASAP7_75t_L g11784 ( 
.A1(n_10973),
.A2(n_11644),
.B(n_10979),
.C(n_11622),
.Y(n_11784)
);

AO21x1_ASAP7_75t_L g11785 ( 
.A1(n_11677),
.A2(n_534),
.B(n_535),
.Y(n_11785)
);

INVx4_ASAP7_75t_L g11786 ( 
.A(n_11012),
.Y(n_11786)
);

BUFx6f_ASAP7_75t_L g11787 ( 
.A(n_11012),
.Y(n_11787)
);

NAND2xp5_ASAP7_75t_L g11788 ( 
.A(n_11139),
.B(n_535),
.Y(n_11788)
);

AND2x2_ASAP7_75t_L g11789 ( 
.A(n_11456),
.B(n_536),
.Y(n_11789)
);

BUFx2_ASAP7_75t_L g11790 ( 
.A(n_11315),
.Y(n_11790)
);

NOR2xp33_ASAP7_75t_L g11791 ( 
.A(n_11615),
.B(n_537),
.Y(n_11791)
);

AOI21xp5_ASAP7_75t_L g11792 ( 
.A1(n_10995),
.A2(n_538),
.B(n_539),
.Y(n_11792)
);

AND2x4_ASAP7_75t_L g11793 ( 
.A(n_11556),
.B(n_538),
.Y(n_11793)
);

O2A1O1Ixp5_ASAP7_75t_L g11794 ( 
.A1(n_11730),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_11794)
);

A2O1A1Ixp33_ASAP7_75t_L g11795 ( 
.A1(n_11561),
.A2(n_543),
.B(n_541),
.C(n_542),
.Y(n_11795)
);

BUFx2_ASAP7_75t_L g11796 ( 
.A(n_11719),
.Y(n_11796)
);

NOR2xp33_ASAP7_75t_L g11797 ( 
.A(n_11628),
.B(n_543),
.Y(n_11797)
);

BUFx3_ASAP7_75t_L g11798 ( 
.A(n_11201),
.Y(n_11798)
);

CKINVDCx16_ASAP7_75t_R g11799 ( 
.A(n_11559),
.Y(n_11799)
);

NAND2xp5_ASAP7_75t_L g11800 ( 
.A(n_11594),
.B(n_544),
.Y(n_11800)
);

O2A1O1Ixp33_ASAP7_75t_L g11801 ( 
.A1(n_11684),
.A2(n_546),
.B(n_544),
.C(n_545),
.Y(n_11801)
);

A2O1A1Ixp33_ASAP7_75t_SL g11802 ( 
.A1(n_11630),
.A2(n_548),
.B(n_545),
.C(n_547),
.Y(n_11802)
);

BUFx6f_ASAP7_75t_L g11803 ( 
.A(n_11572),
.Y(n_11803)
);

O2A1O1Ixp5_ASAP7_75t_L g11804 ( 
.A1(n_11737),
.A2(n_549),
.B(n_547),
.C(n_548),
.Y(n_11804)
);

INVx4_ASAP7_75t_L g11805 ( 
.A(n_11572),
.Y(n_11805)
);

AOI21xp33_ASAP7_75t_L g11806 ( 
.A1(n_11310),
.A2(n_549),
.B(n_550),
.Y(n_11806)
);

INVx2_ASAP7_75t_L g11807 ( 
.A(n_11328),
.Y(n_11807)
);

INVx1_ASAP7_75t_L g11808 ( 
.A(n_10996),
.Y(n_11808)
);

AO21x2_ASAP7_75t_L g11809 ( 
.A1(n_11678),
.A2(n_550),
.B(n_551),
.Y(n_11809)
);

NAND2xp5_ASAP7_75t_L g11810 ( 
.A(n_11440),
.B(n_551),
.Y(n_11810)
);

NAND2xp5_ASAP7_75t_L g11811 ( 
.A(n_11004),
.B(n_552),
.Y(n_11811)
);

AOI21xp5_ASAP7_75t_L g11812 ( 
.A1(n_11027),
.A2(n_552),
.B(n_553),
.Y(n_11812)
);

AOI21xp5_ASAP7_75t_L g11813 ( 
.A1(n_11006),
.A2(n_553),
.B(n_554),
.Y(n_11813)
);

NAND2xp5_ASAP7_75t_L g11814 ( 
.A(n_11643),
.B(n_554),
.Y(n_11814)
);

NAND2xp5_ASAP7_75t_L g11815 ( 
.A(n_11652),
.B(n_555),
.Y(n_11815)
);

NAND2xp5_ASAP7_75t_L g11816 ( 
.A(n_10998),
.B(n_555),
.Y(n_11816)
);

AOI21xp5_ASAP7_75t_L g11817 ( 
.A1(n_11028),
.A2(n_556),
.B(n_557),
.Y(n_11817)
);

NOR2xp33_ASAP7_75t_R g11818 ( 
.A(n_11366),
.B(n_556),
.Y(n_11818)
);

INVx1_ASAP7_75t_L g11819 ( 
.A(n_11557),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11514),
.B(n_557),
.Y(n_11820)
);

OAI22xp5_ASAP7_75t_L g11821 ( 
.A1(n_11385),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_11821)
);

INVx2_ASAP7_75t_L g11822 ( 
.A(n_10999),
.Y(n_11822)
);

AOI21xp5_ASAP7_75t_L g11823 ( 
.A1(n_10967),
.A2(n_558),
.B(n_559),
.Y(n_11823)
);

AOI21xp5_ASAP7_75t_L g11824 ( 
.A1(n_11554),
.A2(n_561),
.B(n_562),
.Y(n_11824)
);

INVx2_ASAP7_75t_SL g11825 ( 
.A(n_11529),
.Y(n_11825)
);

INVx4_ASAP7_75t_L g11826 ( 
.A(n_11661),
.Y(n_11826)
);

AOI21xp5_ASAP7_75t_L g11827 ( 
.A1(n_11555),
.A2(n_561),
.B(n_562),
.Y(n_11827)
);

AOI21xp5_ASAP7_75t_L g11828 ( 
.A1(n_11577),
.A2(n_563),
.B(n_564),
.Y(n_11828)
);

NAND3xp33_ASAP7_75t_L g11829 ( 
.A(n_11681),
.B(n_565),
.C(n_566),
.Y(n_11829)
);

NOR2x1_ASAP7_75t_R g11830 ( 
.A(n_10981),
.B(n_565),
.Y(n_11830)
);

OAI21xp5_ASAP7_75t_L g11831 ( 
.A1(n_11682),
.A2(n_566),
.B(n_567),
.Y(n_11831)
);

INVx1_ASAP7_75t_L g11832 ( 
.A(n_11571),
.Y(n_11832)
);

AOI22xp33_ASAP7_75t_L g11833 ( 
.A1(n_11042),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_11833)
);

NAND2xp5_ASAP7_75t_SL g11834 ( 
.A(n_11060),
.B(n_568),
.Y(n_11834)
);

NOR2x1p5_ASAP7_75t_SL g11835 ( 
.A(n_11067),
.B(n_569),
.Y(n_11835)
);

BUFx2_ASAP7_75t_SL g11836 ( 
.A(n_11454),
.Y(n_11836)
);

INVx3_ASAP7_75t_L g11837 ( 
.A(n_11115),
.Y(n_11837)
);

AND2x4_ASAP7_75t_L g11838 ( 
.A(n_11466),
.B(n_570),
.Y(n_11838)
);

INVx1_ASAP7_75t_L g11839 ( 
.A(n_11588),
.Y(n_11839)
);

AOI21xp5_ASAP7_75t_L g11840 ( 
.A1(n_11578),
.A2(n_571),
.B(n_573),
.Y(n_11840)
);

CKINVDCx5p33_ASAP7_75t_R g11841 ( 
.A(n_11377),
.Y(n_11841)
);

INVx1_ASAP7_75t_L g11842 ( 
.A(n_11592),
.Y(n_11842)
);

INVx3_ASAP7_75t_L g11843 ( 
.A(n_11529),
.Y(n_11843)
);

AOI22xp5_ASAP7_75t_L g11844 ( 
.A1(n_10982),
.A2(n_574),
.B1(n_571),
.B2(n_573),
.Y(n_11844)
);

O2A1O1Ixp33_ASAP7_75t_L g11845 ( 
.A1(n_11569),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_11845)
);

OAI221xp5_ASAP7_75t_L g11846 ( 
.A1(n_11586),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.C(n_579),
.Y(n_11846)
);

NAND2xp5_ASAP7_75t_L g11847 ( 
.A(n_11600),
.B(n_577),
.Y(n_11847)
);

A2O1A1Ixp33_ASAP7_75t_SL g11848 ( 
.A1(n_10984),
.A2(n_580),
.B(n_578),
.C(n_579),
.Y(n_11848)
);

INVx1_ASAP7_75t_L g11849 ( 
.A(n_11624),
.Y(n_11849)
);

NOR2xp33_ASAP7_75t_SL g11850 ( 
.A(n_11485),
.B(n_581),
.Y(n_11850)
);

INVx4_ASAP7_75t_L g11851 ( 
.A(n_11661),
.Y(n_11851)
);

OAI21xp33_ASAP7_75t_L g11852 ( 
.A1(n_11686),
.A2(n_581),
.B(n_582),
.Y(n_11852)
);

OAI21xp33_ASAP7_75t_L g11853 ( 
.A1(n_11696),
.A2(n_582),
.B(n_583),
.Y(n_11853)
);

OAI22xp5_ASAP7_75t_L g11854 ( 
.A1(n_11078),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_11854)
);

OAI22xp5_ASAP7_75t_L g11855 ( 
.A1(n_11119),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_11855)
);

NAND3xp33_ASAP7_75t_SL g11856 ( 
.A(n_11029),
.B(n_586),
.C(n_587),
.Y(n_11856)
);

NOR2xp33_ASAP7_75t_SL g11857 ( 
.A(n_11299),
.B(n_587),
.Y(n_11857)
);

A2O1A1Ixp33_ASAP7_75t_L g11858 ( 
.A1(n_11714),
.A2(n_590),
.B(n_588),
.C(n_589),
.Y(n_11858)
);

INVx1_ASAP7_75t_L g11859 ( 
.A(n_11639),
.Y(n_11859)
);

BUFx6f_ASAP7_75t_L g11860 ( 
.A(n_11713),
.Y(n_11860)
);

A2O1A1Ixp33_ASAP7_75t_L g11861 ( 
.A1(n_11716),
.A2(n_591),
.B(n_588),
.C(n_590),
.Y(n_11861)
);

INVx1_ASAP7_75t_L g11862 ( 
.A(n_11656),
.Y(n_11862)
);

INVx2_ASAP7_75t_L g11863 ( 
.A(n_11007),
.Y(n_11863)
);

INVx2_ASAP7_75t_L g11864 ( 
.A(n_11024),
.Y(n_11864)
);

AOI21xp5_ASAP7_75t_L g11865 ( 
.A1(n_11581),
.A2(n_591),
.B(n_592),
.Y(n_11865)
);

NOR2xp33_ASAP7_75t_L g11866 ( 
.A(n_11632),
.B(n_592),
.Y(n_11866)
);

A2O1A1Ixp33_ASAP7_75t_L g11867 ( 
.A1(n_11718),
.A2(n_596),
.B(n_593),
.C(n_594),
.Y(n_11867)
);

BUFx2_ASAP7_75t_L g11868 ( 
.A(n_11445),
.Y(n_11868)
);

NAND2xp5_ASAP7_75t_SL g11869 ( 
.A(n_11183),
.B(n_593),
.Y(n_11869)
);

NAND3xp33_ASAP7_75t_SL g11870 ( 
.A(n_11126),
.B(n_594),
.C(n_596),
.Y(n_11870)
);

OAI22xp5_ASAP7_75t_L g11871 ( 
.A1(n_11406),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_11871)
);

BUFx6f_ASAP7_75t_L g11872 ( 
.A(n_11713),
.Y(n_11872)
);

BUFx2_ASAP7_75t_L g11873 ( 
.A(n_11747),
.Y(n_11873)
);

OA22x2_ASAP7_75t_L g11874 ( 
.A1(n_11023),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_11874)
);

INVxp67_ASAP7_75t_L g11875 ( 
.A(n_11066),
.Y(n_11875)
);

NOR2xp33_ASAP7_75t_L g11876 ( 
.A(n_11655),
.B(n_601),
.Y(n_11876)
);

AOI21xp5_ASAP7_75t_L g11877 ( 
.A1(n_11582),
.A2(n_601),
.B(n_602),
.Y(n_11877)
);

INVx2_ASAP7_75t_L g11878 ( 
.A(n_11035),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11675),
.Y(n_11879)
);

BUFx6f_ASAP7_75t_L g11880 ( 
.A(n_11742),
.Y(n_11880)
);

AOI21xp5_ASAP7_75t_L g11881 ( 
.A1(n_11584),
.A2(n_602),
.B(n_603),
.Y(n_11881)
);

AO22x1_ASAP7_75t_L g11882 ( 
.A1(n_11021),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_11882)
);

INVx2_ASAP7_75t_L g11883 ( 
.A(n_11041),
.Y(n_11883)
);

INVx1_ASAP7_75t_L g11884 ( 
.A(n_11694),
.Y(n_11884)
);

INVx2_ASAP7_75t_L g11885 ( 
.A(n_11052),
.Y(n_11885)
);

INVx4_ASAP7_75t_L g11886 ( 
.A(n_11742),
.Y(n_11886)
);

INVx2_ASAP7_75t_L g11887 ( 
.A(n_11096),
.Y(n_11887)
);

A2O1A1Ixp33_ASAP7_75t_L g11888 ( 
.A1(n_11727),
.A2(n_607),
.B(n_604),
.C(n_606),
.Y(n_11888)
);

INVx1_ASAP7_75t_L g11889 ( 
.A(n_11703),
.Y(n_11889)
);

BUFx8_ASAP7_75t_L g11890 ( 
.A(n_11699),
.Y(n_11890)
);

NAND2xp5_ASAP7_75t_SL g11891 ( 
.A(n_11183),
.B(n_606),
.Y(n_11891)
);

O2A1O1Ixp33_ASAP7_75t_L g11892 ( 
.A1(n_11680),
.A2(n_609),
.B(n_607),
.C(n_608),
.Y(n_11892)
);

AOI21xp5_ASAP7_75t_L g11893 ( 
.A1(n_11587),
.A2(n_608),
.B(n_609),
.Y(n_11893)
);

INVx2_ASAP7_75t_L g11894 ( 
.A(n_11112),
.Y(n_11894)
);

OAI22xp5_ASAP7_75t_L g11895 ( 
.A1(n_11194),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.Y(n_11895)
);

OR2x6_ASAP7_75t_SL g11896 ( 
.A(n_11237),
.B(n_611),
.Y(n_11896)
);

NOR3xp33_ASAP7_75t_SL g11897 ( 
.A(n_11109),
.B(n_612),
.C(n_613),
.Y(n_11897)
);

OR2x6_ASAP7_75t_L g11898 ( 
.A(n_10968),
.B(n_613),
.Y(n_11898)
);

OAI21x1_ASAP7_75t_L g11899 ( 
.A1(n_11120),
.A2(n_614),
.B(n_615),
.Y(n_11899)
);

INVx2_ASAP7_75t_SL g11900 ( 
.A(n_11235),
.Y(n_11900)
);

CKINVDCx5p33_ASAP7_75t_R g11901 ( 
.A(n_11018),
.Y(n_11901)
);

NOR2xp33_ASAP7_75t_L g11902 ( 
.A(n_11679),
.B(n_614),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_11721),
.Y(n_11903)
);

AOI21xp5_ASAP7_75t_L g11904 ( 
.A1(n_11589),
.A2(n_11601),
.B(n_11595),
.Y(n_11904)
);

O2A1O1Ixp33_ASAP7_75t_L g11905 ( 
.A1(n_11690),
.A2(n_617),
.B(n_615),
.C(n_616),
.Y(n_11905)
);

INVx5_ASAP7_75t_L g11906 ( 
.A(n_11294),
.Y(n_11906)
);

INVx2_ASAP7_75t_L g11907 ( 
.A(n_11123),
.Y(n_11907)
);

OAI22x1_ASAP7_75t_L g11908 ( 
.A1(n_11723),
.A2(n_619),
.B1(n_616),
.B2(n_618),
.Y(n_11908)
);

INVx2_ASAP7_75t_L g11909 ( 
.A(n_11132),
.Y(n_11909)
);

AOI21xp5_ASAP7_75t_L g11910 ( 
.A1(n_11608),
.A2(n_618),
.B(n_619),
.Y(n_11910)
);

NOR2xp33_ASAP7_75t_L g11911 ( 
.A(n_11216),
.B(n_620),
.Y(n_11911)
);

AOI21xp5_ASAP7_75t_L g11912 ( 
.A1(n_11617),
.A2(n_11633),
.B(n_11621),
.Y(n_11912)
);

AND2x4_ASAP7_75t_L g11913 ( 
.A(n_11436),
.B(n_621),
.Y(n_11913)
);

NAND2xp5_ASAP7_75t_SL g11914 ( 
.A(n_11183),
.B(n_11224),
.Y(n_11914)
);

BUFx3_ASAP7_75t_L g11915 ( 
.A(n_11130),
.Y(n_11915)
);

NOR2xp33_ASAP7_75t_L g11916 ( 
.A(n_11038),
.B(n_622),
.Y(n_11916)
);

BUFx2_ASAP7_75t_L g11917 ( 
.A(n_11475),
.Y(n_11917)
);

CKINVDCx5p33_ASAP7_75t_R g11918 ( 
.A(n_11596),
.Y(n_11918)
);

HB1xp67_ASAP7_75t_L g11919 ( 
.A(n_11405),
.Y(n_11919)
);

OA22x2_ASAP7_75t_L g11920 ( 
.A1(n_11657),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_11920)
);

AOI22xp5_ASAP7_75t_L g11921 ( 
.A1(n_11306),
.A2(n_625),
.B1(n_623),
.B2(n_624),
.Y(n_11921)
);

AOI21xp5_ASAP7_75t_L g11922 ( 
.A1(n_11635),
.A2(n_625),
.B(n_626),
.Y(n_11922)
);

AO32x1_ASAP7_75t_L g11923 ( 
.A1(n_10997),
.A2(n_628),
.A3(n_626),
.B1(n_627),
.B2(n_629),
.Y(n_11923)
);

INVxp67_ASAP7_75t_L g11924 ( 
.A(n_11402),
.Y(n_11924)
);

NAND2xp33_ASAP7_75t_SL g11925 ( 
.A(n_11741),
.B(n_629),
.Y(n_11925)
);

O2A1O1Ixp33_ASAP7_75t_L g11926 ( 
.A1(n_11637),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_11926)
);

AOI21xp5_ASAP7_75t_L g11927 ( 
.A1(n_11640),
.A2(n_630),
.B(n_631),
.Y(n_11927)
);

NOR2xp33_ASAP7_75t_L g11928 ( 
.A(n_11531),
.B(n_632),
.Y(n_11928)
);

NAND2xp5_ASAP7_75t_SL g11929 ( 
.A(n_11224),
.B(n_633),
.Y(n_11929)
);

OAI22xp5_ASAP7_75t_L g11930 ( 
.A1(n_11662),
.A2(n_636),
.B1(n_633),
.B2(n_634),
.Y(n_11930)
);

AOI21xp5_ASAP7_75t_L g11931 ( 
.A1(n_11648),
.A2(n_634),
.B(n_637),
.Y(n_11931)
);

NAND2xp5_ASAP7_75t_SL g11932 ( 
.A(n_11224),
.B(n_637),
.Y(n_11932)
);

NAND2x1_ASAP7_75t_L g11933 ( 
.A(n_11380),
.B(n_638),
.Y(n_11933)
);

INVx2_ASAP7_75t_L g11934 ( 
.A(n_11134),
.Y(n_11934)
);

OAI21xp33_ASAP7_75t_L g11935 ( 
.A1(n_11732),
.A2(n_11735),
.B(n_11733),
.Y(n_11935)
);

OAI22xp5_ASAP7_75t_SL g11936 ( 
.A1(n_11269),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11740),
.Y(n_11937)
);

NOR2xp67_ASAP7_75t_SL g11938 ( 
.A(n_11710),
.B(n_639),
.Y(n_11938)
);

A2O1A1Ixp33_ASAP7_75t_SL g11939 ( 
.A1(n_11743),
.A2(n_11751),
.B(n_11746),
.C(n_11162),
.Y(n_11939)
);

BUFx6f_ASAP7_75t_L g11940 ( 
.A(n_11736),
.Y(n_11940)
);

AOI21xp5_ASAP7_75t_L g11941 ( 
.A1(n_11649),
.A2(n_11660),
.B(n_11658),
.Y(n_11941)
);

NOR2xp33_ASAP7_75t_L g11942 ( 
.A(n_11118),
.B(n_641),
.Y(n_11942)
);

NAND2xp5_ASAP7_75t_L g11943 ( 
.A(n_11071),
.B(n_641),
.Y(n_11943)
);

NAND2xp5_ASAP7_75t_SL g11944 ( 
.A(n_11089),
.B(n_642),
.Y(n_11944)
);

HB1xp67_ASAP7_75t_L g11945 ( 
.A(n_11062),
.Y(n_11945)
);

AOI222xp33_ASAP7_75t_L g11946 ( 
.A1(n_11167),
.A2(n_644),
.B1(n_646),
.B2(n_642),
.C1(n_643),
.C2(n_645),
.Y(n_11946)
);

NAND2xp5_ASAP7_75t_L g11947 ( 
.A(n_10990),
.B(n_644),
.Y(n_11947)
);

O2A1O1Ixp33_ASAP7_75t_SL g11948 ( 
.A1(n_11043),
.A2(n_648),
.B(n_646),
.C(n_647),
.Y(n_11948)
);

INVx1_ASAP7_75t_SL g11949 ( 
.A(n_11212),
.Y(n_11949)
);

NAND2xp5_ASAP7_75t_L g11950 ( 
.A(n_11298),
.B(n_647),
.Y(n_11950)
);

NOR2xp33_ASAP7_75t_L g11951 ( 
.A(n_11056),
.B(n_648),
.Y(n_11951)
);

INVx2_ASAP7_75t_L g11952 ( 
.A(n_11164),
.Y(n_11952)
);

INVx2_ASAP7_75t_L g11953 ( 
.A(n_11170),
.Y(n_11953)
);

NAND2xp5_ASAP7_75t_SL g11954 ( 
.A(n_11541),
.B(n_649),
.Y(n_11954)
);

AOI21xp5_ASAP7_75t_L g11955 ( 
.A1(n_11664),
.A2(n_650),
.B(n_651),
.Y(n_11955)
);

NOR2xp33_ASAP7_75t_SL g11956 ( 
.A(n_11563),
.B(n_650),
.Y(n_11956)
);

AOI22xp5_ASAP7_75t_L g11957 ( 
.A1(n_11059),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.Y(n_11957)
);

O2A1O1Ixp33_ASAP7_75t_L g11958 ( 
.A1(n_11093),
.A2(n_655),
.B(n_652),
.C(n_654),
.Y(n_11958)
);

CKINVDCx5p33_ASAP7_75t_R g11959 ( 
.A(n_11262),
.Y(n_11959)
);

AND2x2_ASAP7_75t_L g11960 ( 
.A(n_11527),
.B(n_654),
.Y(n_11960)
);

OAI21xp5_ASAP7_75t_L g11961 ( 
.A1(n_11665),
.A2(n_655),
.B(n_656),
.Y(n_11961)
);

AO32x1_ASAP7_75t_L g11962 ( 
.A1(n_11614),
.A2(n_658),
.A3(n_656),
.B1(n_657),
.B2(n_659),
.Y(n_11962)
);

BUFx3_ASAP7_75t_L g11963 ( 
.A(n_11130),
.Y(n_11963)
);

AOI21xp5_ASAP7_75t_L g11964 ( 
.A1(n_11667),
.A2(n_657),
.B(n_658),
.Y(n_11964)
);

NOR2xp33_ASAP7_75t_R g11965 ( 
.A(n_11462),
.B(n_659),
.Y(n_11965)
);

CKINVDCx10_ASAP7_75t_R g11966 ( 
.A(n_11031),
.Y(n_11966)
);

NAND2xp5_ASAP7_75t_SL g11967 ( 
.A(n_11239),
.B(n_660),
.Y(n_11967)
);

NAND2xp5_ASAP7_75t_L g11968 ( 
.A(n_11279),
.B(n_660),
.Y(n_11968)
);

NAND2xp5_ASAP7_75t_L g11969 ( 
.A(n_11400),
.B(n_661),
.Y(n_11969)
);

AOI21xp5_ASAP7_75t_L g11970 ( 
.A1(n_11669),
.A2(n_661),
.B(n_662),
.Y(n_11970)
);

NAND2xp5_ASAP7_75t_L g11971 ( 
.A(n_11443),
.B(n_663),
.Y(n_11971)
);

OA21x2_ASAP7_75t_L g11972 ( 
.A1(n_11748),
.A2(n_663),
.B(n_664),
.Y(n_11972)
);

NAND2xp5_ASAP7_75t_L g11973 ( 
.A(n_11452),
.B(n_665),
.Y(n_11973)
);

INVxp67_ASAP7_75t_SL g11974 ( 
.A(n_11308),
.Y(n_11974)
);

INVx1_ASAP7_75t_L g11975 ( 
.A(n_11177),
.Y(n_11975)
);

NAND2xp5_ASAP7_75t_L g11976 ( 
.A(n_11336),
.B(n_666),
.Y(n_11976)
);

AOI21x1_ASAP7_75t_L g11977 ( 
.A1(n_11394),
.A2(n_667),
.B(n_668),
.Y(n_11977)
);

INVx1_ASAP7_75t_L g11978 ( 
.A(n_11182),
.Y(n_11978)
);

AOI21xp5_ASAP7_75t_L g11979 ( 
.A1(n_10970),
.A2(n_11616),
.B(n_11558),
.Y(n_11979)
);

NAND2xp5_ASAP7_75t_L g11980 ( 
.A(n_11255),
.B(n_667),
.Y(n_11980)
);

OR2x6_ASAP7_75t_L g11981 ( 
.A(n_11031),
.B(n_11651),
.Y(n_11981)
);

NAND2xp5_ASAP7_75t_SL g11982 ( 
.A(n_11351),
.B(n_668),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_11205),
.Y(n_11983)
);

NOR2xp33_ASAP7_75t_L g11984 ( 
.A(n_11102),
.B(n_669),
.Y(n_11984)
);

AOI21xp5_ASAP7_75t_L g11985 ( 
.A1(n_11674),
.A2(n_669),
.B(n_670),
.Y(n_11985)
);

CKINVDCx20_ASAP7_75t_R g11986 ( 
.A(n_11322),
.Y(n_11986)
);

OAI22xp5_ASAP7_75t_L g11987 ( 
.A1(n_11314),
.A2(n_673),
.B1(n_671),
.B2(n_672),
.Y(n_11987)
);

O2A1O1Ixp5_ASAP7_75t_L g11988 ( 
.A1(n_11009),
.A2(n_674),
.B(n_672),
.C(n_673),
.Y(n_11988)
);

INVx1_ASAP7_75t_L g11989 ( 
.A(n_11221),
.Y(n_11989)
);

O2A1O1Ixp33_ASAP7_75t_L g11990 ( 
.A1(n_11072),
.A2(n_676),
.B(n_674),
.C(n_675),
.Y(n_11990)
);

OAI21xp33_ASAP7_75t_SL g11991 ( 
.A1(n_11609),
.A2(n_675),
.B(n_676),
.Y(n_11991)
);

NAND2xp5_ASAP7_75t_L g11992 ( 
.A(n_10987),
.B(n_677),
.Y(n_11992)
);

OAI21xp5_ASAP7_75t_L g11993 ( 
.A1(n_11346),
.A2(n_678),
.B(n_679),
.Y(n_11993)
);

AOI21xp5_ASAP7_75t_L g11994 ( 
.A1(n_11070),
.A2(n_678),
.B(n_679),
.Y(n_11994)
);

NAND2xp5_ASAP7_75t_SL g11995 ( 
.A(n_11465),
.B(n_680),
.Y(n_11995)
);

NOR2xp33_ASAP7_75t_L g11996 ( 
.A(n_11055),
.B(n_680),
.Y(n_11996)
);

AOI21xp5_ASAP7_75t_L g11997 ( 
.A1(n_11605),
.A2(n_681),
.B(n_682),
.Y(n_11997)
);

INVx1_ASAP7_75t_L g11998 ( 
.A(n_11222),
.Y(n_11998)
);

AOI21xp5_ASAP7_75t_L g11999 ( 
.A1(n_11165),
.A2(n_681),
.B(n_682),
.Y(n_11999)
);

INVx1_ASAP7_75t_L g12000 ( 
.A(n_11228),
.Y(n_12000)
);

OR2x6_ASAP7_75t_L g12001 ( 
.A(n_11651),
.B(n_683),
.Y(n_12001)
);

NAND2xp5_ASAP7_75t_SL g12002 ( 
.A(n_10972),
.B(n_683),
.Y(n_12002)
);

A2O1A1Ixp33_ASAP7_75t_L g12003 ( 
.A1(n_11073),
.A2(n_686),
.B(n_684),
.C(n_685),
.Y(n_12003)
);

NAND3xp33_ASAP7_75t_L g12004 ( 
.A(n_11160),
.B(n_684),
.C(n_685),
.Y(n_12004)
);

OR2x2_ASAP7_75t_L g12005 ( 
.A(n_11231),
.B(n_686),
.Y(n_12005)
);

INVx1_ASAP7_75t_L g12006 ( 
.A(n_10989),
.Y(n_12006)
);

NAND2xp5_ASAP7_75t_L g12007 ( 
.A(n_11017),
.B(n_687),
.Y(n_12007)
);

AOI22xp33_ASAP7_75t_L g12008 ( 
.A1(n_11254),
.A2(n_11280),
.B1(n_11256),
.B2(n_11179),
.Y(n_12008)
);

NAND2xp33_ASAP7_75t_SL g12009 ( 
.A(n_11069),
.B(n_687),
.Y(n_12009)
);

O2A1O1Ixp33_ASAP7_75t_L g12010 ( 
.A1(n_11044),
.A2(n_690),
.B(n_688),
.C(n_689),
.Y(n_12010)
);

INVx1_ASAP7_75t_L g12011 ( 
.A(n_11057),
.Y(n_12011)
);

NAND2xp5_ASAP7_75t_L g12012 ( 
.A(n_11074),
.B(n_688),
.Y(n_12012)
);

OAI22xp5_ASAP7_75t_SL g12013 ( 
.A1(n_11368),
.A2(n_692),
.B1(n_690),
.B2(n_691),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_11110),
.Y(n_12014)
);

INVx2_ASAP7_75t_L g12015 ( 
.A(n_11143),
.Y(n_12015)
);

NOR2xp33_ASAP7_75t_L g12016 ( 
.A(n_10983),
.B(n_692),
.Y(n_12016)
);

NOR2xp33_ASAP7_75t_L g12017 ( 
.A(n_11026),
.B(n_693),
.Y(n_12017)
);

INVx1_ASAP7_75t_L g12018 ( 
.A(n_11154),
.Y(n_12018)
);

AOI21xp5_ASAP7_75t_L g12019 ( 
.A1(n_11220),
.A2(n_694),
.B(n_695),
.Y(n_12019)
);

AOI21xp5_ASAP7_75t_L g12020 ( 
.A1(n_11504),
.A2(n_694),
.B(n_695),
.Y(n_12020)
);

NOR2xp33_ASAP7_75t_L g12021 ( 
.A(n_11399),
.B(n_696),
.Y(n_12021)
);

NAND2xp5_ASAP7_75t_L g12022 ( 
.A(n_11184),
.B(n_697),
.Y(n_12022)
);

NAND3xp33_ASAP7_75t_SL g12023 ( 
.A(n_11193),
.B(n_697),
.C(n_698),
.Y(n_12023)
);

O2A1O1Ixp33_ASAP7_75t_SL g12024 ( 
.A1(n_11113),
.A2(n_701),
.B(n_699),
.C(n_700),
.Y(n_12024)
);

NOR2xp33_ASAP7_75t_L g12025 ( 
.A(n_11403),
.B(n_699),
.Y(n_12025)
);

AOI21xp5_ASAP7_75t_L g12026 ( 
.A1(n_10985),
.A2(n_700),
.B(n_701),
.Y(n_12026)
);

A2O1A1Ixp33_ASAP7_75t_L g12027 ( 
.A1(n_11039),
.A2(n_704),
.B(n_702),
.C(n_703),
.Y(n_12027)
);

AOI22xp33_ASAP7_75t_L g12028 ( 
.A1(n_11495),
.A2(n_705),
.B1(n_702),
.B2(n_703),
.Y(n_12028)
);

AOI21xp5_ASAP7_75t_L g12029 ( 
.A1(n_11153),
.A2(n_705),
.B(n_706),
.Y(n_12029)
);

AOI21xp5_ASAP7_75t_L g12030 ( 
.A1(n_10992),
.A2(n_706),
.B(n_707),
.Y(n_12030)
);

NOR2xp33_ASAP7_75t_L g12031 ( 
.A(n_11297),
.B(n_707),
.Y(n_12031)
);

NAND2xp5_ASAP7_75t_L g12032 ( 
.A(n_11185),
.B(n_708),
.Y(n_12032)
);

OAI21xp33_ASAP7_75t_SL g12033 ( 
.A1(n_11459),
.A2(n_709),
.B(n_710),
.Y(n_12033)
);

INVx2_ASAP7_75t_L g12034 ( 
.A(n_11190),
.Y(n_12034)
);

NAND2xp5_ASAP7_75t_SL g12035 ( 
.A(n_11124),
.B(n_709),
.Y(n_12035)
);

CKINVDCx6p67_ASAP7_75t_R g12036 ( 
.A(n_11709),
.Y(n_12036)
);

BUFx6f_ASAP7_75t_L g12037 ( 
.A(n_10969),
.Y(n_12037)
);

AOI21xp5_ASAP7_75t_L g12038 ( 
.A1(n_11092),
.A2(n_710),
.B(n_711),
.Y(n_12038)
);

OAI22x1_ASAP7_75t_L g12039 ( 
.A1(n_11539),
.A2(n_713),
.B1(n_711),
.B2(n_712),
.Y(n_12039)
);

O2A1O1Ixp33_ASAP7_75t_L g12040 ( 
.A1(n_11331),
.A2(n_716),
.B(n_713),
.C(n_714),
.Y(n_12040)
);

AND2x2_ASAP7_75t_L g12041 ( 
.A(n_11441),
.B(n_714),
.Y(n_12041)
);

CKINVDCx20_ASAP7_75t_R g12042 ( 
.A(n_11376),
.Y(n_12042)
);

NOR3xp33_ASAP7_75t_L g12043 ( 
.A(n_11019),
.B(n_716),
.C(n_717),
.Y(n_12043)
);

OR2x2_ASAP7_75t_SL g12044 ( 
.A(n_11345),
.B(n_717),
.Y(n_12044)
);

NAND2xp5_ASAP7_75t_L g12045 ( 
.A(n_11195),
.B(n_11217),
.Y(n_12045)
);

AOI21xp5_ASAP7_75t_L g12046 ( 
.A1(n_11288),
.A2(n_718),
.B(n_719),
.Y(n_12046)
);

NOR3xp33_ASAP7_75t_L g12047 ( 
.A(n_11343),
.B(n_718),
.C(n_720),
.Y(n_12047)
);

INVx5_ASAP7_75t_L g12048 ( 
.A(n_11416),
.Y(n_12048)
);

CKINVDCx20_ASAP7_75t_R g12049 ( 
.A(n_11534),
.Y(n_12049)
);

BUFx6f_ASAP7_75t_L g12050 ( 
.A(n_11146),
.Y(n_12050)
);

AOI22xp5_ASAP7_75t_L g12051 ( 
.A1(n_11152),
.A2(n_11225),
.B1(n_11244),
.B2(n_11196),
.Y(n_12051)
);

AOI21xp5_ASAP7_75t_L g12052 ( 
.A1(n_10988),
.A2(n_720),
.B(n_721),
.Y(n_12052)
);

AOI21xp5_ASAP7_75t_L g12053 ( 
.A1(n_11008),
.A2(n_11415),
.B(n_11414),
.Y(n_12053)
);

INVx2_ASAP7_75t_L g12054 ( 
.A(n_11603),
.Y(n_12054)
);

NOR2xp33_ASAP7_75t_L g12055 ( 
.A(n_11094),
.B(n_721),
.Y(n_12055)
);

A2O1A1Ixp33_ASAP7_75t_L g12056 ( 
.A1(n_11223),
.A2(n_724),
.B(n_722),
.C(n_723),
.Y(n_12056)
);

INVx2_ASAP7_75t_L g12057 ( 
.A(n_11620),
.Y(n_12057)
);

BUFx3_ASAP7_75t_L g12058 ( 
.A(n_11173),
.Y(n_12058)
);

AOI22xp5_ASAP7_75t_L g12059 ( 
.A1(n_11270),
.A2(n_724),
.B1(n_722),
.B2(n_723),
.Y(n_12059)
);

INVx2_ASAP7_75t_L g12060 ( 
.A(n_11626),
.Y(n_12060)
);

INVx3_ASAP7_75t_L g12061 ( 
.A(n_11339),
.Y(n_12061)
);

INVx1_ASAP7_75t_L g12062 ( 
.A(n_11641),
.Y(n_12062)
);

INVx1_ASAP7_75t_L g12063 ( 
.A(n_11672),
.Y(n_12063)
);

O2A1O1Ixp33_ASAP7_75t_SL g12064 ( 
.A1(n_11448),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_12064)
);

BUFx8_ASAP7_75t_SL g12065 ( 
.A(n_11169),
.Y(n_12065)
);

INVxp67_ASAP7_75t_SL g12066 ( 
.A(n_11313),
.Y(n_12066)
);

INVxp67_ASAP7_75t_L g12067 ( 
.A(n_11513),
.Y(n_12067)
);

NAND2xp5_ASAP7_75t_L g12068 ( 
.A(n_11685),
.B(n_725),
.Y(n_12068)
);

INVx3_ASAP7_75t_SL g12069 ( 
.A(n_11025),
.Y(n_12069)
);

OAI22xp5_ASAP7_75t_SL g12070 ( 
.A1(n_11424),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_12070)
);

OAI22xp5_ASAP7_75t_L g12071 ( 
.A1(n_11451),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_12071)
);

NAND2xp33_ASAP7_75t_SL g12072 ( 
.A(n_11304),
.B(n_730),
.Y(n_12072)
);

INVx2_ASAP7_75t_L g12073 ( 
.A(n_11695),
.Y(n_12073)
);

AND2x4_ASAP7_75t_L g12074 ( 
.A(n_11384),
.B(n_731),
.Y(n_12074)
);

NOR2xp67_ASAP7_75t_SL g12075 ( 
.A(n_11488),
.B(n_732),
.Y(n_12075)
);

AOI21xp5_ASAP7_75t_L g12076 ( 
.A1(n_10974),
.A2(n_732),
.B(n_733),
.Y(n_12076)
);

AOI22xp5_ASAP7_75t_L g12077 ( 
.A1(n_11273),
.A2(n_735),
.B1(n_733),
.B2(n_734),
.Y(n_12077)
);

NOR2xp33_ASAP7_75t_L g12078 ( 
.A(n_11253),
.B(n_11129),
.Y(n_12078)
);

AND2x6_ASAP7_75t_SL g12079 ( 
.A(n_11720),
.B(n_734),
.Y(n_12079)
);

OAI22xp5_ASAP7_75t_SL g12080 ( 
.A1(n_11438),
.A2(n_737),
.B1(n_735),
.B2(n_736),
.Y(n_12080)
);

AOI21xp5_ASAP7_75t_L g12081 ( 
.A1(n_11492),
.A2(n_736),
.B(n_737),
.Y(n_12081)
);

NAND2xp5_ASAP7_75t_L g12082 ( 
.A(n_11712),
.B(n_11725),
.Y(n_12082)
);

INVx1_ASAP7_75t_L g12083 ( 
.A(n_11302),
.Y(n_12083)
);

OAI21xp5_ASAP7_75t_L g12084 ( 
.A1(n_11350),
.A2(n_738),
.B(n_739),
.Y(n_12084)
);

NAND2xp33_ASAP7_75t_L g12085 ( 
.A(n_11382),
.B(n_738),
.Y(n_12085)
);

NAND2xp5_ASAP7_75t_L g12086 ( 
.A(n_11317),
.B(n_739),
.Y(n_12086)
);

OAI22x1_ASAP7_75t_L g12087 ( 
.A1(n_11104),
.A2(n_742),
.B1(n_740),
.B2(n_741),
.Y(n_12087)
);

AO21x1_ASAP7_75t_L g12088 ( 
.A1(n_11095),
.A2(n_741),
.B(n_742),
.Y(n_12088)
);

NAND2xp5_ASAP7_75t_SL g12089 ( 
.A(n_11562),
.B(n_743),
.Y(n_12089)
);

AOI22xp5_ASAP7_75t_L g12090 ( 
.A1(n_11281),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_12090)
);

BUFx4f_ASAP7_75t_L g12091 ( 
.A(n_11025),
.Y(n_12091)
);

NOR2xp33_ASAP7_75t_R g12092 ( 
.A(n_11211),
.B(n_745),
.Y(n_12092)
);

NAND2xp5_ASAP7_75t_L g12093 ( 
.A(n_11335),
.B(n_746),
.Y(n_12093)
);

OAI22x1_ASAP7_75t_L g12094 ( 
.A1(n_11275),
.A2(n_748),
.B1(n_746),
.B2(n_747),
.Y(n_12094)
);

INVx2_ASAP7_75t_L g12095 ( 
.A(n_11425),
.Y(n_12095)
);

AOI21xp5_ASAP7_75t_L g12096 ( 
.A1(n_11145),
.A2(n_747),
.B(n_748),
.Y(n_12096)
);

INVx1_ASAP7_75t_L g12097 ( 
.A(n_11214),
.Y(n_12097)
);

NOR2xp33_ASAP7_75t_L g12098 ( 
.A(n_11574),
.B(n_749),
.Y(n_12098)
);

INVx2_ASAP7_75t_L g12099 ( 
.A(n_11051),
.Y(n_12099)
);

OR2x2_ASAP7_75t_L g12100 ( 
.A(n_11507),
.B(n_750),
.Y(n_12100)
);

CKINVDCx20_ASAP7_75t_R g12101 ( 
.A(n_11036),
.Y(n_12101)
);

NOR2xp33_ASAP7_75t_L g12102 ( 
.A(n_11575),
.B(n_750),
.Y(n_12102)
);

OAI22xp5_ASAP7_75t_L g12103 ( 
.A1(n_11411),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_12103)
);

INVx6_ASAP7_75t_L g12104 ( 
.A(n_11036),
.Y(n_12104)
);

A2O1A1Ixp33_ASAP7_75t_L g12105 ( 
.A1(n_11395),
.A2(n_753),
.B(n_751),
.C(n_752),
.Y(n_12105)
);

INVx2_ASAP7_75t_L g12106 ( 
.A(n_11498),
.Y(n_12106)
);

INVx1_ASAP7_75t_SL g12107 ( 
.A(n_11491),
.Y(n_12107)
);

HB1xp67_ASAP7_75t_L g12108 ( 
.A(n_11509),
.Y(n_12108)
);

INVx2_ASAP7_75t_L g12109 ( 
.A(n_11107),
.Y(n_12109)
);

AOI21xp5_ASAP7_75t_L g12110 ( 
.A1(n_11151),
.A2(n_754),
.B(n_755),
.Y(n_12110)
);

AOI21xp5_ASAP7_75t_L g12111 ( 
.A1(n_11166),
.A2(n_754),
.B(n_755),
.Y(n_12111)
);

INVx2_ASAP7_75t_L g12112 ( 
.A(n_11702),
.Y(n_12112)
);

INVx2_ASAP7_75t_L g12113 ( 
.A(n_11702),
.Y(n_12113)
);

OAI22x1_ASAP7_75t_L g12114 ( 
.A1(n_11705),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_12114)
);

AOI22xp5_ASAP7_75t_L g12115 ( 
.A1(n_11324),
.A2(n_759),
.B1(n_756),
.B2(n_758),
.Y(n_12115)
);

NOR2xp33_ASAP7_75t_L g12116 ( 
.A(n_11576),
.B(n_759),
.Y(n_12116)
);

AOI21xp5_ASAP7_75t_L g12117 ( 
.A1(n_11172),
.A2(n_760),
.B(n_761),
.Y(n_12117)
);

INVx1_ASAP7_75t_L g12118 ( 
.A(n_11282),
.Y(n_12118)
);

NAND2xp5_ASAP7_75t_SL g12119 ( 
.A(n_10975),
.B(n_760),
.Y(n_12119)
);

INVx1_ASAP7_75t_L g12120 ( 
.A(n_11286),
.Y(n_12120)
);

NOR2xp33_ASAP7_75t_L g12121 ( 
.A(n_11647),
.B(n_761),
.Y(n_12121)
);

INVx1_ASAP7_75t_L g12122 ( 
.A(n_11303),
.Y(n_12122)
);

AOI21xp5_ASAP7_75t_L g12123 ( 
.A1(n_11333),
.A2(n_762),
.B(n_763),
.Y(n_12123)
);

OAI21x1_ASAP7_75t_L g12124 ( 
.A1(n_11606),
.A2(n_762),
.B(n_763),
.Y(n_12124)
);

INVx1_ASAP7_75t_L g12125 ( 
.A(n_11305),
.Y(n_12125)
);

INVx2_ASAP7_75t_L g12126 ( 
.A(n_11311),
.Y(n_12126)
);

INVx2_ASAP7_75t_L g12127 ( 
.A(n_11320),
.Y(n_12127)
);

O2A1O1Ixp33_ASAP7_75t_L g12128 ( 
.A1(n_11301),
.A2(n_766),
.B(n_764),
.C(n_765),
.Y(n_12128)
);

AND2x4_ASAP7_75t_L g12129 ( 
.A(n_11156),
.B(n_767),
.Y(n_12129)
);

NOR3xp33_ASAP7_75t_L g12130 ( 
.A(n_11353),
.B(n_767),
.C(n_768),
.Y(n_12130)
);

NOR2xp33_ASAP7_75t_R g12131 ( 
.A(n_11580),
.B(n_769),
.Y(n_12131)
);

BUFx3_ASAP7_75t_L g12132 ( 
.A(n_11173),
.Y(n_12132)
);

NOR2xp33_ASAP7_75t_L g12133 ( 
.A(n_11369),
.B(n_770),
.Y(n_12133)
);

INVx2_ASAP7_75t_L g12134 ( 
.A(n_11321),
.Y(n_12134)
);

O2A1O1Ixp5_ASAP7_75t_L g12135 ( 
.A1(n_11388),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_12135)
);

INVx4_ASAP7_75t_L g12136 ( 
.A(n_11707),
.Y(n_12136)
);

OR2x2_ASAP7_75t_L g12137 ( 
.A(n_11058),
.B(n_771),
.Y(n_12137)
);

INVx3_ASAP7_75t_L g12138 ( 
.A(n_11198),
.Y(n_12138)
);

OR2x6_ASAP7_75t_L g12139 ( 
.A(n_11373),
.B(n_772),
.Y(n_12139)
);

NAND2xp5_ASAP7_75t_L g12140 ( 
.A(n_11704),
.B(n_773),
.Y(n_12140)
);

AND2x2_ASAP7_75t_L g12141 ( 
.A(n_11708),
.B(n_11144),
.Y(n_12141)
);

NAND2xp5_ASAP7_75t_SL g12142 ( 
.A(n_11599),
.B(n_773),
.Y(n_12142)
);

BUFx6f_ASAP7_75t_L g12143 ( 
.A(n_11198),
.Y(n_12143)
);

OAI22xp5_ASAP7_75t_L g12144 ( 
.A1(n_11450),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_12144)
);

NAND2xp5_ASAP7_75t_SL g12145 ( 
.A(n_11446),
.B(n_774),
.Y(n_12145)
);

NAND2xp5_ASAP7_75t_SL g12146 ( 
.A(n_11047),
.B(n_775),
.Y(n_12146)
);

AOI21x1_ASAP7_75t_L g12147 ( 
.A1(n_11341),
.A2(n_11429),
.B(n_11418),
.Y(n_12147)
);

NAND2xp5_ASAP7_75t_L g12148 ( 
.A(n_10976),
.B(n_776),
.Y(n_12148)
);

OAI22xp5_ASAP7_75t_L g12149 ( 
.A1(n_11434),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.Y(n_12149)
);

INVx1_ASAP7_75t_L g12150 ( 
.A(n_11327),
.Y(n_12150)
);

AO21x1_ASAP7_75t_L g12151 ( 
.A1(n_11638),
.A2(n_777),
.B(n_778),
.Y(n_12151)
);

INVx4_ASAP7_75t_L g12152 ( 
.A(n_11122),
.Y(n_12152)
);

AOI21xp5_ASAP7_75t_L g12153 ( 
.A1(n_11010),
.A2(n_780),
.B(n_781),
.Y(n_12153)
);

A2O1A1Ixp33_ASAP7_75t_L g12154 ( 
.A1(n_11050),
.A2(n_782),
.B(n_780),
.C(n_781),
.Y(n_12154)
);

BUFx2_ASAP7_75t_L g12155 ( 
.A(n_11432),
.Y(n_12155)
);

INVxp67_ASAP7_75t_L g12156 ( 
.A(n_11546),
.Y(n_12156)
);

AOI21xp5_ASAP7_75t_L g12157 ( 
.A1(n_11030),
.A2(n_782),
.B(n_783),
.Y(n_12157)
);

INVx4_ASAP7_75t_L g12158 ( 
.A(n_11243),
.Y(n_12158)
);

O2A1O1Ixp33_ASAP7_75t_L g12159 ( 
.A1(n_11319),
.A2(n_786),
.B(n_784),
.C(n_785),
.Y(n_12159)
);

AOI21xp5_ASAP7_75t_L g12160 ( 
.A1(n_11260),
.A2(n_785),
.B(n_786),
.Y(n_12160)
);

AOI21xp5_ASAP7_75t_L g12161 ( 
.A1(n_11264),
.A2(n_787),
.B(n_788),
.Y(n_12161)
);

AOI21xp5_ASAP7_75t_L g12162 ( 
.A1(n_11325),
.A2(n_787),
.B(n_788),
.Y(n_12162)
);

AOI21xp5_ASAP7_75t_L g12163 ( 
.A1(n_11570),
.A2(n_789),
.B(n_790),
.Y(n_12163)
);

NOR2xp33_ASAP7_75t_L g12164 ( 
.A(n_11149),
.B(n_789),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_11174),
.Y(n_12165)
);

INVx3_ASAP7_75t_L g12166 ( 
.A(n_11549),
.Y(n_12166)
);

AOI21xp5_ASAP7_75t_L g12167 ( 
.A1(n_11611),
.A2(n_791),
.B(n_792),
.Y(n_12167)
);

A2O1A1Ixp33_ASAP7_75t_L g12168 ( 
.A1(n_11240),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_12168)
);

NAND2xp5_ASAP7_75t_L g12169 ( 
.A(n_11560),
.B(n_793),
.Y(n_12169)
);

O2A1O1Ixp33_ASAP7_75t_SL g12170 ( 
.A1(n_11367),
.A2(n_796),
.B(n_794),
.C(n_795),
.Y(n_12170)
);

A2O1A1Ixp33_ASAP7_75t_L g12171 ( 
.A1(n_11277),
.A2(n_797),
.B(n_794),
.C(n_796),
.Y(n_12171)
);

OAI22xp5_ASAP7_75t_L g12172 ( 
.A1(n_11565),
.A2(n_799),
.B1(n_797),
.B2(n_798),
.Y(n_12172)
);

INVx2_ASAP7_75t_L g12173 ( 
.A(n_11203),
.Y(n_12173)
);

O2A1O1Ixp5_ASAP7_75t_L g12174 ( 
.A1(n_11431),
.A2(n_800),
.B(n_798),
.C(n_799),
.Y(n_12174)
);

INVx2_ASAP7_75t_L g12175 ( 
.A(n_11208),
.Y(n_12175)
);

NAND2xp5_ASAP7_75t_L g12176 ( 
.A(n_11566),
.B(n_11567),
.Y(n_12176)
);

INVx4_ASAP7_75t_L g12177 ( 
.A(n_11243),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_11210),
.Y(n_12178)
);

NAND2x1p5_ASAP7_75t_L g12179 ( 
.A(n_11463),
.B(n_800),
.Y(n_12179)
);

CKINVDCx20_ASAP7_75t_R g12180 ( 
.A(n_11455),
.Y(n_12180)
);

NAND2xp5_ASAP7_75t_L g12181 ( 
.A(n_11579),
.B(n_801),
.Y(n_12181)
);

AND2x4_ASAP7_75t_L g12182 ( 
.A(n_11505),
.B(n_801),
.Y(n_12182)
);

OAI22xp5_ASAP7_75t_L g12183 ( 
.A1(n_11687),
.A2(n_805),
.B1(n_802),
.B2(n_804),
.Y(n_12183)
);

BUFx8_ASAP7_75t_L g12184 ( 
.A(n_11668),
.Y(n_12184)
);

INVx1_ASAP7_75t_L g12185 ( 
.A(n_11100),
.Y(n_12185)
);

NAND2xp5_ASAP7_75t_L g12186 ( 
.A(n_11591),
.B(n_802),
.Y(n_12186)
);

BUFx6f_ASAP7_75t_L g12187 ( 
.A(n_11263),
.Y(n_12187)
);

AO22x1_ASAP7_75t_L g12188 ( 
.A1(n_11359),
.A2(n_806),
.B1(n_804),
.B2(n_805),
.Y(n_12188)
);

AND2x4_ASAP7_75t_L g12189 ( 
.A(n_11391),
.B(n_806),
.Y(n_12189)
);

BUFx6f_ASAP7_75t_L g12190 ( 
.A(n_11263),
.Y(n_12190)
);

INVx1_ASAP7_75t_L g12191 ( 
.A(n_11334),
.Y(n_12191)
);

OAI21xp5_ASAP7_75t_L g12192 ( 
.A1(n_11360),
.A2(n_807),
.B(n_808),
.Y(n_12192)
);

A2O1A1Ixp33_ASAP7_75t_L g12193 ( 
.A1(n_11284),
.A2(n_809),
.B(n_807),
.C(n_808),
.Y(n_12193)
);

NOR2x1_ASAP7_75t_L g12194 ( 
.A(n_10980),
.B(n_809),
.Y(n_12194)
);

BUFx6f_ASAP7_75t_L g12195 ( 
.A(n_11381),
.Y(n_12195)
);

AOI221xp5_ASAP7_75t_SL g12196 ( 
.A1(n_11489),
.A2(n_812),
.B1(n_810),
.B2(n_811),
.C(n_813),
.Y(n_12196)
);

AND2x2_ASAP7_75t_L g12197 ( 
.A(n_11014),
.B(n_810),
.Y(n_12197)
);

A2O1A1Ixp33_ASAP7_75t_L g12198 ( 
.A1(n_11285),
.A2(n_814),
.B(n_811),
.C(n_812),
.Y(n_12198)
);

INVx2_ASAP7_75t_SL g12199 ( 
.A(n_11187),
.Y(n_12199)
);

AOI21x1_ASAP7_75t_L g12200 ( 
.A1(n_11227),
.A2(n_814),
.B(n_815),
.Y(n_12200)
);

INVx2_ASAP7_75t_L g12201 ( 
.A(n_11340),
.Y(n_12201)
);

BUFx6f_ASAP7_75t_L g12202 ( 
.A(n_11381),
.Y(n_12202)
);

A2O1A1Ixp33_ASAP7_75t_L g12203 ( 
.A1(n_11347),
.A2(n_817),
.B(n_815),
.C(n_816),
.Y(n_12203)
);

INVx2_ASAP7_75t_SL g12204 ( 
.A(n_11250),
.Y(n_12204)
);

BUFx8_ASAP7_75t_L g12205 ( 
.A(n_11447),
.Y(n_12205)
);

BUFx2_ASAP7_75t_L g12206 ( 
.A(n_11447),
.Y(n_12206)
);

AOI21xp5_ASAP7_75t_L g12207 ( 
.A1(n_11618),
.A2(n_816),
.B(n_818),
.Y(n_12207)
);

NAND2xp5_ASAP7_75t_L g12208 ( 
.A(n_11593),
.B(n_819),
.Y(n_12208)
);

NOR3xp33_ASAP7_75t_L g12209 ( 
.A(n_11393),
.B(n_819),
.C(n_820),
.Y(n_12209)
);

A2O1A1Ixp33_ASAP7_75t_L g12210 ( 
.A1(n_11461),
.A2(n_822),
.B(n_820),
.C(n_821),
.Y(n_12210)
);

NOR3xp33_ASAP7_75t_SL g12211 ( 
.A(n_11500),
.B(n_821),
.C(n_822),
.Y(n_12211)
);

AOI22xp5_ASAP7_75t_L g12212 ( 
.A1(n_11711),
.A2(n_826),
.B1(n_823),
.B2(n_825),
.Y(n_12212)
);

OAI21x1_ASAP7_75t_L g12213 ( 
.A1(n_11706),
.A2(n_823),
.B(n_825),
.Y(n_12213)
);

NAND2xp5_ASAP7_75t_SL g12214 ( 
.A(n_11188),
.B(n_826),
.Y(n_12214)
);

NAND2xp5_ASAP7_75t_SL g12215 ( 
.A(n_11192),
.B(n_827),
.Y(n_12215)
);

AOI21xp5_ASAP7_75t_L g12216 ( 
.A1(n_11338),
.A2(n_827),
.B(n_828),
.Y(n_12216)
);

NAND2xp5_ASAP7_75t_L g12217 ( 
.A(n_11597),
.B(n_828),
.Y(n_12217)
);

NAND2xp5_ASAP7_75t_L g12218 ( 
.A(n_11598),
.B(n_829),
.Y(n_12218)
);

BUFx2_ASAP7_75t_L g12219 ( 
.A(n_11171),
.Y(n_12219)
);

INVx2_ASAP7_75t_L g12220 ( 
.A(n_11344),
.Y(n_12220)
);

NAND2xp5_ASAP7_75t_L g12221 ( 
.A(n_11602),
.B(n_829),
.Y(n_12221)
);

INVx5_ASAP7_75t_L g12222 ( 
.A(n_11416),
.Y(n_12222)
);

A2O1A1Ixp33_ASAP7_75t_L g12223 ( 
.A1(n_11471),
.A2(n_832),
.B(n_830),
.C(n_831),
.Y(n_12223)
);

BUFx12f_ASAP7_75t_L g12224 ( 
.A(n_11583),
.Y(n_12224)
);

INVx1_ASAP7_75t_L g12225 ( 
.A(n_11348),
.Y(n_12225)
);

NAND2xp5_ASAP7_75t_SL g12226 ( 
.A(n_11116),
.B(n_830),
.Y(n_12226)
);

AO32x2_ASAP7_75t_L g12227 ( 
.A1(n_11659),
.A2(n_11688),
.A3(n_11689),
.B1(n_11683),
.B2(n_11671),
.Y(n_12227)
);

INVx3_ASAP7_75t_L g12228 ( 
.A(n_11517),
.Y(n_12228)
);

AND2x4_ASAP7_75t_L g12229 ( 
.A(n_11585),
.B(n_831),
.Y(n_12229)
);

BUFx2_ASAP7_75t_L g12230 ( 
.A(n_11482),
.Y(n_12230)
);

NAND2xp5_ASAP7_75t_SL g12231 ( 
.A(n_11215),
.B(n_832),
.Y(n_12231)
);

AOI21xp5_ASAP7_75t_L g12232 ( 
.A1(n_11175),
.A2(n_833),
.B(n_834),
.Y(n_12232)
);

AND2x2_ASAP7_75t_SL g12233 ( 
.A(n_11079),
.B(n_833),
.Y(n_12233)
);

CKINVDCx8_ASAP7_75t_R g12234 ( 
.A(n_11726),
.Y(n_12234)
);

AOI21xp5_ASAP7_75t_L g12235 ( 
.A1(n_11176),
.A2(n_834),
.B(n_835),
.Y(n_12235)
);

A2O1A1Ixp33_ASAP7_75t_L g12236 ( 
.A1(n_11121),
.A2(n_838),
.B(n_836),
.C(n_837),
.Y(n_12236)
);

OR2x6_ASAP7_75t_L g12237 ( 
.A(n_11001),
.B(n_836),
.Y(n_12237)
);

NAND2xp5_ASAP7_75t_L g12238 ( 
.A(n_11604),
.B(n_837),
.Y(n_12238)
);

NAND2xp5_ASAP7_75t_SL g12239 ( 
.A(n_11141),
.B(n_839),
.Y(n_12239)
);

AOI21x1_ASAP7_75t_L g12240 ( 
.A1(n_11090),
.A2(n_839),
.B(n_840),
.Y(n_12240)
);

INVxp67_ASAP7_75t_L g12241 ( 
.A(n_11103),
.Y(n_12241)
);

A2O1A1Ixp33_ASAP7_75t_L g12242 ( 
.A1(n_11508),
.A2(n_842),
.B(n_840),
.C(n_841),
.Y(n_12242)
);

NOR2xp67_ASAP7_75t_L g12243 ( 
.A(n_10993),
.B(n_11003),
.Y(n_12243)
);

BUFx6f_ASAP7_75t_L g12244 ( 
.A(n_11326),
.Y(n_12244)
);

NAND2xp5_ASAP7_75t_L g12245 ( 
.A(n_11607),
.B(n_841),
.Y(n_12245)
);

OA21x2_ASAP7_75t_L g12246 ( 
.A1(n_11734),
.A2(n_842),
.B(n_843),
.Y(n_12246)
);

OAI22xp5_ASAP7_75t_L g12247 ( 
.A1(n_11715),
.A2(n_11738),
.B1(n_11449),
.B2(n_11261),
.Y(n_12247)
);

O2A1O1Ixp33_ASAP7_75t_L g12248 ( 
.A1(n_11186),
.A2(n_846),
.B(n_844),
.C(n_845),
.Y(n_12248)
);

BUFx2_ASAP7_75t_L g12249 ( 
.A(n_11416),
.Y(n_12249)
);

NAND2xp5_ASAP7_75t_L g12250 ( 
.A(n_11612),
.B(n_844),
.Y(n_12250)
);

AOI21xp5_ASAP7_75t_L g12251 ( 
.A1(n_11159),
.A2(n_11140),
.B(n_11131),
.Y(n_12251)
);

INVx1_ASAP7_75t_L g12252 ( 
.A(n_11354),
.Y(n_12252)
);

AOI21x1_ASAP7_75t_L g12253 ( 
.A1(n_11232),
.A2(n_845),
.B(n_846),
.Y(n_12253)
);

INVx8_ASAP7_75t_L g12254 ( 
.A(n_11515),
.Y(n_12254)
);

NOR2xp33_ASAP7_75t_L g12255 ( 
.A(n_11168),
.B(n_847),
.Y(n_12255)
);

INVx1_ASAP7_75t_L g12256 ( 
.A(n_11356),
.Y(n_12256)
);

O2A1O1Ixp33_ASAP7_75t_L g12257 ( 
.A1(n_11300),
.A2(n_849),
.B(n_847),
.C(n_848),
.Y(n_12257)
);

AOI22xp33_ASAP7_75t_L g12258 ( 
.A1(n_11412),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_12258)
);

AOI21xp5_ASAP7_75t_L g12259 ( 
.A1(n_11408),
.A2(n_850),
.B(n_851),
.Y(n_12259)
);

O2A1O1Ixp5_ASAP7_75t_L g12260 ( 
.A1(n_11691),
.A2(n_854),
.B(n_852),
.C(n_853),
.Y(n_12260)
);

INVx1_ASAP7_75t_L g12261 ( 
.A(n_11358),
.Y(n_12261)
);

AOI22xp5_ASAP7_75t_L g12262 ( 
.A1(n_11075),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.Y(n_12262)
);

NOR2xp33_ASAP7_75t_L g12263 ( 
.A(n_11191),
.B(n_855),
.Y(n_12263)
);

NAND2xp5_ASAP7_75t_SL g12264 ( 
.A(n_11258),
.B(n_855),
.Y(n_12264)
);

INVx1_ASAP7_75t_L g12265 ( 
.A(n_11049),
.Y(n_12265)
);

AND2x4_ASAP7_75t_L g12266 ( 
.A(n_11423),
.B(n_856),
.Y(n_12266)
);

NAND2xp5_ASAP7_75t_L g12267 ( 
.A(n_11623),
.B(n_856),
.Y(n_12267)
);

NOR2xp67_ASAP7_75t_L g12268 ( 
.A(n_11013),
.B(n_857),
.Y(n_12268)
);

NOR2xp33_ASAP7_75t_R g12269 ( 
.A(n_11744),
.B(n_857),
.Y(n_12269)
);

AOI21xp5_ASAP7_75t_L g12270 ( 
.A1(n_11233),
.A2(n_858),
.B(n_859),
.Y(n_12270)
);

NAND2xp5_ASAP7_75t_SL g12271 ( 
.A(n_11147),
.B(n_858),
.Y(n_12271)
);

NOR2xp67_ASAP7_75t_L g12272 ( 
.A(n_11016),
.B(n_859),
.Y(n_12272)
);

INVx5_ASAP7_75t_L g12273 ( 
.A(n_11080),
.Y(n_12273)
);

AOI21xp5_ASAP7_75t_L g12274 ( 
.A1(n_11234),
.A2(n_860),
.B(n_861),
.Y(n_12274)
);

BUFx2_ASAP7_75t_SL g12275 ( 
.A(n_11724),
.Y(n_12275)
);

OAI22x1_ASAP7_75t_L g12276 ( 
.A1(n_11467),
.A2(n_863),
.B1(n_860),
.B2(n_862),
.Y(n_12276)
);

INVx1_ASAP7_75t_L g12277 ( 
.A(n_11061),
.Y(n_12277)
);

AOI21xp5_ASAP7_75t_L g12278 ( 
.A1(n_11238),
.A2(n_862),
.B(n_864),
.Y(n_12278)
);

INVx1_ASAP7_75t_L g12279 ( 
.A(n_11077),
.Y(n_12279)
);

AND2x2_ASAP7_75t_L g12280 ( 
.A(n_11568),
.B(n_864),
.Y(n_12280)
);

OAI22xp33_ASAP7_75t_L g12281 ( 
.A1(n_11473),
.A2(n_11439),
.B1(n_11442),
.B2(n_11430),
.Y(n_12281)
);

NOR2x1_ASAP7_75t_L g12282 ( 
.A(n_11088),
.B(n_865),
.Y(n_12282)
);

INVx2_ASAP7_75t_L g12283 ( 
.A(n_11083),
.Y(n_12283)
);

BUFx6f_ASAP7_75t_L g12284 ( 
.A(n_11207),
.Y(n_12284)
);

OAI22xp5_ASAP7_75t_L g12285 ( 
.A1(n_11287),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_12285)
);

NOR3xp33_ASAP7_75t_SL g12286 ( 
.A(n_11476),
.B(n_866),
.C(n_867),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_11033),
.Y(n_12287)
);

NOR2xp33_ASAP7_75t_L g12288 ( 
.A(n_11352),
.B(n_868),
.Y(n_12288)
);

NOR2xp33_ASAP7_75t_L g12289 ( 
.A(n_11613),
.B(n_868),
.Y(n_12289)
);

CKINVDCx5p33_ASAP7_75t_R g12290 ( 
.A(n_11197),
.Y(n_12290)
);

INVx1_ASAP7_75t_L g12291 ( 
.A(n_11034),
.Y(n_12291)
);

BUFx8_ASAP7_75t_L g12292 ( 
.A(n_11427),
.Y(n_12292)
);

NAND2xp5_ASAP7_75t_L g12293 ( 
.A(n_11627),
.B(n_869),
.Y(n_12293)
);

NAND2xp5_ASAP7_75t_SL g12294 ( 
.A(n_11268),
.B(n_869),
.Y(n_12294)
);

NAND2xp5_ASAP7_75t_SL g12295 ( 
.A(n_11251),
.B(n_870),
.Y(n_12295)
);

AOI21x1_ASAP7_75t_L g12296 ( 
.A1(n_11271),
.A2(n_870),
.B(n_871),
.Y(n_12296)
);

BUFx6f_ASAP7_75t_L g12297 ( 
.A(n_11548),
.Y(n_12297)
);

AOI21xp5_ASAP7_75t_L g12298 ( 
.A1(n_11266),
.A2(n_871),
.B(n_872),
.Y(n_12298)
);

INVx1_ASAP7_75t_L g12299 ( 
.A(n_11040),
.Y(n_12299)
);

NAND2xp5_ASAP7_75t_SL g12300 ( 
.A(n_11085),
.B(n_872),
.Y(n_12300)
);

INVx2_ASAP7_75t_L g12301 ( 
.A(n_11045),
.Y(n_12301)
);

AOI21xp5_ASAP7_75t_L g12302 ( 
.A1(n_11272),
.A2(n_873),
.B(n_874),
.Y(n_12302)
);

OAI21xp33_ASAP7_75t_L g12303 ( 
.A1(n_11389),
.A2(n_874),
.B(n_875),
.Y(n_12303)
);

AOI21xp5_ASAP7_75t_L g12304 ( 
.A1(n_11283),
.A2(n_876),
.B(n_877),
.Y(n_12304)
);

INVx3_ASAP7_75t_L g12305 ( 
.A(n_11646),
.Y(n_12305)
);

A2O1A1Ixp33_ASAP7_75t_L g12306 ( 
.A1(n_11525),
.A2(n_879),
.B(n_877),
.C(n_878),
.Y(n_12306)
);

OAI22xp5_ASAP7_75t_L g12307 ( 
.A1(n_11464),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.Y(n_12307)
);

INVx1_ASAP7_75t_L g12308 ( 
.A(n_11236),
.Y(n_12308)
);

AOI22xp5_ASAP7_75t_L g12309 ( 
.A1(n_11728),
.A2(n_882),
.B1(n_880),
.B2(n_881),
.Y(n_12309)
);

HB1xp67_ASAP7_75t_L g12310 ( 
.A(n_11750),
.Y(n_12310)
);

INVx3_ASAP7_75t_L g12311 ( 
.A(n_11515),
.Y(n_12311)
);

INVx1_ASAP7_75t_L g12312 ( 
.A(n_11226),
.Y(n_12312)
);

INVx1_ASAP7_75t_L g12313 ( 
.A(n_11257),
.Y(n_12313)
);

NOR2xp33_ASAP7_75t_L g12314 ( 
.A(n_11246),
.B(n_11015),
.Y(n_12314)
);

O2A1O1Ixp33_ASAP7_75t_L g12315 ( 
.A1(n_11526),
.A2(n_884),
.B(n_881),
.C(n_883),
.Y(n_12315)
);

INVx2_ASAP7_75t_L g12316 ( 
.A(n_11125),
.Y(n_12316)
);

BUFx3_ASAP7_75t_L g12317 ( 
.A(n_11552),
.Y(n_12317)
);

AOI21xp5_ASAP7_75t_L g12318 ( 
.A1(n_11289),
.A2(n_883),
.B(n_884),
.Y(n_12318)
);

BUFx2_ASAP7_75t_L g12319 ( 
.A(n_11189),
.Y(n_12319)
);

BUFx2_ASAP7_75t_L g12320 ( 
.A(n_11293),
.Y(n_12320)
);

INVx2_ASAP7_75t_L g12321 ( 
.A(n_11631),
.Y(n_12321)
);

OR2x2_ASAP7_75t_L g12322 ( 
.A(n_11022),
.B(n_885),
.Y(n_12322)
);

OAI22xp5_ASAP7_75t_L g12323 ( 
.A1(n_11081),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.Y(n_12323)
);

INVx1_ASAP7_75t_L g12324 ( 
.A(n_11257),
.Y(n_12324)
);

NAND2xp5_ASAP7_75t_L g12325 ( 
.A(n_11636),
.B(n_886),
.Y(n_12325)
);

NAND2xp5_ASAP7_75t_SL g12326 ( 
.A(n_11375),
.B(n_887),
.Y(n_12326)
);

NAND2xp5_ASAP7_75t_L g12327 ( 
.A(n_11642),
.B(n_888),
.Y(n_12327)
);

AOI21xp5_ASAP7_75t_L g12328 ( 
.A1(n_11295),
.A2(n_889),
.B(n_890),
.Y(n_12328)
);

BUFx2_ASAP7_75t_L g12329 ( 
.A(n_11453),
.Y(n_12329)
);

NOR2x1_ASAP7_75t_L g12330 ( 
.A(n_11645),
.B(n_11650),
.Y(n_12330)
);

NAND2xp5_ASAP7_75t_L g12331 ( 
.A(n_11653),
.B(n_889),
.Y(n_12331)
);

NOR2xp33_ASAP7_75t_L g12332 ( 
.A(n_11054),
.B(n_890),
.Y(n_12332)
);

O2A1O1Ixp33_ASAP7_75t_L g12333 ( 
.A1(n_11200),
.A2(n_893),
.B(n_891),
.C(n_892),
.Y(n_12333)
);

AOI21xp5_ASAP7_75t_L g12334 ( 
.A1(n_11296),
.A2(n_11307),
.B(n_11099),
.Y(n_12334)
);

NAND2xp5_ASAP7_75t_SL g12335 ( 
.A(n_11426),
.B(n_891),
.Y(n_12335)
);

A2O1A1Ixp33_ASAP7_75t_L g12336 ( 
.A1(n_11378),
.A2(n_894),
.B(n_892),
.C(n_893),
.Y(n_12336)
);

O2A1O1Ixp5_ASAP7_75t_SL g12337 ( 
.A1(n_11480),
.A2(n_897),
.B(n_895),
.C(n_896),
.Y(n_12337)
);

OAI22xp5_ASAP7_75t_L g12338 ( 
.A1(n_11481),
.A2(n_898),
.B1(n_895),
.B2(n_896),
.Y(n_12338)
);

NOR3xp33_ASAP7_75t_SL g12339 ( 
.A(n_11355),
.B(n_898),
.C(n_899),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_SL g12340 ( 
.A(n_11420),
.B(n_899),
.Y(n_12340)
);

INVx1_ASAP7_75t_L g12341 ( 
.A(n_11654),
.Y(n_12341)
);

NAND2xp5_ASAP7_75t_L g12342 ( 
.A(n_11663),
.B(n_11666),
.Y(n_12342)
);

OAI22xp5_ASAP7_75t_L g12343 ( 
.A1(n_11547),
.A2(n_902),
.B1(n_900),
.B2(n_901),
.Y(n_12343)
);

O2A1O1Ixp33_ASAP7_75t_L g12344 ( 
.A1(n_11506),
.A2(n_903),
.B(n_900),
.C(n_901),
.Y(n_12344)
);

BUFx6f_ASAP7_75t_L g12345 ( 
.A(n_11551),
.Y(n_12345)
);

NAND2xp5_ASAP7_75t_SL g12346 ( 
.A(n_11470),
.B(n_903),
.Y(n_12346)
);

BUFx6f_ASAP7_75t_L g12347 ( 
.A(n_11428),
.Y(n_12347)
);

NAND2xp5_ASAP7_75t_L g12348 ( 
.A(n_11670),
.B(n_904),
.Y(n_12348)
);

INVx1_ASAP7_75t_L g12349 ( 
.A(n_11673),
.Y(n_12349)
);

AND2x2_ASAP7_75t_L g12350 ( 
.A(n_11477),
.B(n_904),
.Y(n_12350)
);

NOR2xp33_ASAP7_75t_L g12351 ( 
.A(n_11370),
.B(n_905),
.Y(n_12351)
);

NAND2xp5_ASAP7_75t_L g12352 ( 
.A(n_11676),
.B(n_905),
.Y(n_12352)
);

OAI22xp5_ASAP7_75t_SL g12353 ( 
.A1(n_11543),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_12353)
);

INVx5_ASAP7_75t_L g12354 ( 
.A(n_11478),
.Y(n_12354)
);

AOI21x1_ASAP7_75t_L g12355 ( 
.A1(n_11468),
.A2(n_906),
.B(n_907),
.Y(n_12355)
);

NOR2xp33_ASAP7_75t_R g12356 ( 
.A(n_11520),
.B(n_908),
.Y(n_12356)
);

NAND2xp33_ASAP7_75t_SL g12357 ( 
.A(n_11692),
.B(n_909),
.Y(n_12357)
);

INVx2_ASAP7_75t_L g12358 ( 
.A(n_11693),
.Y(n_12358)
);

NAND2xp5_ASAP7_75t_L g12359 ( 
.A(n_11697),
.B(n_909),
.Y(n_12359)
);

INVx2_ASAP7_75t_L g12360 ( 
.A(n_11698),
.Y(n_12360)
);

AOI21xp5_ASAP7_75t_L g12361 ( 
.A1(n_11048),
.A2(n_910),
.B(n_911),
.Y(n_12361)
);

NOR2xp33_ASAP7_75t_L g12362 ( 
.A(n_11700),
.B(n_910),
.Y(n_12362)
);

AOI22xp5_ASAP7_75t_L g12363 ( 
.A1(n_11407),
.A2(n_913),
.B1(n_911),
.B2(n_912),
.Y(n_12363)
);

OAI22xp5_ASAP7_75t_SL g12364 ( 
.A1(n_11501),
.A2(n_916),
.B1(n_914),
.B2(n_915),
.Y(n_12364)
);

INVx1_ASAP7_75t_L g12365 ( 
.A(n_11701),
.Y(n_12365)
);

NOR2xp33_ASAP7_75t_L g12366 ( 
.A(n_11717),
.B(n_914),
.Y(n_12366)
);

INVx1_ASAP7_75t_L g12367 ( 
.A(n_11722),
.Y(n_12367)
);

OAI22xp5_ASAP7_75t_L g12368 ( 
.A1(n_11528),
.A2(n_919),
.B1(n_917),
.B2(n_918),
.Y(n_12368)
);

BUFx6f_ASAP7_75t_L g12369 ( 
.A(n_11535),
.Y(n_12369)
);

BUFx2_ASAP7_75t_L g12370 ( 
.A(n_11458),
.Y(n_12370)
);

AOI21x1_ASAP7_75t_L g12371 ( 
.A1(n_11421),
.A2(n_917),
.B(n_918),
.Y(n_12371)
);

AOI21xp5_ASAP7_75t_L g12372 ( 
.A1(n_11199),
.A2(n_919),
.B(n_920),
.Y(n_12372)
);

O2A1O1Ixp33_ASAP7_75t_L g12373 ( 
.A1(n_11540),
.A2(n_922),
.B(n_920),
.C(n_921),
.Y(n_12373)
);

AOI21xp5_ASAP7_75t_L g12374 ( 
.A1(n_11204),
.A2(n_921),
.B(n_922),
.Y(n_12374)
);

NAND2xp5_ASAP7_75t_L g12375 ( 
.A(n_11729),
.B(n_923),
.Y(n_12375)
);

NAND2xp5_ASAP7_75t_SL g12376 ( 
.A(n_11731),
.B(n_923),
.Y(n_12376)
);

BUFx2_ASAP7_75t_L g12377 ( 
.A(n_11249),
.Y(n_12377)
);

INVx4_ASAP7_75t_L g12378 ( 
.A(n_11337),
.Y(n_12378)
);

BUFx6f_ASAP7_75t_L g12379 ( 
.A(n_11417),
.Y(n_12379)
);

A2O1A1Ixp33_ASAP7_75t_L g12380 ( 
.A1(n_11497),
.A2(n_926),
.B(n_924),
.C(n_925),
.Y(n_12380)
);

NAND2xp5_ASAP7_75t_L g12381 ( 
.A(n_11739),
.B(n_924),
.Y(n_12381)
);

O2A1O1Ixp33_ASAP7_75t_L g12382 ( 
.A1(n_11209),
.A2(n_928),
.B(n_925),
.C(n_927),
.Y(n_12382)
);

NAND2xp5_ASAP7_75t_L g12383 ( 
.A(n_11404),
.B(n_927),
.Y(n_12383)
);

BUFx6f_ASAP7_75t_L g12384 ( 
.A(n_11276),
.Y(n_12384)
);

NAND2xp5_ASAP7_75t_L g12385 ( 
.A(n_11413),
.B(n_929),
.Y(n_12385)
);

AOI22xp33_ASAP7_75t_L g12386 ( 
.A1(n_11371),
.A2(n_931),
.B1(n_929),
.B2(n_930),
.Y(n_12386)
);

INVx1_ASAP7_75t_L g12387 ( 
.A(n_11242),
.Y(n_12387)
);

AOI21xp5_ASAP7_75t_L g12388 ( 
.A1(n_11101),
.A2(n_930),
.B(n_931),
.Y(n_12388)
);

NAND2xp5_ASAP7_75t_L g12389 ( 
.A(n_11097),
.B(n_932),
.Y(n_12389)
);

NAND2xp5_ASAP7_75t_SL g12390 ( 
.A(n_11433),
.B(n_932),
.Y(n_12390)
);

AOI21x1_ASAP7_75t_SL g12391 ( 
.A1(n_11108),
.A2(n_933),
.B(n_934),
.Y(n_12391)
);

INVxp67_ASAP7_75t_L g12392 ( 
.A(n_11245),
.Y(n_12392)
);

NOR3xp33_ASAP7_75t_L g12393 ( 
.A(n_11020),
.B(n_933),
.C(n_934),
.Y(n_12393)
);

NOR2xp33_ASAP7_75t_L g12394 ( 
.A(n_11374),
.B(n_935),
.Y(n_12394)
);

NAND2xp5_ASAP7_75t_L g12395 ( 
.A(n_11105),
.B(n_936),
.Y(n_12395)
);

NAND2xp5_ASAP7_75t_L g12396 ( 
.A(n_11114),
.B(n_936),
.Y(n_12396)
);

OAI22xp5_ASAP7_75t_L g12397 ( 
.A1(n_11158),
.A2(n_939),
.B1(n_937),
.B2(n_938),
.Y(n_12397)
);

NAND2xp5_ASAP7_75t_L g12398 ( 
.A(n_11117),
.B(n_937),
.Y(n_12398)
);

INVx2_ASAP7_75t_L g12399 ( 
.A(n_11519),
.Y(n_12399)
);

OR2x2_ASAP7_75t_L g12400 ( 
.A(n_11419),
.B(n_939),
.Y(n_12400)
);

NAND2xp5_ASAP7_75t_L g12401 ( 
.A(n_11229),
.B(n_940),
.Y(n_12401)
);

AOI21xp5_ASAP7_75t_L g12402 ( 
.A1(n_11259),
.A2(n_940),
.B(n_941),
.Y(n_12402)
);

AOI21x1_ASAP7_75t_L g12403 ( 
.A1(n_11536),
.A2(n_11625),
.B(n_11573),
.Y(n_12403)
);

AOI21x1_ASAP7_75t_L g12404 ( 
.A1(n_11634),
.A2(n_941),
.B(n_942),
.Y(n_12404)
);

OAI22xp5_ASAP7_75t_L g12405 ( 
.A1(n_11749),
.A2(n_945),
.B1(n_943),
.B2(n_944),
.Y(n_12405)
);

O2A1O1Ixp33_ASAP7_75t_L g12406 ( 
.A1(n_11274),
.A2(n_946),
.B(n_943),
.C(n_945),
.Y(n_12406)
);

NAND2xp5_ASAP7_75t_SL g12407 ( 
.A(n_11437),
.B(n_946),
.Y(n_12407)
);

NAND2xp5_ASAP7_75t_L g12408 ( 
.A(n_11401),
.B(n_947),
.Y(n_12408)
);

AOI21xp5_ASAP7_75t_L g12409 ( 
.A1(n_11063),
.A2(n_947),
.B(n_948),
.Y(n_12409)
);

BUFx6f_ASAP7_75t_L g12410 ( 
.A(n_11247),
.Y(n_12410)
);

A2O1A1Ixp33_ASAP7_75t_SL g12411 ( 
.A1(n_11545),
.A2(n_950),
.B(n_948),
.C(n_949),
.Y(n_12411)
);

BUFx3_ASAP7_75t_L g12412 ( 
.A(n_11150),
.Y(n_12412)
);

AOI21xp5_ASAP7_75t_L g12413 ( 
.A1(n_11065),
.A2(n_949),
.B(n_951),
.Y(n_12413)
);

NAND2xp5_ASAP7_75t_L g12414 ( 
.A(n_11398),
.B(n_11387),
.Y(n_12414)
);

NAND2xp5_ASAP7_75t_L g12415 ( 
.A(n_11435),
.B(n_951),
.Y(n_12415)
);

OAI22x1_ASAP7_75t_L g12416 ( 
.A1(n_11064),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.Y(n_12416)
);

NOR3xp33_ASAP7_75t_SL g12417 ( 
.A(n_11002),
.B(n_953),
.C(n_954),
.Y(n_12417)
);

NOR2xp33_ASAP7_75t_L g12418 ( 
.A(n_11483),
.B(n_955),
.Y(n_12418)
);

A2O1A1Ixp33_ASAP7_75t_L g12419 ( 
.A1(n_11550),
.A2(n_957),
.B(n_955),
.C(n_956),
.Y(n_12419)
);

O2A1O1Ixp33_ASAP7_75t_L g12420 ( 
.A1(n_11076),
.A2(n_959),
.B(n_957),
.C(n_958),
.Y(n_12420)
);

INVx2_ASAP7_75t_L g12421 ( 
.A(n_11390),
.Y(n_12421)
);

O2A1O1Ixp33_ASAP7_75t_L g12422 ( 
.A1(n_11248),
.A2(n_960),
.B(n_958),
.C(n_959),
.Y(n_12422)
);

INVx5_ASAP7_75t_L g12423 ( 
.A(n_11086),
.Y(n_12423)
);

O2A1O1Ixp33_ASAP7_75t_L g12424 ( 
.A1(n_11161),
.A2(n_962),
.B(n_960),
.C(n_961),
.Y(n_12424)
);

NAND2xp5_ASAP7_75t_L g12425 ( 
.A(n_11469),
.B(n_961),
.Y(n_12425)
);

OAI22xp33_ASAP7_75t_L g12426 ( 
.A1(n_11357),
.A2(n_964),
.B1(n_962),
.B2(n_963),
.Y(n_12426)
);

OAI22xp5_ASAP7_75t_L g12427 ( 
.A1(n_11521),
.A2(n_965),
.B1(n_963),
.B2(n_964),
.Y(n_12427)
);

INVxp67_ASAP7_75t_L g12428 ( 
.A(n_11157),
.Y(n_12428)
);

NAND2xp5_ASAP7_75t_L g12429 ( 
.A(n_11472),
.B(n_965),
.Y(n_12429)
);

HB1xp67_ASAP7_75t_L g12430 ( 
.A(n_11537),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_11479),
.Y(n_12431)
);

AOI21xp5_ASAP7_75t_L g12432 ( 
.A1(n_11068),
.A2(n_966),
.B(n_967),
.Y(n_12432)
);

CKINVDCx5p33_ASAP7_75t_R g12433 ( 
.A(n_11493),
.Y(n_12433)
);

BUFx6f_ASAP7_75t_L g12434 ( 
.A(n_11486),
.Y(n_12434)
);

AOI21xp5_ASAP7_75t_L g12435 ( 
.A1(n_11082),
.A2(n_966),
.B(n_967),
.Y(n_12435)
);

OAI22xp5_ASAP7_75t_L g12436 ( 
.A1(n_11490),
.A2(n_970),
.B1(n_968),
.B2(n_969),
.Y(n_12436)
);

NAND2xp5_ASAP7_75t_L g12437 ( 
.A(n_11496),
.B(n_968),
.Y(n_12437)
);

INVx2_ASAP7_75t_L g12438 ( 
.A(n_11291),
.Y(n_12438)
);

BUFx2_ASAP7_75t_L g12439 ( 
.A(n_11502),
.Y(n_12439)
);

AOI21xp5_ASAP7_75t_L g12440 ( 
.A1(n_11084),
.A2(n_969),
.B(n_971),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_11503),
.Y(n_12441)
);

OAI21xp5_ASAP7_75t_L g12442 ( 
.A1(n_11361),
.A2(n_971),
.B(n_972),
.Y(n_12442)
);

INVx1_ASAP7_75t_L g12443 ( 
.A(n_11510),
.Y(n_12443)
);

INVx1_ASAP7_75t_L g12444 ( 
.A(n_11511),
.Y(n_12444)
);

INVx2_ASAP7_75t_L g12445 ( 
.A(n_11318),
.Y(n_12445)
);

OAI21xp33_ASAP7_75t_L g12446 ( 
.A1(n_11512),
.A2(n_974),
.B(n_975),
.Y(n_12446)
);

OAI22xp5_ASAP7_75t_L g12447 ( 
.A1(n_11522),
.A2(n_976),
.B1(n_974),
.B2(n_975),
.Y(n_12447)
);

BUFx6f_ASAP7_75t_L g12448 ( 
.A(n_11524),
.Y(n_12448)
);

CKINVDCx5p33_ASAP7_75t_R g12449 ( 
.A(n_11532),
.Y(n_12449)
);

AOI22xp5_ASAP7_75t_L g12450 ( 
.A1(n_11332),
.A2(n_979),
.B1(n_976),
.B2(n_978),
.Y(n_12450)
);

INVx1_ASAP7_75t_SL g12451 ( 
.A(n_11538),
.Y(n_12451)
);

BUFx2_ASAP7_75t_L g12452 ( 
.A(n_11542),
.Y(n_12452)
);

AND2x2_ASAP7_75t_SL g12453 ( 
.A(n_11544),
.B(n_978),
.Y(n_12453)
);

AND2x4_ASAP7_75t_L g12454 ( 
.A(n_11349),
.B(n_979),
.Y(n_12454)
);

HB1xp67_ASAP7_75t_L g12455 ( 
.A(n_11363),
.Y(n_12455)
);

OR2x2_ASAP7_75t_L g12456 ( 
.A(n_11365),
.B(n_980),
.Y(n_12456)
);

NAND2xp5_ASAP7_75t_L g12457 ( 
.A(n_11396),
.B(n_11397),
.Y(n_12457)
);

NAND2xp5_ASAP7_75t_SL g12458 ( 
.A(n_11444),
.B(n_981),
.Y(n_12458)
);

NOR2xp33_ASAP7_75t_L g12459 ( 
.A(n_11372),
.B(n_981),
.Y(n_12459)
);

INVx1_ASAP7_75t_L g12460 ( 
.A(n_11392),
.Y(n_12460)
);

NOR2xp67_ASAP7_75t_L g12461 ( 
.A(n_11342),
.B(n_982),
.Y(n_12461)
);

AND2x4_ASAP7_75t_L g12462 ( 
.A(n_11553),
.B(n_982),
.Y(n_12462)
);

AOI21xp5_ASAP7_75t_L g12463 ( 
.A1(n_11087),
.A2(n_983),
.B(n_984),
.Y(n_12463)
);

A2O1A1Ixp33_ASAP7_75t_L g12464 ( 
.A1(n_11499),
.A2(n_985),
.B(n_983),
.C(n_984),
.Y(n_12464)
);

OAI22xp5_ASAP7_75t_L g12465 ( 
.A1(n_11516),
.A2(n_987),
.B1(n_985),
.B2(n_986),
.Y(n_12465)
);

INVx1_ASAP7_75t_SL g12466 ( 
.A(n_11457),
.Y(n_12466)
);

A2O1A1Ixp33_ASAP7_75t_SL g12467 ( 
.A1(n_11523),
.A2(n_988),
.B(n_986),
.C(n_987),
.Y(n_12467)
);

INVx2_ASAP7_75t_L g12468 ( 
.A(n_11312),
.Y(n_12468)
);

OAI22xp5_ASAP7_75t_L g12469 ( 
.A1(n_11530),
.A2(n_990),
.B1(n_988),
.B2(n_989),
.Y(n_12469)
);

AOI21xp5_ASAP7_75t_L g12470 ( 
.A1(n_11364),
.A2(n_989),
.B(n_990),
.Y(n_12470)
);

AND2x4_ASAP7_75t_L g12471 ( 
.A(n_11362),
.B(n_991),
.Y(n_12471)
);

INVx1_ASAP7_75t_L g12472 ( 
.A(n_11329),
.Y(n_12472)
);

AOI21xp5_ASAP7_75t_L g12473 ( 
.A1(n_11213),
.A2(n_991),
.B(n_992),
.Y(n_12473)
);

NAND2xp5_ASAP7_75t_L g12474 ( 
.A(n_11533),
.B(n_992),
.Y(n_12474)
);

AOI21xp5_ASAP7_75t_L g12475 ( 
.A1(n_11219),
.A2(n_11230),
.B(n_11181),
.Y(n_12475)
);

NAND2xp5_ASAP7_75t_L g12476 ( 
.A(n_11460),
.B(n_993),
.Y(n_12476)
);

OAI22x1_ASAP7_75t_L g12477 ( 
.A1(n_11474),
.A2(n_995),
.B1(n_993),
.B2(n_994),
.Y(n_12477)
);

OR2x2_ASAP7_75t_L g12478 ( 
.A(n_11484),
.B(n_994),
.Y(n_12478)
);

INVx1_ASAP7_75t_L g12479 ( 
.A(n_11330),
.Y(n_12479)
);

NAND2xp5_ASAP7_75t_L g12480 ( 
.A(n_11494),
.B(n_995),
.Y(n_12480)
);

O2A1O1Ixp33_ASAP7_75t_L g12481 ( 
.A1(n_11011),
.A2(n_998),
.B(n_996),
.C(n_997),
.Y(n_12481)
);

BUFx6f_ASAP7_75t_L g12482 ( 
.A(n_11422),
.Y(n_12482)
);

OAI22xp5_ASAP7_75t_L g12483 ( 
.A1(n_11386),
.A2(n_998),
.B1(n_996),
.B2(n_997),
.Y(n_12483)
);

AOI21xp5_ASAP7_75t_L g12484 ( 
.A1(n_11155),
.A2(n_999),
.B(n_1000),
.Y(n_12484)
);

INVx2_ASAP7_75t_L g12485 ( 
.A(n_11106),
.Y(n_12485)
);

INVx3_ASAP7_75t_L g12486 ( 
.A(n_11409),
.Y(n_12486)
);

OAI21xp33_ASAP7_75t_SL g12487 ( 
.A1(n_11379),
.A2(n_999),
.B(n_1000),
.Y(n_12487)
);

A2O1A1Ixp33_ASAP7_75t_L g12488 ( 
.A1(n_11163),
.A2(n_1003),
.B(n_1001),
.C(n_1002),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_11111),
.Y(n_12489)
);

NAND2xp5_ASAP7_75t_L g12490 ( 
.A(n_11410),
.B(n_1001),
.Y(n_12490)
);

INVx4_ASAP7_75t_L g12491 ( 
.A(n_11241),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_11127),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_11133),
.Y(n_12493)
);

HB1xp67_ASAP7_75t_L g12494 ( 
.A(n_11135),
.Y(n_12494)
);

AOI22xp33_ASAP7_75t_L g12495 ( 
.A1(n_11518),
.A2(n_1004),
.B1(n_1002),
.B2(n_1003),
.Y(n_12495)
);

NAND2xp5_ASAP7_75t_L g12496 ( 
.A(n_11383),
.B(n_1005),
.Y(n_12496)
);

INVx2_ASAP7_75t_L g12497 ( 
.A(n_11137),
.Y(n_12497)
);

O2A1O1Ixp33_ASAP7_75t_L g12498 ( 
.A1(n_11138),
.A2(n_1008),
.B(n_1006),
.C(n_1007),
.Y(n_12498)
);

O2A1O1Ixp5_ASAP7_75t_L g12499 ( 
.A1(n_11098),
.A2(n_1008),
.B(n_1006),
.C(n_1007),
.Y(n_12499)
);

NOR3xp33_ASAP7_75t_SL g12500 ( 
.A(n_11142),
.B(n_1009),
.C(n_1010),
.Y(n_12500)
);

NAND2xp5_ASAP7_75t_SL g12501 ( 
.A(n_11060),
.B(n_1010),
.Y(n_12501)
);

O2A1O1Ixp33_ASAP7_75t_L g12502 ( 
.A1(n_11136),
.A2(n_1013),
.B(n_1011),
.C(n_1012),
.Y(n_12502)
);

INVx5_ASAP7_75t_L g12503 ( 
.A(n_11294),
.Y(n_12503)
);

NAND2xp5_ASAP7_75t_L g12504 ( 
.A(n_11091),
.B(n_1012),
.Y(n_12504)
);

AO21x1_ASAP7_75t_L g12505 ( 
.A1(n_11619),
.A2(n_1013),
.B(n_1014),
.Y(n_12505)
);

AOI21xp5_ASAP7_75t_L g12506 ( 
.A1(n_11619),
.A2(n_1014),
.B(n_1015),
.Y(n_12506)
);

NOR2xp33_ASAP7_75t_L g12507 ( 
.A(n_10971),
.B(n_1015),
.Y(n_12507)
);

NOR2xp33_ASAP7_75t_L g12508 ( 
.A(n_10971),
.B(n_1016),
.Y(n_12508)
);

AOI21xp5_ASAP7_75t_L g12509 ( 
.A1(n_11619),
.A2(n_1017),
.B(n_1018),
.Y(n_12509)
);

NAND2xp5_ASAP7_75t_SL g12510 ( 
.A(n_11060),
.B(n_1018),
.Y(n_12510)
);

NOR2x1_ASAP7_75t_R g12511 ( 
.A(n_11218),
.B(n_1019),
.Y(n_12511)
);

NAND2xp5_ASAP7_75t_SL g12512 ( 
.A(n_11060),
.B(n_1019),
.Y(n_12512)
);

AND2x2_ASAP7_75t_L g12513 ( 
.A(n_11487),
.B(n_1020),
.Y(n_12513)
);

INVx5_ASAP7_75t_L g12514 ( 
.A(n_11294),
.Y(n_12514)
);

A2O1A1Ixp33_ASAP7_75t_L g12515 ( 
.A1(n_10986),
.A2(n_1023),
.B(n_1021),
.C(n_1022),
.Y(n_12515)
);

O2A1O1Ixp33_ASAP7_75t_L g12516 ( 
.A1(n_11136),
.A2(n_1024),
.B(n_1021),
.C(n_1023),
.Y(n_12516)
);

BUFx8_ASAP7_75t_L g12517 ( 
.A(n_11012),
.Y(n_12517)
);

NAND2xp5_ASAP7_75t_SL g12518 ( 
.A(n_11060),
.B(n_1024),
.Y(n_12518)
);

INVx2_ASAP7_75t_L g12519 ( 
.A(n_11267),
.Y(n_12519)
);

INVx2_ASAP7_75t_L g12520 ( 
.A(n_11267),
.Y(n_12520)
);

AND2x4_ASAP7_75t_L g12521 ( 
.A(n_11556),
.B(n_1025),
.Y(n_12521)
);

OAI22xp5_ASAP7_75t_L g12522 ( 
.A1(n_11309),
.A2(n_1027),
.B1(n_1025),
.B2(n_1026),
.Y(n_12522)
);

NAND2xp5_ASAP7_75t_L g12523 ( 
.A(n_11091),
.B(n_1026),
.Y(n_12523)
);

NAND2xp5_ASAP7_75t_L g12524 ( 
.A(n_11091),
.B(n_1027),
.Y(n_12524)
);

OAI22xp5_ASAP7_75t_L g12525 ( 
.A1(n_11309),
.A2(n_1030),
.B1(n_1028),
.B2(n_1029),
.Y(n_12525)
);

AOI21xp5_ASAP7_75t_L g12526 ( 
.A1(n_11619),
.A2(n_1029),
.B(n_1030),
.Y(n_12526)
);

NOR2xp33_ASAP7_75t_L g12527 ( 
.A(n_10971),
.B(n_1031),
.Y(n_12527)
);

INVx5_ASAP7_75t_L g12528 ( 
.A(n_11294),
.Y(n_12528)
);

A2O1A1Ixp33_ASAP7_75t_L g12529 ( 
.A1(n_10986),
.A2(n_1033),
.B(n_1031),
.C(n_1032),
.Y(n_12529)
);

BUFx6f_ASAP7_75t_L g12530 ( 
.A(n_11012),
.Y(n_12530)
);

BUFx4f_ASAP7_75t_SL g12531 ( 
.A(n_11218),
.Y(n_12531)
);

INVx2_ASAP7_75t_L g12532 ( 
.A(n_11267),
.Y(n_12532)
);

AND2x4_ASAP7_75t_L g12533 ( 
.A(n_11556),
.B(n_1032),
.Y(n_12533)
);

AO21x1_ASAP7_75t_L g12534 ( 
.A1(n_11619),
.A2(n_1033),
.B(n_1034),
.Y(n_12534)
);

AOI21xp5_ASAP7_75t_L g12535 ( 
.A1(n_11619),
.A2(n_1034),
.B(n_1035),
.Y(n_12535)
);

NAND2xp5_ASAP7_75t_SL g12536 ( 
.A(n_11060),
.B(n_1035),
.Y(n_12536)
);

A2O1A1Ixp33_ASAP7_75t_L g12537 ( 
.A1(n_10986),
.A2(n_1038),
.B(n_1036),
.C(n_1037),
.Y(n_12537)
);

AOI21xp5_ASAP7_75t_L g12538 ( 
.A1(n_11619),
.A2(n_1036),
.B(n_1038),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_11267),
.Y(n_12539)
);

NOR2xp33_ASAP7_75t_L g12540 ( 
.A(n_10971),
.B(n_1039),
.Y(n_12540)
);

AND2x2_ASAP7_75t_L g12541 ( 
.A(n_11487),
.B(n_1039),
.Y(n_12541)
);

AOI21xp5_ASAP7_75t_L g12542 ( 
.A1(n_11619),
.A2(n_1040),
.B(n_1041),
.Y(n_12542)
);

NAND2xp5_ASAP7_75t_SL g12543 ( 
.A(n_11060),
.B(n_1041),
.Y(n_12543)
);

INVx2_ASAP7_75t_L g12544 ( 
.A(n_11267),
.Y(n_12544)
);

A2O1A1Ixp33_ASAP7_75t_SL g12545 ( 
.A1(n_11561),
.A2(n_1044),
.B(n_1042),
.C(n_1043),
.Y(n_12545)
);

O2A1O1Ixp33_ASAP7_75t_SL g12546 ( 
.A1(n_11136),
.A2(n_1045),
.B(n_1042),
.C(n_1044),
.Y(n_12546)
);

CKINVDCx5p33_ASAP7_75t_R g12547 ( 
.A(n_11590),
.Y(n_12547)
);

OR2x6_ASAP7_75t_L g12548 ( 
.A(n_11005),
.B(n_1045),
.Y(n_12548)
);

OAI22xp5_ASAP7_75t_L g12549 ( 
.A1(n_11309),
.A2(n_1049),
.B1(n_1046),
.B2(n_1047),
.Y(n_12549)
);

AOI21xp5_ASAP7_75t_L g12550 ( 
.A1(n_11619),
.A2(n_1046),
.B(n_1047),
.Y(n_12550)
);

INVx1_ASAP7_75t_SL g12551 ( 
.A(n_11679),
.Y(n_12551)
);

BUFx2_ASAP7_75t_L g12552 ( 
.A(n_11178),
.Y(n_12552)
);

A2O1A1Ixp33_ASAP7_75t_L g12553 ( 
.A1(n_10986),
.A2(n_1052),
.B(n_1050),
.C(n_1051),
.Y(n_12553)
);

AND2x2_ASAP7_75t_L g12554 ( 
.A(n_11487),
.B(n_1050),
.Y(n_12554)
);

NOR3xp33_ASAP7_75t_SL g12555 ( 
.A(n_11366),
.B(n_1051),
.C(n_1052),
.Y(n_12555)
);

OAI22xp5_ASAP7_75t_L g12556 ( 
.A1(n_11309),
.A2(n_1055),
.B1(n_1053),
.B2(n_1054),
.Y(n_12556)
);

O2A1O1Ixp33_ASAP7_75t_SL g12557 ( 
.A1(n_11136),
.A2(n_1056),
.B(n_1053),
.C(n_1055),
.Y(n_12557)
);

INVx1_ASAP7_75t_L g12558 ( 
.A(n_10996),
.Y(n_12558)
);

NAND2xp5_ASAP7_75t_L g12559 ( 
.A(n_11091),
.B(n_1056),
.Y(n_12559)
);

NOR2xp33_ASAP7_75t_L g12560 ( 
.A(n_10971),
.B(n_1057),
.Y(n_12560)
);

INVxp67_ASAP7_75t_L g12561 ( 
.A(n_11315),
.Y(n_12561)
);

CKINVDCx5p33_ASAP7_75t_R g12562 ( 
.A(n_11590),
.Y(n_12562)
);

AOI22xp33_ASAP7_75t_L g12563 ( 
.A1(n_11619),
.A2(n_1059),
.B1(n_1057),
.B2(n_1058),
.Y(n_12563)
);

AOI21xp5_ASAP7_75t_L g12564 ( 
.A1(n_11619),
.A2(n_1058),
.B(n_1060),
.Y(n_12564)
);

INVx1_ASAP7_75t_L g12565 ( 
.A(n_10996),
.Y(n_12565)
);

AOI21x1_ASAP7_75t_L g12566 ( 
.A1(n_11005),
.A2(n_1060),
.B(n_1062),
.Y(n_12566)
);

NAND2xp5_ASAP7_75t_L g12567 ( 
.A(n_11091),
.B(n_1062),
.Y(n_12567)
);

O2A1O1Ixp33_ASAP7_75t_SL g12568 ( 
.A1(n_11136),
.A2(n_1065),
.B(n_1063),
.C(n_1064),
.Y(n_12568)
);

INVx1_ASAP7_75t_L g12569 ( 
.A(n_10996),
.Y(n_12569)
);

INVxp67_ASAP7_75t_L g12570 ( 
.A(n_11315),
.Y(n_12570)
);

INVx3_ASAP7_75t_L g12571 ( 
.A(n_11316),
.Y(n_12571)
);

OAI22xp5_ASAP7_75t_L g12572 ( 
.A1(n_11309),
.A2(n_1066),
.B1(n_1063),
.B2(n_1065),
.Y(n_12572)
);

A2O1A1Ixp33_ASAP7_75t_L g12573 ( 
.A1(n_10986),
.A2(n_1068),
.B(n_1066),
.C(n_1067),
.Y(n_12573)
);

BUFx2_ASAP7_75t_L g12574 ( 
.A(n_11178),
.Y(n_12574)
);

AOI21xp5_ASAP7_75t_L g12575 ( 
.A1(n_11619),
.A2(n_1067),
.B(n_1068),
.Y(n_12575)
);

BUFx2_ASAP7_75t_L g12576 ( 
.A(n_11178),
.Y(n_12576)
);

NAND2xp5_ASAP7_75t_SL g12577 ( 
.A(n_11060),
.B(n_1069),
.Y(n_12577)
);

AOI21xp5_ASAP7_75t_L g12578 ( 
.A1(n_11619),
.A2(n_1069),
.B(n_1070),
.Y(n_12578)
);

AOI21xp5_ASAP7_75t_L g12579 ( 
.A1(n_11619),
.A2(n_1070),
.B(n_1071),
.Y(n_12579)
);

OAI21xp33_ASAP7_75t_L g12580 ( 
.A1(n_10982),
.A2(n_1071),
.B(n_1072),
.Y(n_12580)
);

INVx2_ASAP7_75t_L g12581 ( 
.A(n_11267),
.Y(n_12581)
);

NAND2xp5_ASAP7_75t_L g12582 ( 
.A(n_11091),
.B(n_1072),
.Y(n_12582)
);

INVx1_ASAP7_75t_L g12583 ( 
.A(n_10996),
.Y(n_12583)
);

NOR2xp33_ASAP7_75t_SL g12584 ( 
.A(n_10981),
.B(n_1073),
.Y(n_12584)
);

NOR2xp33_ASAP7_75t_R g12585 ( 
.A(n_11590),
.B(n_1073),
.Y(n_12585)
);

A2O1A1Ixp33_ASAP7_75t_L g12586 ( 
.A1(n_10986),
.A2(n_1076),
.B(n_1074),
.C(n_1075),
.Y(n_12586)
);

NAND2xp5_ASAP7_75t_L g12587 ( 
.A(n_11091),
.B(n_1074),
.Y(n_12587)
);

INVx1_ASAP7_75t_L g12588 ( 
.A(n_10996),
.Y(n_12588)
);

INVx2_ASAP7_75t_L g12589 ( 
.A(n_11267),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_10996),
.Y(n_12590)
);

NAND3xp33_ASAP7_75t_SL g12591 ( 
.A(n_10982),
.B(n_1075),
.C(n_1076),
.Y(n_12591)
);

NAND2xp5_ASAP7_75t_L g12592 ( 
.A(n_11091),
.B(n_1077),
.Y(n_12592)
);

NAND2xp5_ASAP7_75t_SL g12593 ( 
.A(n_11060),
.B(n_1077),
.Y(n_12593)
);

INVx2_ASAP7_75t_L g12594 ( 
.A(n_11267),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_11267),
.Y(n_12595)
);

OAI22xp5_ASAP7_75t_L g12596 ( 
.A1(n_11309),
.A2(n_1080),
.B1(n_1078),
.B2(n_1079),
.Y(n_12596)
);

NAND2xp5_ASAP7_75t_L g12597 ( 
.A(n_11091),
.B(n_1079),
.Y(n_12597)
);

NAND2xp5_ASAP7_75t_L g12598 ( 
.A(n_11091),
.B(n_1081),
.Y(n_12598)
);

INVx6_ASAP7_75t_L g12599 ( 
.A(n_11012),
.Y(n_12599)
);

NAND2xp5_ASAP7_75t_SL g12600 ( 
.A(n_11060),
.B(n_1081),
.Y(n_12600)
);

NOR2xp33_ASAP7_75t_L g12601 ( 
.A(n_10971),
.B(n_1082),
.Y(n_12601)
);

AOI22xp33_ASAP7_75t_SL g12602 ( 
.A1(n_11619),
.A2(n_1084),
.B1(n_1082),
.B2(n_1083),
.Y(n_12602)
);

AOI21xp5_ASAP7_75t_L g12603 ( 
.A1(n_11619),
.A2(n_1083),
.B(n_1084),
.Y(n_12603)
);

INVx2_ASAP7_75t_L g12604 ( 
.A(n_11267),
.Y(n_12604)
);

AOI21xp5_ASAP7_75t_L g12605 ( 
.A1(n_11619),
.A2(n_1085),
.B(n_1086),
.Y(n_12605)
);

NAND2xp5_ASAP7_75t_SL g12606 ( 
.A(n_11060),
.B(n_1085),
.Y(n_12606)
);

O2A1O1Ixp5_ASAP7_75t_L g12607 ( 
.A1(n_10979),
.A2(n_1088),
.B(n_1086),
.C(n_1087),
.Y(n_12607)
);

AOI22xp33_ASAP7_75t_L g12608 ( 
.A1(n_11619),
.A2(n_1089),
.B1(n_1087),
.B2(n_1088),
.Y(n_12608)
);

NAND2xp5_ASAP7_75t_L g12609 ( 
.A(n_11091),
.B(n_1089),
.Y(n_12609)
);

NOR2xp33_ASAP7_75t_L g12610 ( 
.A(n_10971),
.B(n_1090),
.Y(n_12610)
);

NOR2xp33_ASAP7_75t_L g12611 ( 
.A(n_10971),
.B(n_1090),
.Y(n_12611)
);

CKINVDCx5p33_ASAP7_75t_R g12612 ( 
.A(n_11590),
.Y(n_12612)
);

NAND2xp5_ASAP7_75t_L g12613 ( 
.A(n_11091),
.B(n_1091),
.Y(n_12613)
);

A2O1A1Ixp33_ASAP7_75t_L g12614 ( 
.A1(n_10986),
.A2(n_1095),
.B(n_1091),
.C(n_1093),
.Y(n_12614)
);

NOR2xp33_ASAP7_75t_R g12615 ( 
.A(n_11590),
.B(n_1093),
.Y(n_12615)
);

NAND2xp5_ASAP7_75t_SL g12616 ( 
.A(n_11060),
.B(n_1095),
.Y(n_12616)
);

OAI21xp33_ASAP7_75t_SL g12617 ( 
.A1(n_11561),
.A2(n_1096),
.B(n_1097),
.Y(n_12617)
);

AOI21xp5_ASAP7_75t_L g12618 ( 
.A1(n_11619),
.A2(n_1096),
.B(n_1098),
.Y(n_12618)
);

OAI22xp5_ASAP7_75t_L g12619 ( 
.A1(n_11309),
.A2(n_1100),
.B1(n_1098),
.B2(n_1099),
.Y(n_12619)
);

OAI22xp5_ASAP7_75t_L g12620 ( 
.A1(n_11309),
.A2(n_1102),
.B1(n_1100),
.B2(n_1101),
.Y(n_12620)
);

INVx1_ASAP7_75t_L g12621 ( 
.A(n_10996),
.Y(n_12621)
);

INVx4_ASAP7_75t_L g12622 ( 
.A(n_11012),
.Y(n_12622)
);

NAND2xp5_ASAP7_75t_SL g12623 ( 
.A(n_11060),
.B(n_1101),
.Y(n_12623)
);

INVx2_ASAP7_75t_L g12624 ( 
.A(n_11267),
.Y(n_12624)
);

AOI21xp5_ASAP7_75t_L g12625 ( 
.A1(n_11619),
.A2(n_1102),
.B(n_1103),
.Y(n_12625)
);

NAND2xp5_ASAP7_75t_L g12626 ( 
.A(n_11091),
.B(n_1103),
.Y(n_12626)
);

AOI21xp5_ASAP7_75t_L g12627 ( 
.A1(n_11619),
.A2(n_1104),
.B(n_1105),
.Y(n_12627)
);

NOR2xp33_ASAP7_75t_L g12628 ( 
.A(n_10971),
.B(n_1104),
.Y(n_12628)
);

AOI21xp5_ASAP7_75t_L g12629 ( 
.A1(n_11619),
.A2(n_1105),
.B(n_1107),
.Y(n_12629)
);

NOR3xp33_ASAP7_75t_SL g12630 ( 
.A(n_11366),
.B(n_1107),
.C(n_1109),
.Y(n_12630)
);

INVx1_ASAP7_75t_L g12631 ( 
.A(n_10996),
.Y(n_12631)
);

AOI22xp5_ASAP7_75t_L g12632 ( 
.A1(n_11619),
.A2(n_1111),
.B1(n_1109),
.B2(n_1110),
.Y(n_12632)
);

AOI21xp5_ASAP7_75t_L g12633 ( 
.A1(n_11619),
.A2(n_1110),
.B(n_1112),
.Y(n_12633)
);

NAND2xp5_ASAP7_75t_L g12634 ( 
.A(n_11091),
.B(n_1113),
.Y(n_12634)
);

A2O1A1Ixp33_ASAP7_75t_L g12635 ( 
.A1(n_10986),
.A2(n_1115),
.B(n_1113),
.C(n_1114),
.Y(n_12635)
);

A2O1A1Ixp33_ASAP7_75t_L g12636 ( 
.A1(n_10986),
.A2(n_1116),
.B(n_1114),
.C(n_1115),
.Y(n_12636)
);

AOI22xp5_ASAP7_75t_L g12637 ( 
.A1(n_11619),
.A2(n_1118),
.B1(n_1116),
.B2(n_1117),
.Y(n_12637)
);

NAND2xp5_ASAP7_75t_L g12638 ( 
.A(n_11091),
.B(n_1117),
.Y(n_12638)
);

OAI22xp5_ASAP7_75t_L g12639 ( 
.A1(n_11309),
.A2(n_1120),
.B1(n_1118),
.B2(n_1119),
.Y(n_12639)
);

INVx2_ASAP7_75t_L g12640 ( 
.A(n_11267),
.Y(n_12640)
);

AOI21xp5_ASAP7_75t_L g12641 ( 
.A1(n_11619),
.A2(n_1119),
.B(n_1120),
.Y(n_12641)
);

NAND2xp5_ASAP7_75t_L g12642 ( 
.A(n_11091),
.B(n_1121),
.Y(n_12642)
);

NOR2xp33_ASAP7_75t_SL g12643 ( 
.A(n_10981),
.B(n_1121),
.Y(n_12643)
);

CKINVDCx5p33_ASAP7_75t_R g12644 ( 
.A(n_11590),
.Y(n_12644)
);

INVx2_ASAP7_75t_SL g12645 ( 
.A(n_11529),
.Y(n_12645)
);

NOR2xp33_ASAP7_75t_L g12646 ( 
.A(n_10971),
.B(n_1122),
.Y(n_12646)
);

INVx1_ASAP7_75t_L g12647 ( 
.A(n_10996),
.Y(n_12647)
);

NAND2xp5_ASAP7_75t_L g12648 ( 
.A(n_11091),
.B(n_1122),
.Y(n_12648)
);

BUFx2_ASAP7_75t_L g12649 ( 
.A(n_11178),
.Y(n_12649)
);

HB1xp67_ASAP7_75t_L g12650 ( 
.A(n_11180),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_10996),
.Y(n_12651)
);

OAI22xp5_ASAP7_75t_L g12652 ( 
.A1(n_11309),
.A2(n_1125),
.B1(n_1123),
.B2(n_1124),
.Y(n_12652)
);

NAND2xp5_ASAP7_75t_SL g12653 ( 
.A(n_11060),
.B(n_1123),
.Y(n_12653)
);

BUFx2_ASAP7_75t_L g12654 ( 
.A(n_11178),
.Y(n_12654)
);

AOI21xp5_ASAP7_75t_L g12655 ( 
.A1(n_11619),
.A2(n_1124),
.B(n_1125),
.Y(n_12655)
);

BUFx3_ASAP7_75t_L g12656 ( 
.A(n_11316),
.Y(n_12656)
);

NAND2xp5_ASAP7_75t_L g12657 ( 
.A(n_11091),
.B(n_1126),
.Y(n_12657)
);

A2O1A1Ixp33_ASAP7_75t_L g12658 ( 
.A1(n_10986),
.A2(n_1128),
.B(n_1126),
.C(n_1127),
.Y(n_12658)
);

NAND2xp5_ASAP7_75t_L g12659 ( 
.A(n_11091),
.B(n_1127),
.Y(n_12659)
);

NAND2xp33_ASAP7_75t_SL g12660 ( 
.A(n_11741),
.B(n_1128),
.Y(n_12660)
);

A2O1A1Ixp33_ASAP7_75t_L g12661 ( 
.A1(n_10986),
.A2(n_1131),
.B(n_1129),
.C(n_1130),
.Y(n_12661)
);

NOR2xp33_ASAP7_75t_L g12662 ( 
.A(n_10971),
.B(n_1129),
.Y(n_12662)
);

NAND2xp5_ASAP7_75t_L g12663 ( 
.A(n_11091),
.B(n_1130),
.Y(n_12663)
);

NOR2xp33_ASAP7_75t_L g12664 ( 
.A(n_10971),
.B(n_1131),
.Y(n_12664)
);

INVx2_ASAP7_75t_L g12665 ( 
.A(n_11267),
.Y(n_12665)
);

NOR2xp33_ASAP7_75t_L g12666 ( 
.A(n_10971),
.B(n_1132),
.Y(n_12666)
);

NOR3xp33_ASAP7_75t_SL g12667 ( 
.A(n_11366),
.B(n_1134),
.C(n_1135),
.Y(n_12667)
);

AOI21xp5_ASAP7_75t_L g12668 ( 
.A1(n_11619),
.A2(n_1134),
.B(n_1136),
.Y(n_12668)
);

NAND2xp5_ASAP7_75t_L g12669 ( 
.A(n_11091),
.B(n_1136),
.Y(n_12669)
);

INVx1_ASAP7_75t_L g12670 ( 
.A(n_10996),
.Y(n_12670)
);

NOR2xp33_ASAP7_75t_L g12671 ( 
.A(n_10971),
.B(n_1137),
.Y(n_12671)
);

BUFx3_ASAP7_75t_L g12672 ( 
.A(n_11316),
.Y(n_12672)
);

AOI21xp5_ASAP7_75t_L g12673 ( 
.A1(n_11619),
.A2(n_1137),
.B(n_1138),
.Y(n_12673)
);

NOR2xp33_ASAP7_75t_L g12674 ( 
.A(n_10971),
.B(n_1139),
.Y(n_12674)
);

A2O1A1Ixp33_ASAP7_75t_L g12675 ( 
.A1(n_10986),
.A2(n_1141),
.B(n_1139),
.C(n_1140),
.Y(n_12675)
);

INVx3_ASAP7_75t_L g12676 ( 
.A(n_11316),
.Y(n_12676)
);

AOI22xp33_ASAP7_75t_L g12677 ( 
.A1(n_11619),
.A2(n_1143),
.B1(n_1141),
.B2(n_1142),
.Y(n_12677)
);

HB1xp67_ASAP7_75t_L g12678 ( 
.A(n_11180),
.Y(n_12678)
);

AND2x2_ASAP7_75t_L g12679 ( 
.A(n_11487),
.B(n_1143),
.Y(n_12679)
);

NOR2xp33_ASAP7_75t_L g12680 ( 
.A(n_10971),
.B(n_1144),
.Y(n_12680)
);

INVx1_ASAP7_75t_L g12681 ( 
.A(n_10996),
.Y(n_12681)
);

OAI22xp5_ASAP7_75t_L g12682 ( 
.A1(n_11309),
.A2(n_1147),
.B1(n_1145),
.B2(n_1146),
.Y(n_12682)
);

AOI22xp33_ASAP7_75t_L g12683 ( 
.A1(n_11619),
.A2(n_1147),
.B1(n_1145),
.B2(n_1146),
.Y(n_12683)
);

AOI22x1_ASAP7_75t_L g12684 ( 
.A1(n_11677),
.A2(n_1150),
.B1(n_1148),
.B2(n_1149),
.Y(n_12684)
);

OR2x2_ASAP7_75t_L g12685 ( 
.A(n_10996),
.B(n_1148),
.Y(n_12685)
);

OAI22xp5_ASAP7_75t_L g12686 ( 
.A1(n_11309),
.A2(n_1151),
.B1(n_1149),
.B2(n_1150),
.Y(n_12686)
);

NAND2xp5_ASAP7_75t_SL g12687 ( 
.A(n_11060),
.B(n_1151),
.Y(n_12687)
);

NAND2xp5_ASAP7_75t_L g12688 ( 
.A(n_11091),
.B(n_1152),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_10996),
.Y(n_12689)
);

AO31x2_ASAP7_75t_L g12690 ( 
.A1(n_12112),
.A2(n_1154),
.A3(n_1152),
.B(n_1153),
.Y(n_12690)
);

INVx1_ASAP7_75t_L g12691 ( 
.A(n_11975),
.Y(n_12691)
);

OAI21xp33_ASAP7_75t_L g12692 ( 
.A1(n_11935),
.A2(n_1154),
.B(n_1155),
.Y(n_12692)
);

NAND2xp5_ASAP7_75t_L g12693 ( 
.A(n_12561),
.B(n_1155),
.Y(n_12693)
);

INVx2_ASAP7_75t_L g12694 ( 
.A(n_11822),
.Y(n_12694)
);

INVx1_ASAP7_75t_L g12695 ( 
.A(n_11978),
.Y(n_12695)
);

OAI21xp5_ASAP7_75t_L g12696 ( 
.A1(n_11752),
.A2(n_1156),
.B(n_1157),
.Y(n_12696)
);

OA21x2_ASAP7_75t_L g12697 ( 
.A1(n_12313),
.A2(n_1156),
.B(n_1158),
.Y(n_12697)
);

AO31x2_ASAP7_75t_L g12698 ( 
.A1(n_12113),
.A2(n_1161),
.A3(n_1159),
.B(n_1160),
.Y(n_12698)
);

AOI31xp67_ASAP7_75t_L g12699 ( 
.A1(n_11944),
.A2(n_1161),
.A3(n_1159),
.B(n_1160),
.Y(n_12699)
);

AND2x2_ASAP7_75t_L g12700 ( 
.A(n_11777),
.B(n_1162),
.Y(n_12700)
);

NAND2xp5_ASAP7_75t_L g12701 ( 
.A(n_12570),
.B(n_1162),
.Y(n_12701)
);

OAI21x1_ASAP7_75t_L g12702 ( 
.A1(n_12147),
.A2(n_1163),
.B(n_1164),
.Y(n_12702)
);

NAND2xp5_ASAP7_75t_L g12703 ( 
.A(n_11790),
.B(n_1163),
.Y(n_12703)
);

NAND2xp5_ASAP7_75t_L g12704 ( 
.A(n_12678),
.B(n_1164),
.Y(n_12704)
);

AND2x4_ASAP7_75t_L g12705 ( 
.A(n_12552),
.B(n_1165),
.Y(n_12705)
);

OAI21x1_ASAP7_75t_L g12706 ( 
.A1(n_11904),
.A2(n_1165),
.B(n_1166),
.Y(n_12706)
);

BUFx12f_ASAP7_75t_L g12707 ( 
.A(n_11841),
.Y(n_12707)
);

INVx1_ASAP7_75t_L g12708 ( 
.A(n_11983),
.Y(n_12708)
);

AOI21xp5_ASAP7_75t_L g12709 ( 
.A1(n_11912),
.A2(n_1167),
.B(n_1168),
.Y(n_12709)
);

OAI21x1_ASAP7_75t_L g12710 ( 
.A1(n_11941),
.A2(n_1169),
.B(n_1170),
.Y(n_12710)
);

NAND2x1p5_ASAP7_75t_L g12711 ( 
.A(n_12048),
.B(n_1169),
.Y(n_12711)
);

OA21x2_ASAP7_75t_L g12712 ( 
.A1(n_12324),
.A2(n_1170),
.B(n_1171),
.Y(n_12712)
);

INVx1_ASAP7_75t_L g12713 ( 
.A(n_11989),
.Y(n_12713)
);

OAI21x1_ASAP7_75t_L g12714 ( 
.A1(n_12403),
.A2(n_1171),
.B(n_1172),
.Y(n_12714)
);

AOI221x1_ASAP7_75t_L g12715 ( 
.A1(n_12047),
.A2(n_1175),
.B1(n_1173),
.B2(n_1174),
.C(n_1176),
.Y(n_12715)
);

AND2x2_ASAP7_75t_L g12716 ( 
.A(n_12574),
.B(n_1173),
.Y(n_12716)
);

AND2x2_ASAP7_75t_L g12717 ( 
.A(n_12576),
.B(n_1174),
.Y(n_12717)
);

OAI22xp5_ASAP7_75t_L g12718 ( 
.A1(n_12051),
.A2(n_1177),
.B1(n_1175),
.B2(n_1176),
.Y(n_12718)
);

NAND2xp5_ASAP7_75t_SL g12719 ( 
.A(n_12048),
.B(n_1177),
.Y(n_12719)
);

AO31x2_ASAP7_75t_L g12720 ( 
.A1(n_12088),
.A2(n_1180),
.A3(n_1178),
.B(n_1179),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_11783),
.B(n_1178),
.Y(n_12721)
);

NAND2xp5_ASAP7_75t_L g12722 ( 
.A(n_12650),
.B(n_1179),
.Y(n_12722)
);

OAI21x1_ASAP7_75t_L g12723 ( 
.A1(n_12053),
.A2(n_1181),
.B(n_1182),
.Y(n_12723)
);

AOI21x1_ASAP7_75t_L g12724 ( 
.A1(n_11954),
.A2(n_1183),
.B(n_1184),
.Y(n_12724)
);

NAND3xp33_ASAP7_75t_L g12725 ( 
.A(n_11760),
.B(n_1183),
.C(n_1185),
.Y(n_12725)
);

OAI21xp5_ASAP7_75t_L g12726 ( 
.A1(n_11784),
.A2(n_11782),
.B(n_11774),
.Y(n_12726)
);

NAND2xp5_ASAP7_75t_L g12727 ( 
.A(n_12097),
.B(n_12095),
.Y(n_12727)
);

INVx1_ASAP7_75t_L g12728 ( 
.A(n_11998),
.Y(n_12728)
);

AOI21xp5_ASAP7_75t_SL g12729 ( 
.A1(n_11795),
.A2(n_1186),
.B(n_1187),
.Y(n_12729)
);

AOI21xp5_ASAP7_75t_L g12730 ( 
.A1(n_12475),
.A2(n_1186),
.B(n_1187),
.Y(n_12730)
);

AO31x2_ASAP7_75t_L g12731 ( 
.A1(n_11785),
.A2(n_1191),
.A3(n_1189),
.B(n_1190),
.Y(n_12731)
);

OAI21x1_ASAP7_75t_L g12732 ( 
.A1(n_12399),
.A2(n_1189),
.B(n_1190),
.Y(n_12732)
);

NOR2x1_ASAP7_75t_SL g12733 ( 
.A(n_12354),
.B(n_1191),
.Y(n_12733)
);

NAND2xp5_ASAP7_75t_L g12734 ( 
.A(n_12308),
.B(n_1192),
.Y(n_12734)
);

NAND2xp5_ASAP7_75t_L g12735 ( 
.A(n_11770),
.B(n_1193),
.Y(n_12735)
);

AOI21xp5_ASAP7_75t_L g12736 ( 
.A1(n_12334),
.A2(n_1193),
.B(n_1194),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_11771),
.B(n_1194),
.Y(n_12737)
);

AO31x2_ASAP7_75t_L g12738 ( 
.A1(n_12039),
.A2(n_1197),
.A3(n_1195),
.B(n_1196),
.Y(n_12738)
);

AOI21xp5_ASAP7_75t_L g12739 ( 
.A1(n_11939),
.A2(n_1195),
.B(n_1196),
.Y(n_12739)
);

INVx3_ASAP7_75t_L g12740 ( 
.A(n_11798),
.Y(n_12740)
);

NAND2xp5_ASAP7_75t_L g12741 ( 
.A(n_11779),
.B(n_1197),
.Y(n_12741)
);

INVx2_ASAP7_75t_L g12742 ( 
.A(n_11863),
.Y(n_12742)
);

NAND2xp5_ASAP7_75t_L g12743 ( 
.A(n_12649),
.B(n_1198),
.Y(n_12743)
);

NAND2xp5_ASAP7_75t_L g12744 ( 
.A(n_12654),
.B(n_1198),
.Y(n_12744)
);

OA21x2_ASAP7_75t_L g12745 ( 
.A1(n_11899),
.A2(n_1199),
.B(n_1200),
.Y(n_12745)
);

NAND3xp33_ASAP7_75t_L g12746 ( 
.A(n_11829),
.B(n_1199),
.C(n_1200),
.Y(n_12746)
);

OAI21x1_ASAP7_75t_L g12747 ( 
.A1(n_12316),
.A2(n_1201),
.B(n_1202),
.Y(n_12747)
);

OA21x2_ASAP7_75t_L g12748 ( 
.A1(n_11794),
.A2(n_11950),
.B(n_11974),
.Y(n_12748)
);

HB1xp67_ASAP7_75t_L g12749 ( 
.A(n_12108),
.Y(n_12749)
);

OAI21x1_ASAP7_75t_L g12750 ( 
.A1(n_12240),
.A2(n_1201),
.B(n_1202),
.Y(n_12750)
);

INVx2_ASAP7_75t_L g12751 ( 
.A(n_11864),
.Y(n_12751)
);

BUFx6f_ASAP7_75t_L g12752 ( 
.A(n_12037),
.Y(n_12752)
);

OAI21x1_ASAP7_75t_L g12753 ( 
.A1(n_12421),
.A2(n_1203),
.B(n_1204),
.Y(n_12753)
);

AOI21xp5_ASAP7_75t_L g12754 ( 
.A1(n_11979),
.A2(n_1203),
.B(n_1204),
.Y(n_12754)
);

OAI21x1_ASAP7_75t_L g12755 ( 
.A1(n_12472),
.A2(n_1205),
.B(n_1206),
.Y(n_12755)
);

AOI21xp5_ASAP7_75t_L g12756 ( 
.A1(n_12066),
.A2(n_1205),
.B(n_1206),
.Y(n_12756)
);

AOI21xp5_ASAP7_75t_L g12757 ( 
.A1(n_11961),
.A2(n_1207),
.B(n_1208),
.Y(n_12757)
);

INVx1_ASAP7_75t_L g12758 ( 
.A(n_12000),
.Y(n_12758)
);

OAI21x1_ASAP7_75t_L g12759 ( 
.A1(n_12479),
.A2(n_1207),
.B(n_1208),
.Y(n_12759)
);

INVx5_ASAP7_75t_L g12760 ( 
.A(n_12065),
.Y(n_12760)
);

OAI21x1_ASAP7_75t_L g12761 ( 
.A1(n_11977),
.A2(n_1209),
.B(n_1210),
.Y(n_12761)
);

INVx1_ASAP7_75t_SL g12762 ( 
.A(n_11873),
.Y(n_12762)
);

NOR2xp33_ASAP7_75t_L g12763 ( 
.A(n_12345),
.B(n_1209),
.Y(n_12763)
);

OAI21x1_ASAP7_75t_L g12764 ( 
.A1(n_12468),
.A2(n_1210),
.B(n_1211),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_11808),
.B(n_1211),
.Y(n_12765)
);

NAND2xp5_ASAP7_75t_L g12766 ( 
.A(n_11819),
.B(n_1212),
.Y(n_12766)
);

AO31x2_ASAP7_75t_L g12767 ( 
.A1(n_12505),
.A2(n_12534),
.A3(n_12151),
.B(n_12529),
.Y(n_12767)
);

BUFx2_ASAP7_75t_L g12768 ( 
.A(n_11796),
.Y(n_12768)
);

NAND2xp5_ASAP7_75t_L g12769 ( 
.A(n_11832),
.B(n_1212),
.Y(n_12769)
);

INVx1_ASAP7_75t_SL g12770 ( 
.A(n_12551),
.Y(n_12770)
);

BUFx6f_ASAP7_75t_L g12771 ( 
.A(n_12037),
.Y(n_12771)
);

AOI21xp5_ASAP7_75t_L g12772 ( 
.A1(n_12251),
.A2(n_1213),
.B(n_1214),
.Y(n_12772)
);

AOI21xp5_ASAP7_75t_L g12773 ( 
.A1(n_12335),
.A2(n_1214),
.B(n_1215),
.Y(n_12773)
);

A2O1A1Ixp33_ASAP7_75t_L g12774 ( 
.A1(n_12040),
.A2(n_1218),
.B(n_1216),
.C(n_1217),
.Y(n_12774)
);

NAND2xp5_ASAP7_75t_L g12775 ( 
.A(n_11839),
.B(n_1216),
.Y(n_12775)
);

AOI21xp5_ASAP7_75t_L g12776 ( 
.A1(n_12506),
.A2(n_1217),
.B(n_1218),
.Y(n_12776)
);

INVxp67_ASAP7_75t_L g12777 ( 
.A(n_12370),
.Y(n_12777)
);

AOI21xp5_ASAP7_75t_L g12778 ( 
.A1(n_12509),
.A2(n_1219),
.B(n_1220),
.Y(n_12778)
);

OAI21x1_ASAP7_75t_L g12779 ( 
.A1(n_12253),
.A2(n_1219),
.B(n_1220),
.Y(n_12779)
);

INVx3_ASAP7_75t_L g12780 ( 
.A(n_11837),
.Y(n_12780)
);

NAND2xp5_ASAP7_75t_SL g12781 ( 
.A(n_12222),
.B(n_1221),
.Y(n_12781)
);

NOR2xp33_ASAP7_75t_L g12782 ( 
.A(n_12345),
.B(n_1222),
.Y(n_12782)
);

OAI21x1_ASAP7_75t_L g12783 ( 
.A1(n_12296),
.A2(n_1222),
.B(n_1223),
.Y(n_12783)
);

AOI21xp5_ASAP7_75t_L g12784 ( 
.A1(n_12526),
.A2(n_1223),
.B(n_1224),
.Y(n_12784)
);

AOI21xp5_ASAP7_75t_L g12785 ( 
.A1(n_12535),
.A2(n_1224),
.B(n_1225),
.Y(n_12785)
);

AOI21xp5_ASAP7_75t_L g12786 ( 
.A1(n_12538),
.A2(n_1226),
.B(n_1227),
.Y(n_12786)
);

NAND3xp33_ASAP7_75t_SL g12787 ( 
.A(n_12130),
.B(n_1227),
.C(n_1228),
.Y(n_12787)
);

AOI21xp5_ASAP7_75t_L g12788 ( 
.A1(n_12542),
.A2(n_1228),
.B(n_1229),
.Y(n_12788)
);

INVx2_ASAP7_75t_L g12789 ( 
.A(n_11878),
.Y(n_12789)
);

NOR2xp67_ASAP7_75t_L g12790 ( 
.A(n_11906),
.B(n_1229),
.Y(n_12790)
);

INVx1_ASAP7_75t_L g12791 ( 
.A(n_11883),
.Y(n_12791)
);

OAI22xp5_ASAP7_75t_L g12792 ( 
.A1(n_12008),
.A2(n_11844),
.B1(n_12273),
.B2(n_12077),
.Y(n_12792)
);

NOR2xp33_ASAP7_75t_L g12793 ( 
.A(n_12273),
.B(n_1230),
.Y(n_12793)
);

OAI22xp5_ASAP7_75t_L g12794 ( 
.A1(n_12059),
.A2(n_1232),
.B1(n_1230),
.B2(n_1231),
.Y(n_12794)
);

OAI21x1_ASAP7_75t_L g12795 ( 
.A1(n_12200),
.A2(n_12355),
.B(n_11914),
.Y(n_12795)
);

A2O1A1Ixp33_ASAP7_75t_L g12796 ( 
.A1(n_12580),
.A2(n_1233),
.B(n_1231),
.C(n_1232),
.Y(n_12796)
);

OAI21x1_ASAP7_75t_L g12797 ( 
.A1(n_12404),
.A2(n_1233),
.B(n_1234),
.Y(n_12797)
);

OAI21xp5_ASAP7_75t_L g12798 ( 
.A1(n_11792),
.A2(n_1234),
.B(n_1235),
.Y(n_12798)
);

AO31x2_ASAP7_75t_L g12799 ( 
.A1(n_12515),
.A2(n_1238),
.A3(n_1236),
.B(n_1237),
.Y(n_12799)
);

AOI21xp33_ASAP7_75t_L g12800 ( 
.A1(n_11946),
.A2(n_1236),
.B(n_1237),
.Y(n_12800)
);

AOI21xp5_ASAP7_75t_L g12801 ( 
.A1(n_12550),
.A2(n_12575),
.B(n_12564),
.Y(n_12801)
);

BUFx2_ASAP7_75t_L g12802 ( 
.A(n_11917),
.Y(n_12802)
);

INVx2_ASAP7_75t_L g12803 ( 
.A(n_11885),
.Y(n_12803)
);

AND2x4_ASAP7_75t_L g12804 ( 
.A(n_12067),
.B(n_1238),
.Y(n_12804)
);

AO21x2_ASAP7_75t_L g12805 ( 
.A1(n_11945),
.A2(n_1239),
.B(n_1240),
.Y(n_12805)
);

OAI21x1_ASAP7_75t_L g12806 ( 
.A1(n_12124),
.A2(n_1239),
.B(n_1240),
.Y(n_12806)
);

NOR4xp25_ASAP7_75t_L g12807 ( 
.A(n_12281),
.B(n_1243),
.C(n_1241),
.D(n_1242),
.Y(n_12807)
);

AOI21xp5_ASAP7_75t_L g12808 ( 
.A1(n_12578),
.A2(n_1241),
.B(n_1242),
.Y(n_12808)
);

AOI21xp5_ASAP7_75t_L g12809 ( 
.A1(n_12579),
.A2(n_1243),
.B(n_1244),
.Y(n_12809)
);

OAI21x1_ASAP7_75t_L g12810 ( 
.A1(n_12371),
.A2(n_1244),
.B(n_1245),
.Y(n_12810)
);

A2O1A1Ixp33_ASAP7_75t_L g12811 ( 
.A1(n_12373),
.A2(n_1247),
.B(n_1245),
.C(n_1246),
.Y(n_12811)
);

NAND2x1p5_ASAP7_75t_L g12812 ( 
.A(n_12222),
.B(n_1246),
.Y(n_12812)
);

AOI21xp5_ASAP7_75t_L g12813 ( 
.A1(n_12603),
.A2(n_1247),
.B(n_1248),
.Y(n_12813)
);

OAI21xp5_ASAP7_75t_L g12814 ( 
.A1(n_11812),
.A2(n_11817),
.B(n_11813),
.Y(n_12814)
);

AOI21xp5_ASAP7_75t_L g12815 ( 
.A1(n_12605),
.A2(n_1249),
.B(n_1250),
.Y(n_12815)
);

NAND2xp5_ASAP7_75t_L g12816 ( 
.A(n_11842),
.B(n_1250),
.Y(n_12816)
);

A2O1A1Ixp33_ASAP7_75t_L g12817 ( 
.A1(n_11754),
.A2(n_12502),
.B(n_12516),
.C(n_12618),
.Y(n_12817)
);

AOI21xp5_ASAP7_75t_L g12818 ( 
.A1(n_12625),
.A2(n_1251),
.B(n_1252),
.Y(n_12818)
);

AOI21x1_ASAP7_75t_SL g12819 ( 
.A1(n_12474),
.A2(n_1252),
.B(n_1254),
.Y(n_12819)
);

OAI21x1_ASAP7_75t_L g12820 ( 
.A1(n_11768),
.A2(n_1255),
.B(n_1256),
.Y(n_12820)
);

AOI21xp5_ASAP7_75t_L g12821 ( 
.A1(n_12627),
.A2(n_1255),
.B(n_1256),
.Y(n_12821)
);

AOI21xp33_ASAP7_75t_L g12822 ( 
.A1(n_11993),
.A2(n_1257),
.B(n_1258),
.Y(n_12822)
);

AO22x2_ASAP7_75t_L g12823 ( 
.A1(n_11849),
.A2(n_1260),
.B1(n_1258),
.B2(n_1259),
.Y(n_12823)
);

AO31x2_ASAP7_75t_L g12824 ( 
.A1(n_12537),
.A2(n_1262),
.A3(n_1259),
.B(n_1261),
.Y(n_12824)
);

AND2x4_ASAP7_75t_L g12825 ( 
.A(n_11924),
.B(n_1261),
.Y(n_12825)
);

BUFx4_ASAP7_75t_SL g12826 ( 
.A(n_11986),
.Y(n_12826)
);

OAI21x1_ASAP7_75t_L g12827 ( 
.A1(n_12213),
.A2(n_1262),
.B(n_1263),
.Y(n_12827)
);

INVx1_ASAP7_75t_L g12828 ( 
.A(n_11887),
.Y(n_12828)
);

OAI21x1_ASAP7_75t_L g12829 ( 
.A1(n_12489),
.A2(n_1263),
.B(n_1264),
.Y(n_12829)
);

OAI21x1_ASAP7_75t_L g12830 ( 
.A1(n_12492),
.A2(n_1264),
.B(n_1265),
.Y(n_12830)
);

HB1xp67_ASAP7_75t_L g12831 ( 
.A(n_11919),
.Y(n_12831)
);

CKINVDCx8_ASAP7_75t_R g12832 ( 
.A(n_11799),
.Y(n_12832)
);

INVx2_ASAP7_75t_L g12833 ( 
.A(n_11894),
.Y(n_12833)
);

OAI21x1_ASAP7_75t_SL g12834 ( 
.A1(n_11831),
.A2(n_1265),
.B(n_1266),
.Y(n_12834)
);

OA21x2_ASAP7_75t_L g12835 ( 
.A1(n_12231),
.A2(n_1267),
.B(n_1268),
.Y(n_12835)
);

OAI21x1_ASAP7_75t_L g12836 ( 
.A1(n_12493),
.A2(n_1267),
.B(n_1269),
.Y(n_12836)
);

INVx1_ASAP7_75t_L g12837 ( 
.A(n_11907),
.Y(n_12837)
);

OAI21x1_ASAP7_75t_L g12838 ( 
.A1(n_12566),
.A2(n_1269),
.B(n_1270),
.Y(n_12838)
);

AO21x1_ASAP7_75t_L g12839 ( 
.A1(n_11925),
.A2(n_12660),
.B(n_12072),
.Y(n_12839)
);

INVx1_ASAP7_75t_L g12840 ( 
.A(n_11909),
.Y(n_12840)
);

OAI21x1_ASAP7_75t_SL g12841 ( 
.A1(n_12333),
.A2(n_1271),
.B(n_1272),
.Y(n_12841)
);

INVx1_ASAP7_75t_L g12842 ( 
.A(n_11934),
.Y(n_12842)
);

INVx1_ASAP7_75t_L g12843 ( 
.A(n_11952),
.Y(n_12843)
);

NAND2xp5_ASAP7_75t_L g12844 ( 
.A(n_11859),
.B(n_1272),
.Y(n_12844)
);

OAI22xp5_ASAP7_75t_L g12845 ( 
.A1(n_12090),
.A2(n_1275),
.B1(n_1273),
.B2(n_1274),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_11862),
.B(n_1273),
.Y(n_12846)
);

INVxp67_ASAP7_75t_L g12847 ( 
.A(n_12377),
.Y(n_12847)
);

OAI21xp5_ASAP7_75t_L g12848 ( 
.A1(n_11823),
.A2(n_1274),
.B(n_1275),
.Y(n_12848)
);

NOR2xp67_ASAP7_75t_SL g12849 ( 
.A(n_12234),
.B(n_12629),
.Y(n_12849)
);

INVx1_ASAP7_75t_L g12850 ( 
.A(n_11953),
.Y(n_12850)
);

INVx1_ASAP7_75t_L g12851 ( 
.A(n_11807),
.Y(n_12851)
);

OA21x2_ASAP7_75t_L g12852 ( 
.A1(n_11800),
.A2(n_1276),
.B(n_1277),
.Y(n_12852)
);

OAI21xp5_ASAP7_75t_L g12853 ( 
.A1(n_11824),
.A2(n_1276),
.B(n_1277),
.Y(n_12853)
);

NAND2xp5_ASAP7_75t_SL g12854 ( 
.A(n_12354),
.B(n_1278),
.Y(n_12854)
);

OAI21x1_ASAP7_75t_L g12855 ( 
.A1(n_12485),
.A2(n_1278),
.B(n_1279),
.Y(n_12855)
);

OAI21x1_ASAP7_75t_L g12856 ( 
.A1(n_12497),
.A2(n_1280),
.B(n_1281),
.Y(n_12856)
);

INVx1_ASAP7_75t_L g12857 ( 
.A(n_11879),
.Y(n_12857)
);

OAI21xp5_ASAP7_75t_L g12858 ( 
.A1(n_11827),
.A2(n_1280),
.B(n_1281),
.Y(n_12858)
);

A2O1A1Ixp33_ASAP7_75t_L g12859 ( 
.A1(n_12633),
.A2(n_1284),
.B(n_1282),
.C(n_1283),
.Y(n_12859)
);

AND2x2_ASAP7_75t_L g12860 ( 
.A(n_11868),
.B(n_1282),
.Y(n_12860)
);

OAI21x1_ASAP7_75t_L g12861 ( 
.A1(n_12430),
.A2(n_1283),
.B(n_1284),
.Y(n_12861)
);

AND2x2_ASAP7_75t_L g12862 ( 
.A(n_11836),
.B(n_1285),
.Y(n_12862)
);

INVx1_ASAP7_75t_L g12863 ( 
.A(n_11884),
.Y(n_12863)
);

NAND2xp5_ASAP7_75t_L g12864 ( 
.A(n_11889),
.B(n_1285),
.Y(n_12864)
);

NAND2xp5_ASAP7_75t_L g12865 ( 
.A(n_11903),
.B(n_1286),
.Y(n_12865)
);

OAI21x1_ASAP7_75t_L g12866 ( 
.A1(n_11828),
.A2(n_1286),
.B(n_1287),
.Y(n_12866)
);

BUFx6f_ASAP7_75t_L g12867 ( 
.A(n_12050),
.Y(n_12867)
);

OR2x2_ASAP7_75t_L g12868 ( 
.A(n_11937),
.B(n_1287),
.Y(n_12868)
);

OAI21xp5_ASAP7_75t_L g12869 ( 
.A1(n_11840),
.A2(n_1288),
.B(n_1289),
.Y(n_12869)
);

AO31x2_ASAP7_75t_L g12870 ( 
.A1(n_12553),
.A2(n_1290),
.A3(n_1288),
.B(n_1289),
.Y(n_12870)
);

OAI21x1_ASAP7_75t_L g12871 ( 
.A1(n_11865),
.A2(n_1290),
.B(n_1291),
.Y(n_12871)
);

AO32x2_ASAP7_75t_L g12872 ( 
.A1(n_12353),
.A2(n_1294),
.A3(n_1292),
.B1(n_1293),
.B2(n_1295),
.Y(n_12872)
);

CKINVDCx8_ASAP7_75t_R g12873 ( 
.A(n_12290),
.Y(n_12873)
);

OAI21x1_ASAP7_75t_L g12874 ( 
.A1(n_11877),
.A2(n_1293),
.B(n_1294),
.Y(n_12874)
);

OAI22xp5_ASAP7_75t_L g12875 ( 
.A1(n_12115),
.A2(n_12637),
.B1(n_12632),
.B2(n_12608),
.Y(n_12875)
);

NAND2xp5_ASAP7_75t_L g12876 ( 
.A(n_12558),
.B(n_1295),
.Y(n_12876)
);

INVx1_ASAP7_75t_L g12877 ( 
.A(n_12565),
.Y(n_12877)
);

NAND2xp5_ASAP7_75t_L g12878 ( 
.A(n_12569),
.B(n_1296),
.Y(n_12878)
);

NAND2xp5_ASAP7_75t_L g12879 ( 
.A(n_12583),
.B(n_1296),
.Y(n_12879)
);

OAI21x1_ASAP7_75t_L g12880 ( 
.A1(n_11881),
.A2(n_11910),
.B(n_11893),
.Y(n_12880)
);

NAND3xp33_ASAP7_75t_L g12881 ( 
.A(n_11922),
.B(n_1297),
.C(n_1298),
.Y(n_12881)
);

NAND2xp5_ASAP7_75t_L g12882 ( 
.A(n_12588),
.B(n_1299),
.Y(n_12882)
);

AOI22xp5_ASAP7_75t_L g12883 ( 
.A1(n_12209),
.A2(n_1302),
.B1(n_1300),
.B2(n_1301),
.Y(n_12883)
);

OAI21x1_ASAP7_75t_L g12884 ( 
.A1(n_11927),
.A2(n_1300),
.B(n_1302),
.Y(n_12884)
);

AOI21xp5_ASAP7_75t_L g12885 ( 
.A1(n_12641),
.A2(n_12668),
.B(n_12655),
.Y(n_12885)
);

AOI22xp5_ASAP7_75t_L g12886 ( 
.A1(n_12591),
.A2(n_1305),
.B1(n_1303),
.B2(n_1304),
.Y(n_12886)
);

AND2x2_ASAP7_75t_L g12887 ( 
.A(n_12590),
.B(n_1303),
.Y(n_12887)
);

AOI221x1_ASAP7_75t_L g12888 ( 
.A1(n_12673),
.A2(n_1306),
.B1(n_1304),
.B2(n_1305),
.C(n_1307),
.Y(n_12888)
);

OAI21x1_ASAP7_75t_L g12889 ( 
.A1(n_11931),
.A2(n_1306),
.B(n_1307),
.Y(n_12889)
);

NAND2xp5_ASAP7_75t_SL g12890 ( 
.A(n_12423),
.B(n_12243),
.Y(n_12890)
);

BUFx6f_ASAP7_75t_L g12891 ( 
.A(n_12050),
.Y(n_12891)
);

NAND3xp33_ASAP7_75t_SL g12892 ( 
.A(n_12043),
.B(n_1308),
.C(n_1309),
.Y(n_12892)
);

NAND2xp5_ASAP7_75t_L g12893 ( 
.A(n_12621),
.B(n_1308),
.Y(n_12893)
);

A2O1A1Ixp33_ASAP7_75t_L g12894 ( 
.A1(n_12315),
.A2(n_1312),
.B(n_1310),
.C(n_1311),
.Y(n_12894)
);

INVx1_ASAP7_75t_L g12895 ( 
.A(n_12631),
.Y(n_12895)
);

CKINVDCx5p33_ASAP7_75t_R g12896 ( 
.A(n_12547),
.Y(n_12896)
);

AOI21xp5_ASAP7_75t_L g12897 ( 
.A1(n_12494),
.A2(n_1310),
.B(n_1311),
.Y(n_12897)
);

AOI21xp5_ASAP7_75t_L g12898 ( 
.A1(n_11955),
.A2(n_1312),
.B(n_1313),
.Y(n_12898)
);

OAI21x1_ASAP7_75t_L g12899 ( 
.A1(n_11964),
.A2(n_1313),
.B(n_1314),
.Y(n_12899)
);

NAND2xp5_ASAP7_75t_L g12900 ( 
.A(n_12647),
.B(n_1314),
.Y(n_12900)
);

AOI21xp5_ASAP7_75t_L g12901 ( 
.A1(n_11970),
.A2(n_1315),
.B(n_1316),
.Y(n_12901)
);

AOI21xp5_ASAP7_75t_L g12902 ( 
.A1(n_11802),
.A2(n_1315),
.B(n_1316),
.Y(n_12902)
);

NAND2xp5_ASAP7_75t_L g12903 ( 
.A(n_12651),
.B(n_1317),
.Y(n_12903)
);

NAND2xp5_ASAP7_75t_L g12904 ( 
.A(n_12670),
.B(n_1317),
.Y(n_12904)
);

INVx2_ASAP7_75t_L g12905 ( 
.A(n_12681),
.Y(n_12905)
);

AO31x2_ASAP7_75t_L g12906 ( 
.A1(n_12573),
.A2(n_1320),
.A3(n_1318),
.B(n_1319),
.Y(n_12906)
);

OR2x2_ASAP7_75t_L g12907 ( 
.A(n_12689),
.B(n_1318),
.Y(n_12907)
);

AND2x4_ASAP7_75t_L g12908 ( 
.A(n_12099),
.B(n_1319),
.Y(n_12908)
);

AOI21xp5_ASAP7_75t_L g12909 ( 
.A1(n_12545),
.A2(n_12146),
.B(n_12084),
.Y(n_12909)
);

INVxp67_ASAP7_75t_SL g12910 ( 
.A(n_11757),
.Y(n_12910)
);

INVx2_ASAP7_75t_SL g12911 ( 
.A(n_12104),
.Y(n_12911)
);

CKINVDCx14_ASAP7_75t_R g12912 ( 
.A(n_12269),
.Y(n_12912)
);

NAND2xp5_ASAP7_75t_L g12913 ( 
.A(n_12321),
.B(n_1321),
.Y(n_12913)
);

NOR2xp67_ASAP7_75t_L g12914 ( 
.A(n_11906),
.B(n_1322),
.Y(n_12914)
);

OAI21xp33_ASAP7_75t_L g12915 ( 
.A1(n_11852),
.A2(n_1322),
.B(n_1323),
.Y(n_12915)
);

AOI21xp5_ASAP7_75t_L g12916 ( 
.A1(n_12192),
.A2(n_1323),
.B(n_1324),
.Y(n_12916)
);

NAND2xp5_ASAP7_75t_L g12917 ( 
.A(n_12358),
.B(n_1324),
.Y(n_12917)
);

INVx3_ASAP7_75t_L g12918 ( 
.A(n_12143),
.Y(n_12918)
);

NAND2xp5_ASAP7_75t_SL g12919 ( 
.A(n_12423),
.B(n_1325),
.Y(n_12919)
);

AO22x2_ASAP7_75t_L g12920 ( 
.A1(n_11895),
.A2(n_1327),
.B1(n_1325),
.B2(n_1326),
.Y(n_12920)
);

NOR2xp33_ASAP7_75t_L g12921 ( 
.A(n_12078),
.B(n_1326),
.Y(n_12921)
);

AO32x2_ASAP7_75t_L g12922 ( 
.A1(n_12013),
.A2(n_12364),
.A3(n_12080),
.B1(n_12070),
.B2(n_12378),
.Y(n_12922)
);

AOI21xp5_ASAP7_75t_L g12923 ( 
.A1(n_12442),
.A2(n_1328),
.B(n_1329),
.Y(n_12923)
);

INVx1_ASAP7_75t_L g12924 ( 
.A(n_12006),
.Y(n_12924)
);

NAND2xp5_ASAP7_75t_L g12925 ( 
.A(n_12360),
.B(n_1328),
.Y(n_12925)
);

A2O1A1Ixp33_ASAP7_75t_L g12926 ( 
.A1(n_11958),
.A2(n_1331),
.B(n_1329),
.C(n_1330),
.Y(n_12926)
);

AO31x2_ASAP7_75t_L g12927 ( 
.A1(n_12586),
.A2(n_1332),
.A3(n_1330),
.B(n_1331),
.Y(n_12927)
);

NOR4xp25_ASAP7_75t_L g12928 ( 
.A(n_12145),
.B(n_1334),
.C(n_1332),
.D(n_1333),
.Y(n_12928)
);

INVx2_ASAP7_75t_SL g12929 ( 
.A(n_12104),
.Y(n_12929)
);

AO31x2_ASAP7_75t_L g12930 ( 
.A1(n_12614),
.A2(n_1335),
.A3(n_1333),
.B(n_1334),
.Y(n_12930)
);

BUFx3_ASAP7_75t_L g12931 ( 
.A(n_12517),
.Y(n_12931)
);

NAND2xp5_ASAP7_75t_L g12932 ( 
.A(n_12341),
.B(n_1335),
.Y(n_12932)
);

INVx1_ASAP7_75t_L g12933 ( 
.A(n_12011),
.Y(n_12933)
);

INVx2_ASAP7_75t_L g12934 ( 
.A(n_11766),
.Y(n_12934)
);

NAND2xp5_ASAP7_75t_L g12935 ( 
.A(n_12349),
.B(n_1336),
.Y(n_12935)
);

AND2x2_ASAP7_75t_L g12936 ( 
.A(n_12439),
.B(n_1336),
.Y(n_12936)
);

AOI21xp5_ASAP7_75t_L g12937 ( 
.A1(n_11956),
.A2(n_1337),
.B(n_1338),
.Y(n_12937)
);

AO31x2_ASAP7_75t_L g12938 ( 
.A1(n_12635),
.A2(n_1339),
.A3(n_1337),
.B(n_1338),
.Y(n_12938)
);

INVxp67_ASAP7_75t_SL g12939 ( 
.A(n_12519),
.Y(n_12939)
);

OAI21x1_ASAP7_75t_L g12940 ( 
.A1(n_12076),
.A2(n_1339),
.B(n_1340),
.Y(n_12940)
);

NAND2xp5_ASAP7_75t_L g12941 ( 
.A(n_12365),
.B(n_1340),
.Y(n_12941)
);

BUFx3_ASAP7_75t_L g12942 ( 
.A(n_11890),
.Y(n_12942)
);

AND2x2_ASAP7_75t_SL g12943 ( 
.A(n_12233),
.B(n_1341),
.Y(n_12943)
);

HB1xp67_ASAP7_75t_L g12944 ( 
.A(n_12520),
.Y(n_12944)
);

NAND2xp5_ASAP7_75t_L g12945 ( 
.A(n_12367),
.B(n_1341),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12018),
.Y(n_12946)
);

OAI21x1_ASAP7_75t_L g12947 ( 
.A1(n_12026),
.A2(n_1342),
.B(n_1343),
.Y(n_12947)
);

INVx1_ASAP7_75t_L g12948 ( 
.A(n_12062),
.Y(n_12948)
);

OA22x2_ASAP7_75t_L g12949 ( 
.A1(n_12548),
.A2(n_1344),
.B1(n_1342),
.B2(n_1343),
.Y(n_12949)
);

AO31x2_ASAP7_75t_L g12950 ( 
.A1(n_12636),
.A2(n_1346),
.A3(n_1344),
.B(n_1345),
.Y(n_12950)
);

NAND2xp5_ASAP7_75t_L g12951 ( 
.A(n_12173),
.B(n_1345),
.Y(n_12951)
);

NAND2xp5_ASAP7_75t_L g12952 ( 
.A(n_12175),
.B(n_12201),
.Y(n_12952)
);

NAND2x1_ASAP7_75t_L g12953 ( 
.A(n_12014),
.B(n_1346),
.Y(n_12953)
);

A2O1A1Ixp33_ASAP7_75t_L g12954 ( 
.A1(n_11990),
.A2(n_1349),
.B(n_1347),
.C(n_1348),
.Y(n_12954)
);

NAND2xp5_ASAP7_75t_L g12955 ( 
.A(n_12220),
.B(n_1348),
.Y(n_12955)
);

AOI22xp33_ASAP7_75t_SL g12956 ( 
.A1(n_12247),
.A2(n_1351),
.B1(n_1349),
.B2(n_1350),
.Y(n_12956)
);

NAND2xp5_ASAP7_75t_L g12957 ( 
.A(n_12126),
.B(n_1350),
.Y(n_12957)
);

INVxp67_ASAP7_75t_L g12958 ( 
.A(n_12230),
.Y(n_12958)
);

NAND2xp5_ASAP7_75t_SL g12959 ( 
.A(n_12330),
.B(n_1351),
.Y(n_12959)
);

OR2x2_ASAP7_75t_L g12960 ( 
.A(n_12109),
.B(n_1352),
.Y(n_12960)
);

INVx3_ASAP7_75t_L g12961 ( 
.A(n_12143),
.Y(n_12961)
);

AO31x2_ASAP7_75t_L g12962 ( 
.A1(n_12658),
.A2(n_1355),
.A3(n_1352),
.B(n_1354),
.Y(n_12962)
);

AND2x2_ASAP7_75t_L g12963 ( 
.A(n_12452),
.B(n_1354),
.Y(n_12963)
);

AOI21xp5_ASAP7_75t_L g12964 ( 
.A1(n_11981),
.A2(n_1355),
.B(n_1357),
.Y(n_12964)
);

BUFx3_ASAP7_75t_L g12965 ( 
.A(n_12205),
.Y(n_12965)
);

NOR2xp33_ASAP7_75t_L g12966 ( 
.A(n_11875),
.B(n_1357),
.Y(n_12966)
);

BUFx2_ASAP7_75t_L g12967 ( 
.A(n_12185),
.Y(n_12967)
);

NAND2xp5_ASAP7_75t_L g12968 ( 
.A(n_12127),
.B(n_1358),
.Y(n_12968)
);

OAI21x1_ASAP7_75t_L g12969 ( 
.A1(n_11985),
.A2(n_1358),
.B(n_1359),
.Y(n_12969)
);

NOR2x1_ASAP7_75t_SL g12970 ( 
.A(n_11981),
.B(n_1359),
.Y(n_12970)
);

AO31x2_ASAP7_75t_L g12971 ( 
.A1(n_12661),
.A2(n_1362),
.A3(n_1360),
.B(n_1361),
.Y(n_12971)
);

NAND2xp5_ASAP7_75t_L g12972 ( 
.A(n_12134),
.B(n_1361),
.Y(n_12972)
);

NAND2xp5_ASAP7_75t_L g12973 ( 
.A(n_12165),
.B(n_12178),
.Y(n_12973)
);

AND2x6_ASAP7_75t_SL g12974 ( 
.A(n_11928),
.B(n_1362),
.Y(n_12974)
);

OAI21x1_ASAP7_75t_SL g12975 ( 
.A1(n_11781),
.A2(n_1363),
.B(n_1364),
.Y(n_12975)
);

OAI21xp5_ASAP7_75t_L g12976 ( 
.A1(n_12153),
.A2(n_1363),
.B(n_1364),
.Y(n_12976)
);

INVx1_ASAP7_75t_L g12977 ( 
.A(n_12063),
.Y(n_12977)
);

INVx2_ASAP7_75t_L g12978 ( 
.A(n_12532),
.Y(n_12978)
);

INVx2_ASAP7_75t_L g12979 ( 
.A(n_12539),
.Y(n_12979)
);

OAI22xp5_ASAP7_75t_L g12980 ( 
.A1(n_12563),
.A2(n_1367),
.B1(n_1365),
.B2(n_1366),
.Y(n_12980)
);

OAI21x1_ASAP7_75t_L g12981 ( 
.A1(n_12372),
.A2(n_1365),
.B(n_1366),
.Y(n_12981)
);

INVx3_ASAP7_75t_L g12982 ( 
.A(n_11915),
.Y(n_12982)
);

OAI21xp33_ASAP7_75t_L g12983 ( 
.A1(n_11853),
.A2(n_1368),
.B(n_1369),
.Y(n_12983)
);

NAND2xp5_ASAP7_75t_L g12984 ( 
.A(n_12191),
.B(n_1368),
.Y(n_12984)
);

AOI211x1_ASAP7_75t_L g12985 ( 
.A1(n_12188),
.A2(n_1372),
.B(n_1370),
.C(n_1371),
.Y(n_12985)
);

OAI21x1_ASAP7_75t_L g12986 ( 
.A1(n_12374),
.A2(n_1370),
.B(n_1371),
.Y(n_12986)
);

OAI21x1_ASAP7_75t_L g12987 ( 
.A1(n_12388),
.A2(n_1372),
.B(n_1373),
.Y(n_12987)
);

NAND2xp5_ASAP7_75t_L g12988 ( 
.A(n_12225),
.B(n_1373),
.Y(n_12988)
);

INVxp67_ASAP7_75t_SL g12989 ( 
.A(n_12544),
.Y(n_12989)
);

INVx1_ASAP7_75t_L g12990 ( 
.A(n_12083),
.Y(n_12990)
);

INVxp67_ASAP7_75t_SL g12991 ( 
.A(n_12581),
.Y(n_12991)
);

OAI21x1_ASAP7_75t_L g12992 ( 
.A1(n_12081),
.A2(n_1374),
.B(n_1375),
.Y(n_12992)
);

OAI21x1_ASAP7_75t_L g12993 ( 
.A1(n_12030),
.A2(n_1374),
.B(n_1375),
.Y(n_12993)
);

NOR2xp67_ASAP7_75t_SL g12994 ( 
.A(n_12020),
.B(n_1376),
.Y(n_12994)
);

BUFx4_ASAP7_75t_SL g12995 ( 
.A(n_12042),
.Y(n_12995)
);

NAND2xp5_ASAP7_75t_L g12996 ( 
.A(n_12252),
.B(n_1376),
.Y(n_12996)
);

INVx1_ASAP7_75t_L g12997 ( 
.A(n_12589),
.Y(n_12997)
);

OAI21x1_ASAP7_75t_L g12998 ( 
.A1(n_12486),
.A2(n_12157),
.B(n_12110),
.Y(n_12998)
);

NAND2xp5_ASAP7_75t_L g12999 ( 
.A(n_12256),
.B(n_1377),
.Y(n_12999)
);

NAND2xp5_ASAP7_75t_L g13000 ( 
.A(n_12261),
.B(n_1377),
.Y(n_13000)
);

OAI21x1_ASAP7_75t_L g13001 ( 
.A1(n_12096),
.A2(n_1378),
.B(n_1379),
.Y(n_13001)
);

AOI21x1_ASAP7_75t_L g13002 ( 
.A1(n_12226),
.A2(n_1378),
.B(n_1380),
.Y(n_13002)
);

OAI21x1_ASAP7_75t_SL g13003 ( 
.A1(n_11994),
.A2(n_1380),
.B(n_1381),
.Y(n_13003)
);

BUFx10_ASAP7_75t_L g13004 ( 
.A(n_11959),
.Y(n_13004)
);

NAND2xp5_ASAP7_75t_L g13005 ( 
.A(n_12265),
.B(n_1381),
.Y(n_13005)
);

A2O1A1Ixp33_ASAP7_75t_L g13006 ( 
.A1(n_11801),
.A2(n_1384),
.B(n_1382),
.C(n_1383),
.Y(n_13006)
);

NAND2xp5_ASAP7_75t_L g13007 ( 
.A(n_12283),
.B(n_1382),
.Y(n_13007)
);

OAI22xp5_ASAP7_75t_L g13008 ( 
.A1(n_12677),
.A2(n_1385),
.B1(n_1383),
.B2(n_1384),
.Y(n_13008)
);

AND2x2_ASAP7_75t_L g13009 ( 
.A(n_12141),
.B(n_1385),
.Y(n_13009)
);

OAI21x1_ASAP7_75t_L g13010 ( 
.A1(n_12473),
.A2(n_1386),
.B(n_1387),
.Y(n_13010)
);

OAI22xp5_ASAP7_75t_L g13011 ( 
.A1(n_12683),
.A2(n_1389),
.B1(n_1386),
.B2(n_1388),
.Y(n_13011)
);

BUFx4f_ASAP7_75t_SL g13012 ( 
.A(n_12049),
.Y(n_13012)
);

BUFx3_ASAP7_75t_L g13013 ( 
.A(n_12101),
.Y(n_13013)
);

OAI21x1_ASAP7_75t_SL g13014 ( 
.A1(n_12019),
.A2(n_1388),
.B(n_1389),
.Y(n_13014)
);

BUFx10_ASAP7_75t_L g13015 ( 
.A(n_12562),
.Y(n_13015)
);

OAI21x1_ASAP7_75t_L g13016 ( 
.A1(n_12409),
.A2(n_1390),
.B(n_1391),
.Y(n_13016)
);

BUFx2_ASAP7_75t_L g13017 ( 
.A(n_12219),
.Y(n_13017)
);

AO31x2_ASAP7_75t_L g13018 ( 
.A1(n_12675),
.A2(n_1392),
.A3(n_1390),
.B(n_1391),
.Y(n_13018)
);

AND2x2_ASAP7_75t_L g13019 ( 
.A(n_12384),
.B(n_1392),
.Y(n_13019)
);

AOI21xp5_ASAP7_75t_L g13020 ( 
.A1(n_12466),
.A2(n_1393),
.B(n_1394),
.Y(n_13020)
);

OAI21x1_ASAP7_75t_L g13021 ( 
.A1(n_12413),
.A2(n_1393),
.B(n_1394),
.Y(n_13021)
);

OA22x2_ASAP7_75t_L g13022 ( 
.A1(n_12548),
.A2(n_1397),
.B1(n_1395),
.B2(n_1396),
.Y(n_13022)
);

OAI21xp5_ASAP7_75t_L g13023 ( 
.A1(n_11999),
.A2(n_1395),
.B(n_1397),
.Y(n_13023)
);

INVx4_ASAP7_75t_L g13024 ( 
.A(n_12091),
.Y(n_13024)
);

NAND2xp5_ASAP7_75t_L g13025 ( 
.A(n_12301),
.B(n_1398),
.Y(n_13025)
);

OAI21x1_ASAP7_75t_L g13026 ( 
.A1(n_12432),
.A2(n_12440),
.B(n_12435),
.Y(n_13026)
);

OAI21xp5_ASAP7_75t_L g13027 ( 
.A1(n_12038),
.A2(n_12052),
.B(n_12216),
.Y(n_13027)
);

O2A1O1Ixp5_ASAP7_75t_L g13028 ( 
.A1(n_11882),
.A2(n_1400),
.B(n_1398),
.C(n_1399),
.Y(n_13028)
);

INVx1_ASAP7_75t_L g13029 ( 
.A(n_12594),
.Y(n_13029)
);

OAI21x1_ASAP7_75t_L g13030 ( 
.A1(n_12463),
.A2(n_1399),
.B(n_1401),
.Y(n_13030)
);

INVx1_ASAP7_75t_L g13031 ( 
.A(n_12595),
.Y(n_13031)
);

AOI21xp5_ASAP7_75t_L g13032 ( 
.A1(n_12085),
.A2(n_1401),
.B(n_1402),
.Y(n_13032)
);

A2O1A1Ixp33_ASAP7_75t_L g13033 ( 
.A1(n_11845),
.A2(n_1404),
.B(n_1402),
.C(n_1403),
.Y(n_13033)
);

NAND2xp5_ASAP7_75t_L g13034 ( 
.A(n_12118),
.B(n_1403),
.Y(n_13034)
);

OAI21xp5_ASAP7_75t_L g13035 ( 
.A1(n_12160),
.A2(n_1404),
.B(n_1405),
.Y(n_13035)
);

NAND2xp5_ASAP7_75t_L g13036 ( 
.A(n_12120),
.B(n_1405),
.Y(n_13036)
);

NAND2xp5_ASAP7_75t_L g13037 ( 
.A(n_12122),
.B(n_1406),
.Y(n_13037)
);

AOI21xp5_ASAP7_75t_L g13038 ( 
.A1(n_11834),
.A2(n_1406),
.B(n_1407),
.Y(n_13038)
);

NAND2xp5_ASAP7_75t_L g13039 ( 
.A(n_12125),
.B(n_1408),
.Y(n_13039)
);

INVx1_ASAP7_75t_L g13040 ( 
.A(n_12604),
.Y(n_13040)
);

INVx2_ASAP7_75t_L g13041 ( 
.A(n_12624),
.Y(n_13041)
);

AOI21xp5_ASAP7_75t_L g13042 ( 
.A1(n_12501),
.A2(n_1408),
.B(n_1409),
.Y(n_13042)
);

AOI22xp5_ASAP7_75t_L g13043 ( 
.A1(n_11856),
.A2(n_1411),
.B1(n_1409),
.B2(n_1410),
.Y(n_13043)
);

NAND2xp5_ASAP7_75t_L g13044 ( 
.A(n_12150),
.B(n_1410),
.Y(n_13044)
);

AND2x4_ASAP7_75t_L g13045 ( 
.A(n_12640),
.B(n_1411),
.Y(n_13045)
);

OAI21xp5_ASAP7_75t_L g13046 ( 
.A1(n_12161),
.A2(n_1412),
.B(n_1413),
.Y(n_13046)
);

NOR2xp33_ASAP7_75t_L g13047 ( 
.A(n_12176),
.B(n_1412),
.Y(n_13047)
);

INVx1_ASAP7_75t_SL g13048 ( 
.A(n_11949),
.Y(n_13048)
);

NAND2x1p5_ASAP7_75t_L g13049 ( 
.A(n_12249),
.B(n_1413),
.Y(n_13049)
);

OR2x2_ASAP7_75t_L g13050 ( 
.A(n_12387),
.B(n_1414),
.Y(n_13050)
);

A2O1A1Ixp33_ASAP7_75t_L g13051 ( 
.A1(n_11892),
.A2(n_1416),
.B(n_1414),
.C(n_1415),
.Y(n_13051)
);

AND2x2_ASAP7_75t_L g13052 ( 
.A(n_12384),
.B(n_1415),
.Y(n_13052)
);

OAI21x1_ASAP7_75t_L g13053 ( 
.A1(n_12402),
.A2(n_1416),
.B(n_1417),
.Y(n_13053)
);

NAND2xp5_ASAP7_75t_L g13054 ( 
.A(n_12277),
.B(n_1417),
.Y(n_13054)
);

NAND2xp5_ASAP7_75t_L g13055 ( 
.A(n_12279),
.B(n_1418),
.Y(n_13055)
);

AND2x2_ASAP7_75t_L g13056 ( 
.A(n_12410),
.B(n_1418),
.Y(n_13056)
);

NOR2xp33_ASAP7_75t_L g13057 ( 
.A(n_12342),
.B(n_1419),
.Y(n_13057)
);

OAI21xp5_ASAP7_75t_L g13058 ( 
.A1(n_12123),
.A2(n_1419),
.B(n_1420),
.Y(n_13058)
);

OAI21xp5_ASAP7_75t_L g13059 ( 
.A1(n_12232),
.A2(n_1420),
.B(n_1421),
.Y(n_13059)
);

AOI21x1_ASAP7_75t_L g13060 ( 
.A1(n_11967),
.A2(n_12320),
.B(n_11938),
.Y(n_13060)
);

OAI21x1_ASAP7_75t_L g13061 ( 
.A1(n_12117),
.A2(n_1422),
.B(n_1423),
.Y(n_13061)
);

INVx3_ASAP7_75t_L g13062 ( 
.A(n_11963),
.Y(n_13062)
);

AND2x2_ASAP7_75t_L g13063 ( 
.A(n_12410),
.B(n_1422),
.Y(n_13063)
);

OR2x2_ASAP7_75t_L g13064 ( 
.A(n_12451),
.B(n_1423),
.Y(n_13064)
);

NAND2xp5_ASAP7_75t_L g13065 ( 
.A(n_12287),
.B(n_1424),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_12665),
.Y(n_13066)
);

OAI21x1_ASAP7_75t_L g13067 ( 
.A1(n_12270),
.A2(n_1424),
.B(n_1425),
.Y(n_13067)
);

NOR2xp67_ASAP7_75t_L g13068 ( 
.A(n_12503),
.B(n_1425),
.Y(n_13068)
);

OAI21xp33_ASAP7_75t_L g13069 ( 
.A1(n_12617),
.A2(n_1426),
.B(n_1427),
.Y(n_13069)
);

NAND2xp5_ASAP7_75t_L g13070 ( 
.A(n_12291),
.B(n_1426),
.Y(n_13070)
);

NAND2xp5_ASAP7_75t_SL g13071 ( 
.A(n_12329),
.B(n_1428),
.Y(n_13071)
);

AO31x2_ASAP7_75t_L g13072 ( 
.A1(n_12154),
.A2(n_1431),
.A3(n_1429),
.B(n_1430),
.Y(n_13072)
);

OAI22x1_ASAP7_75t_L g13073 ( 
.A1(n_11982),
.A2(n_1432),
.B1(n_1430),
.B2(n_1431),
.Y(n_13073)
);

OAI21xp5_ASAP7_75t_L g13074 ( 
.A1(n_12235),
.A2(n_1432),
.B(n_1433),
.Y(n_13074)
);

A2O1A1Ixp33_ASAP7_75t_L g13075 ( 
.A1(n_11905),
.A2(n_1435),
.B(n_1433),
.C(n_1434),
.Y(n_13075)
);

AND2x2_ASAP7_75t_L g13076 ( 
.A(n_12379),
.B(n_1434),
.Y(n_13076)
);

NAND2xp5_ASAP7_75t_L g13077 ( 
.A(n_12299),
.B(n_1435),
.Y(n_13077)
);

INVx1_ASAP7_75t_L g13078 ( 
.A(n_12015),
.Y(n_13078)
);

OAI21x1_ASAP7_75t_L g13079 ( 
.A1(n_12274),
.A2(n_1436),
.B(n_1437),
.Y(n_13079)
);

OAI21xp5_ASAP7_75t_L g13080 ( 
.A1(n_12470),
.A2(n_1436),
.B(n_1437),
.Y(n_13080)
);

OAI21x1_ASAP7_75t_L g13081 ( 
.A1(n_12278),
.A2(n_1438),
.B(n_1439),
.Y(n_13081)
);

OAI21x1_ASAP7_75t_L g13082 ( 
.A1(n_12298),
.A2(n_1438),
.B(n_1439),
.Y(n_13082)
);

BUFx2_ASAP7_75t_L g13083 ( 
.A(n_12156),
.Y(n_13083)
);

NAND2xp5_ASAP7_75t_L g13084 ( 
.A(n_12392),
.B(n_1440),
.Y(n_13084)
);

CKINVDCx20_ASAP7_75t_R g13085 ( 
.A(n_12531),
.Y(n_13085)
);

NAND2x1p5_ASAP7_75t_L g13086 ( 
.A(n_12319),
.B(n_1440),
.Y(n_13086)
);

BUFx6f_ASAP7_75t_L g13087 ( 
.A(n_12187),
.Y(n_13087)
);

INVx3_ASAP7_75t_L g13088 ( 
.A(n_12058),
.Y(n_13088)
);

OAI21x1_ASAP7_75t_L g13089 ( 
.A1(n_12302),
.A2(n_1441),
.B(n_1442),
.Y(n_13089)
);

NAND2xp5_ASAP7_75t_L g13090 ( 
.A(n_12241),
.B(n_1441),
.Y(n_13090)
);

OAI21x1_ASAP7_75t_L g13091 ( 
.A1(n_12304),
.A2(n_1443),
.B(n_1444),
.Y(n_13091)
);

NOR2xp33_ASAP7_75t_L g13092 ( 
.A(n_11753),
.B(n_12507),
.Y(n_13092)
);

NAND2xp5_ASAP7_75t_L g13093 ( 
.A(n_12428),
.B(n_12312),
.Y(n_13093)
);

AOI22xp5_ASAP7_75t_L g13094 ( 
.A1(n_11870),
.A2(n_1446),
.B1(n_1443),
.B2(n_1445),
.Y(n_13094)
);

AOI21xp5_ASAP7_75t_L g13095 ( 
.A1(n_12510),
.A2(n_1445),
.B(n_1446),
.Y(n_13095)
);

AOI21xp5_ASAP7_75t_L g13096 ( 
.A1(n_12512),
.A2(n_1447),
.B(n_1448),
.Y(n_13096)
);

AOI21xp5_ASAP7_75t_L g13097 ( 
.A1(n_12518),
.A2(n_1449),
.B(n_1450),
.Y(n_13097)
);

OR2x6_ASAP7_75t_L g13098 ( 
.A(n_12254),
.B(n_1449),
.Y(n_13098)
);

OAI21x1_ASAP7_75t_L g13099 ( 
.A1(n_12318),
.A2(n_1450),
.B(n_1451),
.Y(n_13099)
);

NAND2xp5_ASAP7_75t_SL g13100 ( 
.A(n_12482),
.B(n_1452),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_12034),
.Y(n_13101)
);

NAND2x1_ASAP7_75t_L g13102 ( 
.A(n_12054),
.B(n_1452),
.Y(n_13102)
);

OAI22xp5_ASAP7_75t_L g13103 ( 
.A1(n_12212),
.A2(n_1455),
.B1(n_1453),
.B2(n_1454),
.Y(n_13103)
);

NAND2x1p5_ASAP7_75t_L g13104 ( 
.A(n_12491),
.B(n_1453),
.Y(n_13104)
);

NAND2xp5_ASAP7_75t_L g13105 ( 
.A(n_12310),
.B(n_1456),
.Y(n_13105)
);

AOI21xp5_ASAP7_75t_L g13106 ( 
.A1(n_12536),
.A2(n_12577),
.B(n_12543),
.Y(n_13106)
);

INVx4_ASAP7_75t_L g13107 ( 
.A(n_12069),
.Y(n_13107)
);

AND2x4_ASAP7_75t_L g13108 ( 
.A(n_12106),
.B(n_12057),
.Y(n_13108)
);

AOI21xp5_ASAP7_75t_L g13109 ( 
.A1(n_12593),
.A2(n_1456),
.B(n_1457),
.Y(n_13109)
);

OAI21xp5_ASAP7_75t_L g13110 ( 
.A1(n_12328),
.A2(n_1457),
.B(n_1458),
.Y(n_13110)
);

INVx2_ASAP7_75t_L g13111 ( 
.A(n_12060),
.Y(n_13111)
);

NAND2x1p5_ASAP7_75t_L g13112 ( 
.A(n_12503),
.B(n_1458),
.Y(n_13112)
);

INVx4_ASAP7_75t_L g13113 ( 
.A(n_12187),
.Y(n_13113)
);

INVx1_ASAP7_75t_L g13114 ( 
.A(n_12073),
.Y(n_13114)
);

AO21x2_ASAP7_75t_L g13115 ( 
.A1(n_11806),
.A2(n_1459),
.B(n_1460),
.Y(n_13115)
);

NAND2xp5_ASAP7_75t_L g13116 ( 
.A(n_12045),
.B(n_1459),
.Y(n_13116)
);

INVx2_ASAP7_75t_L g13117 ( 
.A(n_12082),
.Y(n_13117)
);

OAI21xp5_ASAP7_75t_L g13118 ( 
.A1(n_12029),
.A2(n_1461),
.B(n_1462),
.Y(n_13118)
);

OAI21xp5_ASAP7_75t_L g13119 ( 
.A1(n_12361),
.A2(n_1461),
.B(n_1462),
.Y(n_13119)
);

OAI21x1_ASAP7_75t_L g13120 ( 
.A1(n_12259),
.A2(n_1463),
.B(n_1464),
.Y(n_13120)
);

OAI21x1_ASAP7_75t_L g13121 ( 
.A1(n_12111),
.A2(n_1463),
.B(n_1464),
.Y(n_13121)
);

NAND2xp5_ASAP7_75t_L g13122 ( 
.A(n_12431),
.B(n_1465),
.Y(n_13122)
);

NOR2xp33_ASAP7_75t_SL g13123 ( 
.A(n_12152),
.B(n_1465),
.Y(n_13123)
);

AO21x1_ASAP7_75t_L g13124 ( 
.A1(n_12357),
.A2(n_1466),
.B(n_1467),
.Y(n_13124)
);

NAND2xp5_ASAP7_75t_L g13125 ( 
.A(n_12441),
.B(n_1466),
.Y(n_13125)
);

INVx8_ASAP7_75t_L g13126 ( 
.A(n_11763),
.Y(n_13126)
);

AOI22xp5_ASAP7_75t_L g13127 ( 
.A1(n_12023),
.A2(n_1469),
.B1(n_1467),
.B2(n_1468),
.Y(n_13127)
);

BUFx2_ASAP7_75t_SL g13128 ( 
.A(n_12180),
.Y(n_13128)
);

BUFx2_ASAP7_75t_L g13129 ( 
.A(n_12206),
.Y(n_13129)
);

BUFx2_ASAP7_75t_L g13130 ( 
.A(n_12311),
.Y(n_13130)
);

OAI21x1_ASAP7_75t_L g13131 ( 
.A1(n_12484),
.A2(n_1468),
.B(n_1469),
.Y(n_13131)
);

OAI21xp5_ASAP7_75t_L g13132 ( 
.A1(n_11858),
.A2(n_1470),
.B(n_1471),
.Y(n_13132)
);

AOI21x1_ASAP7_75t_L g13133 ( 
.A1(n_12600),
.A2(n_1471),
.B(n_1472),
.Y(n_13133)
);

NAND2xp5_ASAP7_75t_L g13134 ( 
.A(n_12443),
.B(n_1473),
.Y(n_13134)
);

AOI21xp5_ASAP7_75t_L g13135 ( 
.A1(n_12606),
.A2(n_1473),
.B(n_1474),
.Y(n_13135)
);

OAI21xp5_ASAP7_75t_SL g13136 ( 
.A1(n_11921),
.A2(n_1474),
.B(n_1475),
.Y(n_13136)
);

OAI21x1_ASAP7_75t_L g13137 ( 
.A1(n_12499),
.A2(n_1476),
.B(n_1477),
.Y(n_13137)
);

OAI21x1_ASAP7_75t_SL g13138 ( 
.A1(n_11926),
.A2(n_1477),
.B(n_1479),
.Y(n_13138)
);

A2O1A1Ixp33_ASAP7_75t_L g13139 ( 
.A1(n_12010),
.A2(n_1482),
.B(n_1480),
.C(n_1481),
.Y(n_13139)
);

AOI21xp33_ASAP7_75t_L g13140 ( 
.A1(n_12033),
.A2(n_1480),
.B(n_1482),
.Y(n_13140)
);

INVx5_ASAP7_75t_L g13141 ( 
.A(n_11763),
.Y(n_13141)
);

AOI22xp33_ASAP7_75t_L g13142 ( 
.A1(n_12684),
.A2(n_1485),
.B1(n_1483),
.B2(n_1484),
.Y(n_13142)
);

AND2x2_ASAP7_75t_L g13143 ( 
.A(n_12379),
.B(n_1483),
.Y(n_13143)
);

OAI21x1_ASAP7_75t_L g13144 ( 
.A1(n_12616),
.A2(n_1485),
.B(n_1486),
.Y(n_13144)
);

OAI21x1_ASAP7_75t_L g13145 ( 
.A1(n_12623),
.A2(n_1486),
.B(n_1487),
.Y(n_13145)
);

INVx1_ASAP7_75t_L g13146 ( 
.A(n_11816),
.Y(n_13146)
);

NAND2xp5_ASAP7_75t_SL g13147 ( 
.A(n_12482),
.B(n_1487),
.Y(n_13147)
);

NAND2xp5_ASAP7_75t_L g13148 ( 
.A(n_12444),
.B(n_1488),
.Y(n_13148)
);

INVx4_ASAP7_75t_L g13149 ( 
.A(n_12190),
.Y(n_13149)
);

NAND2xp5_ASAP7_75t_L g13150 ( 
.A(n_12412),
.B(n_1488),
.Y(n_13150)
);

INVx1_ASAP7_75t_L g13151 ( 
.A(n_11847),
.Y(n_13151)
);

OAI21xp5_ASAP7_75t_L g13152 ( 
.A1(n_11861),
.A2(n_1489),
.B(n_1490),
.Y(n_13152)
);

A2O1A1Ixp33_ASAP7_75t_L g13153 ( 
.A1(n_12128),
.A2(n_1491),
.B(n_1489),
.C(n_1490),
.Y(n_13153)
);

OA21x2_ASAP7_75t_L g13154 ( 
.A1(n_12135),
.A2(n_1491),
.B(n_1492),
.Y(n_13154)
);

OAI21xp5_ASAP7_75t_L g13155 ( 
.A1(n_11867),
.A2(n_1492),
.B(n_1493),
.Y(n_13155)
);

INVx2_ASAP7_75t_L g13156 ( 
.A(n_12005),
.Y(n_13156)
);

AOI21xp5_ASAP7_75t_L g13157 ( 
.A1(n_12653),
.A2(n_1493),
.B(n_1494),
.Y(n_13157)
);

NAND2xp5_ASAP7_75t_L g13158 ( 
.A(n_12414),
.B(n_1495),
.Y(n_13158)
);

OAI21x1_ASAP7_75t_L g13159 ( 
.A1(n_12687),
.A2(n_1495),
.B(n_1496),
.Y(n_13159)
);

OAI21xp5_ASAP7_75t_L g13160 ( 
.A1(n_11888),
.A2(n_12046),
.B(n_12464),
.Y(n_13160)
);

AOI22xp5_ASAP7_75t_L g13161 ( 
.A1(n_12303),
.A2(n_1498),
.B1(n_1496),
.B2(n_1497),
.Y(n_13161)
);

AOI22x1_ASAP7_75t_L g13162 ( 
.A1(n_12094),
.A2(n_1502),
.B1(n_1499),
.B2(n_1501),
.Y(n_13162)
);

AOI22xp5_ASAP7_75t_L g13163 ( 
.A1(n_12237),
.A2(n_1502),
.B1(n_1499),
.B2(n_1501),
.Y(n_13163)
);

OAI21x1_ASAP7_75t_SL g13164 ( 
.A1(n_12159),
.A2(n_1503),
.B(n_1504),
.Y(n_13164)
);

OAI22xp5_ASAP7_75t_L g13165 ( 
.A1(n_12105),
.A2(n_1505),
.B1(n_1503),
.B2(n_1504),
.Y(n_13165)
);

NOR2xp67_ASAP7_75t_SL g13166 ( 
.A(n_11997),
.B(n_1505),
.Y(n_13166)
);

AOI21xp5_ASAP7_75t_L g13167 ( 
.A1(n_12214),
.A2(n_1506),
.B(n_1507),
.Y(n_13167)
);

NAND2xp5_ASAP7_75t_L g13168 ( 
.A(n_12031),
.B(n_1506),
.Y(n_13168)
);

INVx1_ASAP7_75t_SL g13169 ( 
.A(n_12107),
.Y(n_13169)
);

OA21x2_ASAP7_75t_L g13170 ( 
.A1(n_12174),
.A2(n_1507),
.B(n_1508),
.Y(n_13170)
);

OAI21x1_ASAP7_75t_L g13171 ( 
.A1(n_11933),
.A2(n_1508),
.B(n_1509),
.Y(n_13171)
);

AOI21x1_ASAP7_75t_L g13172 ( 
.A1(n_11869),
.A2(n_1509),
.B(n_1510),
.Y(n_13172)
);

INVxp67_ASAP7_75t_SL g13173 ( 
.A(n_12455),
.Y(n_13173)
);

OAI21xp5_ASAP7_75t_L g13174 ( 
.A1(n_12461),
.A2(n_1510),
.B(n_1511),
.Y(n_13174)
);

NAND2xp5_ASAP7_75t_L g13175 ( 
.A(n_12041),
.B(n_1511),
.Y(n_13175)
);

OA21x2_ASAP7_75t_L g13176 ( 
.A1(n_12196),
.A2(n_11988),
.B(n_11804),
.Y(n_13176)
);

OAI21xp5_ASAP7_75t_L g13177 ( 
.A1(n_12004),
.A2(n_1512),
.B(n_1513),
.Y(n_13177)
);

BUFx5_ASAP7_75t_L g13178 ( 
.A(n_12460),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_11976),
.Y(n_13179)
);

AOI21xp5_ASAP7_75t_SL g13180 ( 
.A1(n_12237),
.A2(n_1513),
.B(n_1515),
.Y(n_13180)
);

OAI21x1_ASAP7_75t_L g13181 ( 
.A1(n_12457),
.A2(n_1515),
.B(n_1516),
.Y(n_13181)
);

NAND2xp5_ASAP7_75t_SL g13182 ( 
.A(n_12438),
.B(n_1517),
.Y(n_13182)
);

OA22x2_ASAP7_75t_L g13183 ( 
.A1(n_11898),
.A2(n_12001),
.B1(n_11929),
.B2(n_11932),
.Y(n_13183)
);

NAND3x1_ASAP7_75t_L g13184 ( 
.A(n_12282),
.B(n_1517),
.C(n_1519),
.Y(n_13184)
);

OA21x2_ASAP7_75t_L g13185 ( 
.A1(n_11775),
.A2(n_1519),
.B(n_1520),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_12317),
.B(n_1520),
.Y(n_13186)
);

NAND2xp5_ASAP7_75t_L g13187 ( 
.A(n_11758),
.B(n_1521),
.Y(n_13187)
);

AO21x1_ASAP7_75t_L g13188 ( 
.A1(n_12009),
.A2(n_1521),
.B(n_1522),
.Y(n_13188)
);

INVx2_ASAP7_75t_L g13189 ( 
.A(n_11773),
.Y(n_13189)
);

NAND2xp5_ASAP7_75t_L g13190 ( 
.A(n_12504),
.B(n_1522),
.Y(n_13190)
);

INVxp67_ASAP7_75t_L g13191 ( 
.A(n_12434),
.Y(n_13191)
);

A2O1A1Ixp33_ASAP7_75t_L g13192 ( 
.A1(n_12248),
.A2(n_12257),
.B(n_12344),
.C(n_12481),
.Y(n_13192)
);

AOI21xp5_ASAP7_75t_L g13193 ( 
.A1(n_12215),
.A2(n_1523),
.B(n_1524),
.Y(n_13193)
);

AOI21xp33_ASAP7_75t_L g13194 ( 
.A1(n_12467),
.A2(n_1523),
.B(n_1525),
.Y(n_13194)
);

A2O1A1Ixp33_ASAP7_75t_L g13195 ( 
.A1(n_12211),
.A2(n_1528),
.B(n_1526),
.C(n_1527),
.Y(n_13195)
);

CKINVDCx5p33_ASAP7_75t_R g13196 ( 
.A(n_12612),
.Y(n_13196)
);

AOI21xp5_ASAP7_75t_L g13197 ( 
.A1(n_12326),
.A2(n_1527),
.B(n_1528),
.Y(n_13197)
);

OAI21xp5_ASAP7_75t_L g13198 ( 
.A1(n_12168),
.A2(n_1529),
.B(n_1530),
.Y(n_13198)
);

INVx1_ASAP7_75t_L g13199 ( 
.A(n_12685),
.Y(n_13199)
);

O2A1O1Ixp5_ASAP7_75t_L g13200 ( 
.A1(n_12144),
.A2(n_1531),
.B(n_1529),
.C(n_1530),
.Y(n_13200)
);

NAND2x1_ASAP7_75t_L g13201 ( 
.A(n_12445),
.B(n_1531),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_11780),
.Y(n_13202)
);

NAND2xp5_ASAP7_75t_SL g13203 ( 
.A(n_12514),
.B(n_1532),
.Y(n_13203)
);

BUFx2_ASAP7_75t_L g13204 ( 
.A(n_12254),
.Y(n_13204)
);

NAND2xp5_ASAP7_75t_SL g13205 ( 
.A(n_12514),
.B(n_1532),
.Y(n_13205)
);

NAND2xp5_ASAP7_75t_L g13206 ( 
.A(n_12523),
.B(n_1533),
.Y(n_13206)
);

OAI21x1_ASAP7_75t_L g13207 ( 
.A1(n_12246),
.A2(n_1533),
.B(n_1534),
.Y(n_13207)
);

INVxp67_ASAP7_75t_L g13208 ( 
.A(n_12434),
.Y(n_13208)
);

AOI21xp5_ASAP7_75t_L g13209 ( 
.A1(n_12390),
.A2(n_1534),
.B(n_1535),
.Y(n_13209)
);

CKINVDCx5p33_ASAP7_75t_R g13210 ( 
.A(n_12644),
.Y(n_13210)
);

AND2x2_ASAP7_75t_L g13211 ( 
.A(n_12448),
.B(n_1535),
.Y(n_13211)
);

AOI21xp5_ASAP7_75t_L g13212 ( 
.A1(n_12407),
.A2(n_1536),
.B(n_1537),
.Y(n_13212)
);

AO32x2_ASAP7_75t_L g13213 ( 
.A1(n_11987),
.A2(n_11821),
.A3(n_12525),
.B1(n_12522),
.B2(n_11854),
.Y(n_13213)
);

NAND2xp5_ASAP7_75t_L g13214 ( 
.A(n_12524),
.B(n_1537),
.Y(n_13214)
);

NOR2xp33_ASAP7_75t_L g13215 ( 
.A(n_12508),
.B(n_1538),
.Y(n_13215)
);

OAI21x1_ASAP7_75t_L g13216 ( 
.A1(n_12391),
.A2(n_1538),
.B(n_1539),
.Y(n_13216)
);

NAND2xp5_ASAP7_75t_L g13217 ( 
.A(n_12559),
.B(n_1539),
.Y(n_13217)
);

INVx1_ASAP7_75t_L g13218 ( 
.A(n_11992),
.Y(n_13218)
);

OAI22xp5_ASAP7_75t_L g13219 ( 
.A1(n_12028),
.A2(n_12258),
.B1(n_12602),
.B2(n_12363),
.Y(n_13219)
);

OAI21x1_ASAP7_75t_L g13220 ( 
.A1(n_12458),
.A2(n_1540),
.B(n_1541),
.Y(n_13220)
);

OAI21xp5_ASAP7_75t_L g13221 ( 
.A1(n_12171),
.A2(n_1540),
.B(n_1541),
.Y(n_13221)
);

AOI21xp5_ASAP7_75t_L g13222 ( 
.A1(n_11848),
.A2(n_1542),
.B(n_1543),
.Y(n_13222)
);

NAND2xp5_ASAP7_75t_L g13223 ( 
.A(n_12567),
.B(n_1542),
.Y(n_13223)
);

OAI21x1_ASAP7_75t_L g13224 ( 
.A1(n_12163),
.A2(n_1544),
.B(n_1545),
.Y(n_13224)
);

AND2x4_ASAP7_75t_L g13225 ( 
.A(n_11900),
.B(n_1544),
.Y(n_13225)
);

OAI21x1_ASAP7_75t_L g13226 ( 
.A1(n_12167),
.A2(n_1545),
.B(n_1547),
.Y(n_13226)
);

OAI21xp5_ASAP7_75t_L g13227 ( 
.A1(n_12193),
.A2(n_1548),
.B(n_1549),
.Y(n_13227)
);

NAND2xp5_ASAP7_75t_L g13228 ( 
.A(n_12582),
.B(n_1548),
.Y(n_13228)
);

OAI21x1_ASAP7_75t_L g13229 ( 
.A1(n_12207),
.A2(n_1549),
.B(n_1550),
.Y(n_13229)
);

OAI21x1_ASAP7_75t_L g13230 ( 
.A1(n_12162),
.A2(n_1551),
.B(n_1553),
.Y(n_13230)
);

OAI21x1_ASAP7_75t_L g13231 ( 
.A1(n_12476),
.A2(n_1551),
.B(n_1553),
.Y(n_13231)
);

OAI21x1_ASAP7_75t_L g13232 ( 
.A1(n_12480),
.A2(n_1554),
.B(n_1555),
.Y(n_13232)
);

NAND2xp5_ASAP7_75t_L g13233 ( 
.A(n_12587),
.B(n_1554),
.Y(n_13233)
);

CKINVDCx11_ASAP7_75t_R g13234 ( 
.A(n_11896),
.Y(n_13234)
);

AND2x2_ASAP7_75t_L g13235 ( 
.A(n_12448),
.B(n_1555),
.Y(n_13235)
);

OAI21x1_ASAP7_75t_L g13236 ( 
.A1(n_12490),
.A2(n_1556),
.B(n_1557),
.Y(n_13236)
);

NAND2xp5_ASAP7_75t_L g13237 ( 
.A(n_12592),
.B(n_1556),
.Y(n_13237)
);

BUFx8_ASAP7_75t_L g13238 ( 
.A(n_12155),
.Y(n_13238)
);

NAND2xp5_ASAP7_75t_L g13239 ( 
.A(n_12597),
.B(n_12598),
.Y(n_13239)
);

NAND2xp5_ASAP7_75t_L g13240 ( 
.A(n_12609),
.B(n_1557),
.Y(n_13240)
);

AOI21xp5_ASAP7_75t_L g13241 ( 
.A1(n_12607),
.A2(n_1558),
.B(n_1559),
.Y(n_13241)
);

NAND2xp5_ASAP7_75t_SL g13242 ( 
.A(n_12528),
.B(n_1558),
.Y(n_13242)
);

AOI21xp5_ASAP7_75t_L g13243 ( 
.A1(n_12295),
.A2(n_1559),
.B(n_1560),
.Y(n_13243)
);

INVx2_ASAP7_75t_SL g13244 ( 
.A(n_12190),
.Y(n_13244)
);

A2O1A1Ixp33_ASAP7_75t_L g13245 ( 
.A1(n_12498),
.A2(n_1563),
.B(n_1561),
.C(n_1562),
.Y(n_13245)
);

NAND2xp5_ASAP7_75t_L g13246 ( 
.A(n_12613),
.B(n_1562),
.Y(n_13246)
);

NAND2xp5_ASAP7_75t_L g13247 ( 
.A(n_12626),
.B(n_12634),
.Y(n_13247)
);

BUFx2_ASAP7_75t_L g13248 ( 
.A(n_12224),
.Y(n_13248)
);

INVxp67_ASAP7_75t_SL g13249 ( 
.A(n_12228),
.Y(n_13249)
);

AND2x4_ASAP7_75t_L g13250 ( 
.A(n_12166),
.B(n_12528),
.Y(n_13250)
);

INVxp67_ASAP7_75t_SL g13251 ( 
.A(n_12007),
.Y(n_13251)
);

NAND2xp5_ASAP7_75t_SL g13252 ( 
.A(n_12347),
.B(n_1564),
.Y(n_13252)
);

OAI21xp5_ASAP7_75t_L g13253 ( 
.A1(n_12198),
.A2(n_12336),
.B(n_12488),
.Y(n_13253)
);

INVx1_ASAP7_75t_L g13254 ( 
.A(n_12012),
.Y(n_13254)
);

INVx2_ASAP7_75t_SL g13255 ( 
.A(n_12195),
.Y(n_13255)
);

AOI21xp5_ASAP7_75t_L g13256 ( 
.A1(n_12546),
.A2(n_1564),
.B(n_1565),
.Y(n_13256)
);

NAND2xp5_ASAP7_75t_L g13257 ( 
.A(n_12638),
.B(n_1565),
.Y(n_13257)
);

OAI21x1_ASAP7_75t_L g13258 ( 
.A1(n_12496),
.A2(n_1566),
.B(n_1567),
.Y(n_13258)
);

INVx4_ASAP7_75t_L g13259 ( 
.A(n_12195),
.Y(n_13259)
);

OAI21x1_ASAP7_75t_SL g13260 ( 
.A1(n_12420),
.A2(n_1568),
.B(n_1569),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_11838),
.Y(n_13261)
);

CKINVDCx5p33_ASAP7_75t_R g13262 ( 
.A(n_11901),
.Y(n_13262)
);

AOI22xp33_ASAP7_75t_L g13263 ( 
.A1(n_12393),
.A2(n_1572),
.B1(n_1568),
.B2(n_1570),
.Y(n_13263)
);

INVx1_ASAP7_75t_L g13264 ( 
.A(n_12022),
.Y(n_13264)
);

AOI21x1_ASAP7_75t_SL g13265 ( 
.A1(n_12148),
.A2(n_1570),
.B(n_1572),
.Y(n_13265)
);

NAND2x1_ASAP7_75t_L g13266 ( 
.A(n_11898),
.B(n_1573),
.Y(n_13266)
);

AND2x2_ASAP7_75t_L g13267 ( 
.A(n_12347),
.B(n_1573),
.Y(n_13267)
);

AOI21xp5_ASAP7_75t_L g13268 ( 
.A1(n_12557),
.A2(n_1574),
.B(n_1575),
.Y(n_13268)
);

OAI21x1_ASAP7_75t_L g13269 ( 
.A1(n_12032),
.A2(n_1574),
.B(n_1576),
.Y(n_13269)
);

BUFx2_ASAP7_75t_L g13270 ( 
.A(n_12158),
.Y(n_13270)
);

AOI21xp5_ASAP7_75t_L g13271 ( 
.A1(n_12568),
.A2(n_1576),
.B(n_1577),
.Y(n_13271)
);

AND2x4_ASAP7_75t_L g13272 ( 
.A(n_12199),
.B(n_1577),
.Y(n_13272)
);

INVx2_ASAP7_75t_SL g13273 ( 
.A(n_12202),
.Y(n_13273)
);

AOI22xp5_ASAP7_75t_L g13274 ( 
.A1(n_11930),
.A2(n_1580),
.B1(n_1578),
.B2(n_1579),
.Y(n_13274)
);

AOI221xp5_ASAP7_75t_L g13275 ( 
.A1(n_12397),
.A2(n_1580),
.B1(n_1578),
.B2(n_1579),
.C(n_1581),
.Y(n_13275)
);

OAI21x1_ASAP7_75t_L g13276 ( 
.A1(n_12068),
.A2(n_1581),
.B(n_1582),
.Y(n_13276)
);

OR2x2_ASAP7_75t_L g13277 ( 
.A(n_11767),
.B(n_1582),
.Y(n_13277)
);

OR2x2_ASAP7_75t_L g13278 ( 
.A(n_11769),
.B(n_11772),
.Y(n_13278)
);

NOR2xp33_ASAP7_75t_L g13279 ( 
.A(n_12527),
.B(n_1583),
.Y(n_13279)
);

NAND2xp5_ASAP7_75t_L g13280 ( 
.A(n_12642),
.B(n_1583),
.Y(n_13280)
);

A2O1A1Ixp33_ASAP7_75t_L g13281 ( 
.A1(n_12382),
.A2(n_1586),
.B(n_1584),
.C(n_1585),
.Y(n_13281)
);

INVx1_ASAP7_75t_L g13282 ( 
.A(n_12086),
.Y(n_13282)
);

OA22x2_ASAP7_75t_L g13283 ( 
.A1(n_12001),
.A2(n_1588),
.B1(n_1584),
.B2(n_1587),
.Y(n_13283)
);

INVx5_ASAP7_75t_L g13284 ( 
.A(n_12202),
.Y(n_13284)
);

AND2x2_ASAP7_75t_L g13285 ( 
.A(n_12369),
.B(n_1589),
.Y(n_13285)
);

NAND2xp5_ASAP7_75t_L g13286 ( 
.A(n_12648),
.B(n_1589),
.Y(n_13286)
);

INVx1_ASAP7_75t_L g13287 ( 
.A(n_12093),
.Y(n_13287)
);

OAI21x1_ASAP7_75t_L g13288 ( 
.A1(n_12337),
.A2(n_1590),
.B(n_1591),
.Y(n_13288)
);

OAI21x1_ASAP7_75t_L g13289 ( 
.A1(n_12478),
.A2(n_1590),
.B(n_1591),
.Y(n_13289)
);

BUFx2_ASAP7_75t_L g13290 ( 
.A(n_12177),
.Y(n_13290)
);

AND2x2_ASAP7_75t_L g13291 ( 
.A(n_12369),
.B(n_1592),
.Y(n_13291)
);

AOI21xp5_ASAP7_75t_L g13292 ( 
.A1(n_11948),
.A2(n_1593),
.B(n_1594),
.Y(n_13292)
);

NAND2xp5_ASAP7_75t_L g13293 ( 
.A(n_12657),
.B(n_1593),
.Y(n_13293)
);

O2A1O1Ixp5_ASAP7_75t_L g13294 ( 
.A1(n_11855),
.A2(n_1597),
.B(n_1595),
.C(n_1596),
.Y(n_13294)
);

AOI21xp5_ASAP7_75t_L g13295 ( 
.A1(n_12002),
.A2(n_1596),
.B(n_1597),
.Y(n_13295)
);

NAND2xp5_ASAP7_75t_L g13296 ( 
.A(n_12659),
.B(n_1598),
.Y(n_13296)
);

OAI21xp5_ASAP7_75t_L g13297 ( 
.A1(n_11991),
.A2(n_12260),
.B(n_12210),
.Y(n_13297)
);

AOI21xp5_ASAP7_75t_L g13298 ( 
.A1(n_12294),
.A2(n_1598),
.B(n_1599),
.Y(n_13298)
);

OAI22xp5_ASAP7_75t_L g13299 ( 
.A1(n_11833),
.A2(n_1601),
.B1(n_1599),
.B2(n_1600),
.Y(n_13299)
);

INVx5_ASAP7_75t_L g13300 ( 
.A(n_12079),
.Y(n_13300)
);

AOI21xp5_ASAP7_75t_L g13301 ( 
.A1(n_12271),
.A2(n_1601),
.B(n_1602),
.Y(n_13301)
);

OAI21x1_ASAP7_75t_L g13302 ( 
.A1(n_12179),
.A2(n_1602),
.B(n_1603),
.Y(n_13302)
);

INVx2_ASAP7_75t_L g13303 ( 
.A(n_12100),
.Y(n_13303)
);

NAND2xp5_ASAP7_75t_L g13304 ( 
.A(n_12663),
.B(n_1603),
.Y(n_13304)
);

AO31x2_ASAP7_75t_L g13305 ( 
.A1(n_12223),
.A2(n_1607),
.A3(n_1604),
.B(n_1605),
.Y(n_13305)
);

AND2x4_ASAP7_75t_L g13306 ( 
.A(n_12204),
.B(n_1604),
.Y(n_13306)
);

AOI21xp5_ASAP7_75t_SL g13307 ( 
.A1(n_12203),
.A2(n_1605),
.B(n_1607),
.Y(n_13307)
);

NAND2xp5_ASAP7_75t_L g13308 ( 
.A(n_12669),
.B(n_1608),
.Y(n_13308)
);

AOI211x1_ASAP7_75t_L g13309 ( 
.A1(n_11846),
.A2(n_11755),
.B(n_12376),
.C(n_12436),
.Y(n_13309)
);

AO31x2_ASAP7_75t_L g13310 ( 
.A1(n_12242),
.A2(n_1611),
.A3(n_1609),
.B(n_1610),
.Y(n_13310)
);

INVx2_ASAP7_75t_L g13311 ( 
.A(n_11810),
.Y(n_13311)
);

OAI21x1_ASAP7_75t_SL g13312 ( 
.A1(n_12422),
.A2(n_1609),
.B(n_1611),
.Y(n_13312)
);

A2O1A1Ixp33_ASAP7_75t_L g13313 ( 
.A1(n_12306),
.A2(n_1614),
.B(n_1612),
.C(n_1613),
.Y(n_13313)
);

NOR2xp33_ASAP7_75t_L g13314 ( 
.A(n_12540),
.B(n_1612),
.Y(n_13314)
);

NAND2xp5_ASAP7_75t_SL g13315 ( 
.A(n_12244),
.B(n_12061),
.Y(n_13315)
);

INVxp67_ASAP7_75t_L g13316 ( 
.A(n_11811),
.Y(n_13316)
);

BUFx2_ASAP7_75t_L g13317 ( 
.A(n_12132),
.Y(n_13317)
);

OAI21x1_ASAP7_75t_L g13318 ( 
.A1(n_12340),
.A2(n_1613),
.B(n_1615),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_11971),
.Y(n_13319)
);

AND2x2_ASAP7_75t_L g13320 ( 
.A(n_11764),
.B(n_1615),
.Y(n_13320)
);

BUFx3_ASAP7_75t_L g13321 ( 
.A(n_12184),
.Y(n_13321)
);

BUFx3_ASAP7_75t_L g13322 ( 
.A(n_11940),
.Y(n_13322)
);

OAI21x1_ASAP7_75t_SL g13323 ( 
.A1(n_12424),
.A2(n_1616),
.B(n_1617),
.Y(n_13323)
);

INVx1_ASAP7_75t_L g13324 ( 
.A(n_11973),
.Y(n_13324)
);

NAND2x1p5_ASAP7_75t_L g13325 ( 
.A(n_11891),
.B(n_1616),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_11969),
.Y(n_13326)
);

NAND2xp5_ASAP7_75t_L g13327 ( 
.A(n_12688),
.B(n_1617),
.Y(n_13327)
);

OAI21x1_ASAP7_75t_L g13328 ( 
.A1(n_12346),
.A2(n_1618),
.B(n_1619),
.Y(n_13328)
);

OAI22xp5_ASAP7_75t_L g13329 ( 
.A1(n_12339),
.A2(n_1620),
.B1(n_1618),
.B2(n_1619),
.Y(n_13329)
);

A2O1A1Ixp33_ASAP7_75t_L g13330 ( 
.A1(n_12406),
.A2(n_1622),
.B(n_1620),
.C(n_1621),
.Y(n_13330)
);

OAI22xp5_ASAP7_75t_L g13331 ( 
.A1(n_11957),
.A2(n_1624),
.B1(n_1621),
.B2(n_1622),
.Y(n_13331)
);

NAND2xp5_ASAP7_75t_SL g13332 ( 
.A(n_12244),
.B(n_1624),
.Y(n_13332)
);

BUFx2_ASAP7_75t_L g13333 ( 
.A(n_11843),
.Y(n_13333)
);

NAND2xp5_ASAP7_75t_L g13334 ( 
.A(n_12560),
.B(n_1625),
.Y(n_13334)
);

AOI21xp5_ASAP7_75t_L g13335 ( 
.A1(n_12411),
.A2(n_1625),
.B(n_1626),
.Y(n_13335)
);

OR2x2_ASAP7_75t_L g13336 ( 
.A(n_11814),
.B(n_1626),
.Y(n_13336)
);

OAI21x1_ASAP7_75t_L g13337 ( 
.A1(n_12483),
.A2(n_1627),
.B(n_1628),
.Y(n_13337)
);

NAND2xp5_ASAP7_75t_SL g13338 ( 
.A(n_12194),
.B(n_1627),
.Y(n_13338)
);

INVx3_ASAP7_75t_L g13339 ( 
.A(n_12138),
.Y(n_13339)
);

OAI21x1_ASAP7_75t_L g13340 ( 
.A1(n_12119),
.A2(n_1628),
.B(n_1629),
.Y(n_13340)
);

OAI22xp5_ASAP7_75t_L g13341 ( 
.A1(n_12044),
.A2(n_1631),
.B1(n_1629),
.B2(n_1630),
.Y(n_13341)
);

NAND2xp5_ASAP7_75t_L g13342 ( 
.A(n_12601),
.B(n_1630),
.Y(n_13342)
);

OR2x2_ASAP7_75t_L g13343 ( 
.A(n_11815),
.B(n_1631),
.Y(n_13343)
);

NAND2xp5_ASAP7_75t_SL g13344 ( 
.A(n_12284),
.B(n_1632),
.Y(n_13344)
);

NAND2xp5_ASAP7_75t_L g13345 ( 
.A(n_12610),
.B(n_12611),
.Y(n_13345)
);

AOI21xp5_ASAP7_75t_L g13346 ( 
.A1(n_12064),
.A2(n_1632),
.B(n_1633),
.Y(n_13346)
);

A2O1A1Ixp33_ASAP7_75t_L g13347 ( 
.A1(n_12500),
.A2(n_1635),
.B(n_1633),
.C(n_1634),
.Y(n_13347)
);

INVx3_ASAP7_75t_L g13348 ( 
.A(n_11761),
.Y(n_13348)
);

NAND2xp5_ASAP7_75t_L g13349 ( 
.A(n_12628),
.B(n_1634),
.Y(n_13349)
);

INVx5_ASAP7_75t_L g13350 ( 
.A(n_11940),
.Y(n_13350)
);

NOR2xp33_ASAP7_75t_L g13351 ( 
.A(n_12646),
.B(n_1635),
.Y(n_13351)
);

NAND2xp5_ASAP7_75t_L g13352 ( 
.A(n_12662),
.B(n_1636),
.Y(n_13352)
);

OAI21x1_ASAP7_75t_L g13353 ( 
.A1(n_12142),
.A2(n_1636),
.B(n_1637),
.Y(n_13353)
);

AOI21xp5_ASAP7_75t_L g13354 ( 
.A1(n_11923),
.A2(n_1637),
.B(n_1638),
.Y(n_13354)
);

INVx1_ASAP7_75t_SL g13355 ( 
.A(n_11825),
.Y(n_13355)
);

AOI21x1_ASAP7_75t_L g13356 ( 
.A1(n_12089),
.A2(n_1638),
.B(n_1639),
.Y(n_13356)
);

NAND2xp5_ASAP7_75t_L g13357 ( 
.A(n_12664),
.B(n_1640),
.Y(n_13357)
);

OAI21xp5_ASAP7_75t_L g13358 ( 
.A1(n_12487),
.A2(n_1640),
.B(n_1641),
.Y(n_13358)
);

OAI21x1_ASAP7_75t_L g13359 ( 
.A1(n_11943),
.A2(n_1642),
.B(n_1643),
.Y(n_13359)
);

NAND2xp5_ASAP7_75t_L g13360 ( 
.A(n_12666),
.B(n_1642),
.Y(n_13360)
);

AOI21xp5_ASAP7_75t_L g13361 ( 
.A1(n_11923),
.A2(n_1643),
.B(n_1644),
.Y(n_13361)
);

NAND2xp5_ASAP7_75t_L g13362 ( 
.A(n_12671),
.B(n_1644),
.Y(n_13362)
);

AO31x2_ASAP7_75t_L g13363 ( 
.A1(n_12003),
.A2(n_1647),
.A3(n_1645),
.B(n_1646),
.Y(n_13363)
);

AOI21xp5_ASAP7_75t_L g13364 ( 
.A1(n_11962),
.A2(n_1645),
.B(n_1646),
.Y(n_13364)
);

INVx8_ASAP7_75t_L g13365 ( 
.A(n_11787),
.Y(n_13365)
);

OAI21x1_ASAP7_75t_L g13366 ( 
.A1(n_11947),
.A2(n_1647),
.B(n_1648),
.Y(n_13366)
);

NAND2xp5_ASAP7_75t_L g13367 ( 
.A(n_12674),
.B(n_1648),
.Y(n_13367)
);

OAI21x1_ASAP7_75t_L g13368 ( 
.A1(n_12469),
.A2(n_1649),
.B(n_1650),
.Y(n_13368)
);

NAND2xp5_ASAP7_75t_L g13369 ( 
.A(n_12680),
.B(n_1650),
.Y(n_13369)
);

OAI21x1_ASAP7_75t_L g13370 ( 
.A1(n_12300),
.A2(n_1651),
.B(n_1652),
.Y(n_13370)
);

INVx1_ASAP7_75t_L g13371 ( 
.A(n_11968),
.Y(n_13371)
);

INVxp67_ASAP7_75t_SL g13372 ( 
.A(n_11972),
.Y(n_13372)
);

NAND2xp5_ASAP7_75t_L g13373 ( 
.A(n_12362),
.B(n_1651),
.Y(n_13373)
);

OAI21x1_ASAP7_75t_L g13374 ( 
.A1(n_12465),
.A2(n_1652),
.B(n_1653),
.Y(n_13374)
);

OAI21xp5_ASAP7_75t_L g13375 ( 
.A1(n_12236),
.A2(n_1654),
.B(n_1655),
.Y(n_13375)
);

NAND2xp5_ASAP7_75t_L g13376 ( 
.A(n_12366),
.B(n_11788),
.Y(n_13376)
);

INVx2_ASAP7_75t_L g13377 ( 
.A(n_11913),
.Y(n_13377)
);

BUFx6f_ASAP7_75t_L g13378 ( 
.A(n_11787),
.Y(n_13378)
);

NAND2xp5_ASAP7_75t_SL g13379 ( 
.A(n_12284),
.B(n_1654),
.Y(n_13379)
);

INVx2_ASAP7_75t_SL g13380 ( 
.A(n_12645),
.Y(n_13380)
);

OAI21x1_ASAP7_75t_L g13381 ( 
.A1(n_12239),
.A2(n_1655),
.B(n_1656),
.Y(n_13381)
);

AOI22xp33_ASAP7_75t_SL g13382 ( 
.A1(n_11857),
.A2(n_1658),
.B1(n_1656),
.B2(n_1657),
.Y(n_13382)
);

AO21x1_ASAP7_75t_L g13383 ( 
.A1(n_12133),
.A2(n_1657),
.B(n_1658),
.Y(n_13383)
);

INVx2_ASAP7_75t_L g13384 ( 
.A(n_11820),
.Y(n_13384)
);

OAI22xp5_ASAP7_75t_L g13385 ( 
.A1(n_12386),
.A2(n_12417),
.B1(n_12419),
.B2(n_12380),
.Y(n_13385)
);

OAI21x1_ASAP7_75t_L g13386 ( 
.A1(n_12264),
.A2(n_1659),
.B(n_1660),
.Y(n_13386)
);

NAND2xp5_ASAP7_75t_L g13387 ( 
.A(n_11911),
.B(n_1659),
.Y(n_13387)
);

NAND2x1_ASAP7_75t_L g13388 ( 
.A(n_12139),
.B(n_1660),
.Y(n_13388)
);

INVx1_ASAP7_75t_L g13389 ( 
.A(n_11789),
.Y(n_13389)
);

OAI21x1_ASAP7_75t_L g13390 ( 
.A1(n_12456),
.A2(n_1661),
.B(n_1662),
.Y(n_13390)
);

AOI21x1_ASAP7_75t_L g13391 ( 
.A1(n_12075),
.A2(n_1661),
.B(n_1662),
.Y(n_13391)
);

OAI21xp5_ASAP7_75t_L g13392 ( 
.A1(n_12056),
.A2(n_1663),
.B(n_1664),
.Y(n_13392)
);

AOI21xp5_ASAP7_75t_L g13393 ( 
.A1(n_11962),
.A2(n_1663),
.B(n_1664),
.Y(n_13393)
);

NAND2xp5_ASAP7_75t_L g13394 ( 
.A(n_12169),
.B(n_1665),
.Y(n_13394)
);

NAND2xp5_ASAP7_75t_L g13395 ( 
.A(n_12181),
.B(n_1665),
.Y(n_13395)
);

AO31x2_ASAP7_75t_L g13396 ( 
.A1(n_12027),
.A2(n_1668),
.A3(n_1666),
.B(n_1667),
.Y(n_13396)
);

AO31x2_ASAP7_75t_L g13397 ( 
.A1(n_12477),
.A2(n_1669),
.A3(n_1666),
.B(n_1668),
.Y(n_13397)
);

AND2x2_ASAP7_75t_L g13398 ( 
.A(n_12314),
.B(n_1669),
.Y(n_13398)
);

NAND2xp5_ASAP7_75t_L g13399 ( 
.A(n_12186),
.B(n_1670),
.Y(n_13399)
);

AND2x2_ASAP7_75t_SL g13400 ( 
.A(n_12584),
.B(n_1670),
.Y(n_13400)
);

NOR4xp25_ASAP7_75t_L g13401 ( 
.A(n_12035),
.B(n_1673),
.C(n_1671),
.D(n_1672),
.Y(n_13401)
);

AO31x2_ASAP7_75t_L g13402 ( 
.A1(n_12114),
.A2(n_1673),
.A3(n_1671),
.B(n_1672),
.Y(n_13402)
);

INVx1_ASAP7_75t_L g13403 ( 
.A(n_11960),
.Y(n_13403)
);

OAI21xp5_ASAP7_75t_L g13404 ( 
.A1(n_12459),
.A2(n_12017),
.B(n_12016),
.Y(n_13404)
);

OAI22xp5_ASAP7_75t_L g13405 ( 
.A1(n_12309),
.A2(n_12262),
.B1(n_11874),
.B2(n_11920),
.Y(n_13405)
);

INVx1_ASAP7_75t_L g13406 ( 
.A(n_11980),
.Y(n_13406)
);

OAI21x1_ASAP7_75t_L g13407 ( 
.A1(n_12495),
.A2(n_1674),
.B(n_1676),
.Y(n_13407)
);

AOI21xp5_ASAP7_75t_L g13408 ( 
.A1(n_12024),
.A2(n_1674),
.B(n_1676),
.Y(n_13408)
);

OAI21x1_ASAP7_75t_L g13409 ( 
.A1(n_12208),
.A2(n_1677),
.B(n_1678),
.Y(n_13409)
);

OAI21x1_ASAP7_75t_L g13410 ( 
.A1(n_12217),
.A2(n_1677),
.B(n_1678),
.Y(n_13410)
);

AOI21x1_ASAP7_75t_SL g13411 ( 
.A1(n_12218),
.A2(n_1679),
.B(n_1680),
.Y(n_13411)
);

AOI21xp5_ASAP7_75t_L g13412 ( 
.A1(n_12170),
.A2(n_1680),
.B(n_1681),
.Y(n_13412)
);

OAI22xp5_ASAP7_75t_L g13413 ( 
.A1(n_11871),
.A2(n_1683),
.B1(n_1681),
.B2(n_1682),
.Y(n_13413)
);

OAI21xp5_ASAP7_75t_SL g13414 ( 
.A1(n_12098),
.A2(n_1682),
.B(n_1683),
.Y(n_13414)
);

OAI21x1_ASAP7_75t_L g13415 ( 
.A1(n_12221),
.A2(n_1684),
.B(n_1685),
.Y(n_13415)
);

CKINVDCx5p33_ASAP7_75t_R g13416 ( 
.A(n_11918),
.Y(n_13416)
);

NAND2xp5_ASAP7_75t_L g13417 ( 
.A(n_12238),
.B(n_1684),
.Y(n_13417)
);

AO22x2_ASAP7_75t_L g13418 ( 
.A1(n_12549),
.A2(n_1688),
.B1(n_1686),
.B2(n_1687),
.Y(n_13418)
);

OAI21x1_ASAP7_75t_L g13419 ( 
.A1(n_12245),
.A2(n_1686),
.B(n_1687),
.Y(n_13419)
);

INVx1_ASAP7_75t_L g13420 ( 
.A(n_12137),
.Y(n_13420)
);

NAND2xp5_ASAP7_75t_L g13421 ( 
.A(n_12250),
.B(n_1688),
.Y(n_13421)
);

AOI21xp5_ASAP7_75t_L g13422 ( 
.A1(n_11809),
.A2(n_1689),
.B(n_1690),
.Y(n_13422)
);

OAI21x1_ASAP7_75t_L g13423 ( 
.A1(n_12267),
.A2(n_1689),
.B(n_1690),
.Y(n_13423)
);

AOI22xp5_ASAP7_75t_L g13424 ( 
.A1(n_12368),
.A2(n_12572),
.B1(n_12596),
.B2(n_12556),
.Y(n_13424)
);

BUFx12f_ASAP7_75t_SL g13425 ( 
.A(n_11803),
.Y(n_13425)
);

NOR2x1_ASAP7_75t_SL g13426 ( 
.A(n_12275),
.B(n_12139),
.Y(n_13426)
);

O2A1O1Ixp5_ASAP7_75t_L g13427 ( 
.A1(n_12619),
.A2(n_1693),
.B(n_1691),
.C(n_1692),
.Y(n_13427)
);

OAI21xp5_ASAP7_75t_L g13428 ( 
.A1(n_12102),
.A2(n_1691),
.B(n_1692),
.Y(n_13428)
);

INVx2_ASAP7_75t_L g13429 ( 
.A(n_11793),
.Y(n_13429)
);

A2O1A1Ixp33_ASAP7_75t_L g13430 ( 
.A1(n_12446),
.A2(n_1695),
.B(n_1693),
.C(n_1694),
.Y(n_13430)
);

OAI21xp5_ASAP7_75t_L g13431 ( 
.A1(n_12116),
.A2(n_1694),
.B(n_1695),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_12433),
.B(n_1696),
.Y(n_13432)
);

INVx2_ASAP7_75t_SL g13433 ( 
.A(n_12599),
.Y(n_13433)
);

AOI21xp5_ASAP7_75t_SL g13434 ( 
.A1(n_11995),
.A2(n_1697),
.B(n_1698),
.Y(n_13434)
);

AO21x1_ASAP7_75t_L g13435 ( 
.A1(n_12643),
.A2(n_1697),
.B(n_1698),
.Y(n_13435)
);

OAI222xp33_ASAP7_75t_L g13436 ( 
.A1(n_12620),
.A2(n_1701),
.B1(n_1703),
.B2(n_1699),
.C1(n_1700),
.C2(n_1702),
.Y(n_13436)
);

BUFx3_ASAP7_75t_L g13437 ( 
.A(n_12599),
.Y(n_13437)
);

OAI21x1_ASAP7_75t_L g13438 ( 
.A1(n_12293),
.A2(n_1699),
.B(n_1701),
.Y(n_13438)
);

INVxp67_ASAP7_75t_SL g13439 ( 
.A(n_11996),
.Y(n_13439)
);

AO21x1_ASAP7_75t_L g13440 ( 
.A1(n_12351),
.A2(n_12255),
.B(n_12164),
.Y(n_13440)
);

OAI22xp5_ASAP7_75t_L g13441 ( 
.A1(n_12450),
.A2(n_12652),
.B1(n_12682),
.B2(n_12639),
.Y(n_13441)
);

OAI22x1_ASAP7_75t_L g13442 ( 
.A1(n_12521),
.A2(n_1704),
.B1(n_1702),
.B2(n_1703),
.Y(n_13442)
);

AND2x2_ASAP7_75t_L g13443 ( 
.A(n_11756),
.B(n_1704),
.Y(n_13443)
);

AOI21xp5_ASAP7_75t_L g13444 ( 
.A1(n_12686),
.A2(n_1705),
.B(n_1706),
.Y(n_13444)
);

NAND2xp33_ASAP7_75t_L g13445 ( 
.A(n_11897),
.B(n_1706),
.Y(n_13445)
);

NAND2xp5_ASAP7_75t_L g13446 ( 
.A(n_12325),
.B(n_1707),
.Y(n_13446)
);

AOI21xp5_ASAP7_75t_SL g13447 ( 
.A1(n_12471),
.A2(n_1707),
.B(n_1708),
.Y(n_13447)
);

OAI21x1_ASAP7_75t_L g13448 ( 
.A1(n_12327),
.A2(n_1708),
.B(n_1709),
.Y(n_13448)
);

AOI21x1_ASAP7_75t_L g13449 ( 
.A1(n_11908),
.A2(n_1709),
.B(n_1710),
.Y(n_13449)
);

AND2x2_ASAP7_75t_L g13450 ( 
.A(n_12513),
.B(n_1710),
.Y(n_13450)
);

INVx1_ASAP7_75t_L g13451 ( 
.A(n_11835),
.Y(n_13451)
);

INVx1_ASAP7_75t_L g13452 ( 
.A(n_12400),
.Y(n_13452)
);

AO31x2_ASAP7_75t_L g13453 ( 
.A1(n_12087),
.A2(n_1713),
.A3(n_1711),
.B(n_1712),
.Y(n_13453)
);

INVx6_ASAP7_75t_SL g13454 ( 
.A(n_12533),
.Y(n_13454)
);

NAND2xp5_ASAP7_75t_L g13455 ( 
.A(n_12331),
.B(n_1711),
.Y(n_13455)
);

INVx3_ASAP7_75t_SL g13456 ( 
.A(n_12036),
.Y(n_13456)
);

AND2x2_ASAP7_75t_L g13457 ( 
.A(n_12541),
.B(n_1712),
.Y(n_13457)
);

INVx1_ASAP7_75t_L g13458 ( 
.A(n_12322),
.Y(n_13458)
);

BUFx3_ASAP7_75t_L g13459 ( 
.A(n_11803),
.Y(n_13459)
);

OAI21x1_ASAP7_75t_L g13460 ( 
.A1(n_12348),
.A2(n_1713),
.B(n_1714),
.Y(n_13460)
);

AO31x2_ASAP7_75t_L g13461 ( 
.A1(n_12276),
.A2(n_1716),
.A3(n_1714),
.B(n_1715),
.Y(n_13461)
);

INVx2_ASAP7_75t_SL g13462 ( 
.A(n_12571),
.Y(n_13462)
);

INVx2_ASAP7_75t_L g13463 ( 
.A(n_12129),
.Y(n_13463)
);

BUFx2_ASAP7_75t_L g13464 ( 
.A(n_12676),
.Y(n_13464)
);

NAND2x1_ASAP7_75t_L g13465 ( 
.A(n_12305),
.B(n_1717),
.Y(n_13465)
);

OAI21x1_ASAP7_75t_L g13466 ( 
.A1(n_12352),
.A2(n_1717),
.B(n_1718),
.Y(n_13466)
);

INVxp67_ASAP7_75t_L g13467 ( 
.A(n_12359),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_12375),
.Y(n_13468)
);

INVx1_ASAP7_75t_L g13469 ( 
.A(n_12381),
.Y(n_13469)
);

INVx1_ASAP7_75t_L g13470 ( 
.A(n_12074),
.Y(n_13470)
);

NAND2xp5_ASAP7_75t_L g13471 ( 
.A(n_12394),
.B(n_1718),
.Y(n_13471)
);

AOI21xp5_ASAP7_75t_L g13472 ( 
.A1(n_12071),
.A2(n_1719),
.B(n_1720),
.Y(n_13472)
);

OAI21xp5_ASAP7_75t_L g13473 ( 
.A1(n_12121),
.A2(n_1719),
.B(n_1720),
.Y(n_13473)
);

INVx1_ASAP7_75t_L g13474 ( 
.A(n_12389),
.Y(n_13474)
);

AO32x2_ASAP7_75t_L g13475 ( 
.A1(n_11936),
.A2(n_1724),
.A3(n_1721),
.B1(n_1723),
.B2(n_1725),
.Y(n_13475)
);

BUFx3_ASAP7_75t_L g13476 ( 
.A(n_12707),
.Y(n_13476)
);

HB1xp67_ASAP7_75t_L g13477 ( 
.A(n_12831),
.Y(n_13477)
);

BUFx3_ASAP7_75t_L g13478 ( 
.A(n_13238),
.Y(n_13478)
);

OAI21x1_ASAP7_75t_L g13479 ( 
.A1(n_12795),
.A2(n_12405),
.B(n_12396),
.Y(n_13479)
);

BUFx4_ASAP7_75t_SL g13480 ( 
.A(n_13085),
.Y(n_13480)
);

INVx6_ASAP7_75t_L g13481 ( 
.A(n_13004),
.Y(n_13481)
);

BUFx6f_ASAP7_75t_L g13482 ( 
.A(n_13087),
.Y(n_13482)
);

INVxp67_ASAP7_75t_SL g13483 ( 
.A(n_12749),
.Y(n_13483)
);

BUFx2_ASAP7_75t_L g13484 ( 
.A(n_13017),
.Y(n_13484)
);

AND2x4_ASAP7_75t_L g13485 ( 
.A(n_13130),
.B(n_12656),
.Y(n_13485)
);

BUFx4_ASAP7_75t_SL g13486 ( 
.A(n_12931),
.Y(n_13486)
);

BUFx3_ASAP7_75t_L g13487 ( 
.A(n_12942),
.Y(n_13487)
);

INVx1_ASAP7_75t_L g13488 ( 
.A(n_12691),
.Y(n_13488)
);

AO21x2_ASAP7_75t_L g13489 ( 
.A1(n_13372),
.A2(n_12356),
.B(n_11965),
.Y(n_13489)
);

BUFx3_ASAP7_75t_L g13490 ( 
.A(n_13321),
.Y(n_13490)
);

INVxp67_ASAP7_75t_SL g13491 ( 
.A(n_13173),
.Y(n_13491)
);

BUFx3_ASAP7_75t_L g13492 ( 
.A(n_12760),
.Y(n_13492)
);

HB1xp67_ASAP7_75t_L g13493 ( 
.A(n_12944),
.Y(n_13493)
);

BUFx3_ASAP7_75t_L g13494 ( 
.A(n_12760),
.Y(n_13494)
);

INVx6_ASAP7_75t_L g13495 ( 
.A(n_13015),
.Y(n_13495)
);

INVx1_ASAP7_75t_SL g13496 ( 
.A(n_13456),
.Y(n_13496)
);

BUFx6f_ASAP7_75t_L g13497 ( 
.A(n_13087),
.Y(n_13497)
);

NOR2x1_ASAP7_75t_R g13498 ( 
.A(n_13300),
.B(n_12136),
.Y(n_13498)
);

OAI21xp5_ASAP7_75t_L g13499 ( 
.A1(n_12726),
.A2(n_12055),
.B(n_12263),
.Y(n_13499)
);

INVx1_ASAP7_75t_L g13500 ( 
.A(n_12695),
.Y(n_13500)
);

OAI21x1_ASAP7_75t_L g13501 ( 
.A1(n_12998),
.A2(n_12398),
.B(n_12395),
.Y(n_13501)
);

INVx6_ASAP7_75t_L g13502 ( 
.A(n_13107),
.Y(n_13502)
);

INVxp67_ASAP7_75t_SL g13503 ( 
.A(n_12777),
.Y(n_13503)
);

NAND2xp5_ASAP7_75t_L g13504 ( 
.A(n_13251),
.B(n_11902),
.Y(n_13504)
);

BUFx3_ASAP7_75t_L g13505 ( 
.A(n_12965),
.Y(n_13505)
);

OAI21x1_ASAP7_75t_L g13506 ( 
.A1(n_12706),
.A2(n_12401),
.B(n_12408),
.Y(n_13506)
);

OR2x6_ASAP7_75t_L g13507 ( 
.A(n_13126),
.B(n_12672),
.Y(n_13507)
);

INVx1_ASAP7_75t_L g13508 ( 
.A(n_12708),
.Y(n_13508)
);

BUFx5_ASAP7_75t_L g13509 ( 
.A(n_13250),
.Y(n_13509)
);

OA21x2_ASAP7_75t_L g13510 ( 
.A1(n_12890),
.A2(n_12415),
.B(n_12385),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_12713),
.Y(n_13511)
);

OAI21x1_ASAP7_75t_L g13512 ( 
.A1(n_12710),
.A2(n_12383),
.B(n_12447),
.Y(n_13512)
);

BUFx6f_ASAP7_75t_L g13513 ( 
.A(n_13378),
.Y(n_13513)
);

INVx2_ASAP7_75t_L g13514 ( 
.A(n_12802),
.Y(n_13514)
);

BUFx5_ASAP7_75t_L g13515 ( 
.A(n_13437),
.Y(n_13515)
);

AO21x2_ASAP7_75t_L g13516 ( 
.A1(n_13451),
.A2(n_12272),
.B(n_12268),
.Y(n_13516)
);

AND2x4_ASAP7_75t_L g13517 ( 
.A(n_12768),
.B(n_12297),
.Y(n_13517)
);

INVx2_ASAP7_75t_SL g13518 ( 
.A(n_13350),
.Y(n_13518)
);

INVx2_ASAP7_75t_SL g13519 ( 
.A(n_13350),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_12728),
.Y(n_13520)
);

AND2x4_ASAP7_75t_L g13521 ( 
.A(n_13129),
.B(n_12297),
.Y(n_13521)
);

OAI21x1_ASAP7_75t_L g13522 ( 
.A1(n_12723),
.A2(n_12429),
.B(n_12425),
.Y(n_13522)
);

OAI21xp5_ASAP7_75t_L g13523 ( 
.A1(n_12801),
.A2(n_11916),
.B(n_11984),
.Y(n_13523)
);

OAI21x1_ASAP7_75t_L g13524 ( 
.A1(n_12880),
.A2(n_13026),
.B(n_12714),
.Y(n_13524)
);

INVx2_ASAP7_75t_L g13525 ( 
.A(n_12905),
.Y(n_13525)
);

BUFx2_ASAP7_75t_SL g13526 ( 
.A(n_12832),
.Y(n_13526)
);

INVx2_ASAP7_75t_SL g13527 ( 
.A(n_13322),
.Y(n_13527)
);

INVx1_ASAP7_75t_L g13528 ( 
.A(n_12758),
.Y(n_13528)
);

NOR2xp67_ASAP7_75t_SL g13529 ( 
.A(n_13180),
.B(n_12449),
.Y(n_13529)
);

AO21x2_ASAP7_75t_L g13530 ( 
.A1(n_12696),
.A2(n_11778),
.B(n_11765),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_12910),
.Y(n_13531)
);

AND2x4_ASAP7_75t_L g13532 ( 
.A(n_12762),
.B(n_11786),
.Y(n_13532)
);

OAI21x1_ASAP7_75t_L g13533 ( 
.A1(n_12814),
.A2(n_12437),
.B(n_12343),
.Y(n_13533)
);

CKINVDCx11_ASAP7_75t_R g13534 ( 
.A(n_12873),
.Y(n_13534)
);

NAND2x1p5_ASAP7_75t_L g13535 ( 
.A(n_13141),
.B(n_12266),
.Y(n_13535)
);

NOR2xp33_ASAP7_75t_SL g13536 ( 
.A(n_13300),
.B(n_11762),
.Y(n_13536)
);

AND2x2_ASAP7_75t_L g13537 ( 
.A(n_12967),
.B(n_12847),
.Y(n_13537)
);

AOI22xp33_ASAP7_75t_SL g13538 ( 
.A1(n_12792),
.A2(n_12453),
.B1(n_11850),
.B2(n_12021),
.Y(n_13538)
);

INVx1_ASAP7_75t_L g13539 ( 
.A(n_12939),
.Y(n_13539)
);

AO21x2_ASAP7_75t_L g13540 ( 
.A1(n_12765),
.A2(n_12615),
.B(n_12585),
.Y(n_13540)
);

INVx1_ASAP7_75t_SL g13541 ( 
.A(n_13270),
.Y(n_13541)
);

AO21x2_ASAP7_75t_L g13542 ( 
.A1(n_12766),
.A2(n_11818),
.B(n_12092),
.Y(n_13542)
);

BUFx3_ASAP7_75t_L g13543 ( 
.A(n_13012),
.Y(n_13543)
);

AOI22x1_ASAP7_75t_L g13544 ( 
.A1(n_13032),
.A2(n_12416),
.B1(n_12182),
.B2(n_12189),
.Y(n_13544)
);

INVx1_ASAP7_75t_L g13545 ( 
.A(n_12989),
.Y(n_13545)
);

INVx2_ASAP7_75t_SL g13546 ( 
.A(n_13317),
.Y(n_13546)
);

BUFx2_ASAP7_75t_R g13547 ( 
.A(n_13128),
.Y(n_13547)
);

OAI21x1_ASAP7_75t_L g13548 ( 
.A1(n_13027),
.A2(n_12427),
.B(n_12140),
.Y(n_13548)
);

OAI21x1_ASAP7_75t_L g13549 ( 
.A1(n_13207),
.A2(n_12338),
.B(n_11776),
.Y(n_13549)
);

OAI21x1_ASAP7_75t_L g13550 ( 
.A1(n_12885),
.A2(n_11791),
.B(n_11759),
.Y(n_13550)
);

INVx2_ASAP7_75t_SL g13551 ( 
.A(n_13348),
.Y(n_13551)
);

OAI21x1_ASAP7_75t_L g13552 ( 
.A1(n_12736),
.A2(n_11866),
.B(n_11797),
.Y(n_13552)
);

BUFx3_ASAP7_75t_L g13553 ( 
.A(n_13013),
.Y(n_13553)
);

OAI21x1_ASAP7_75t_L g13554 ( 
.A1(n_12730),
.A2(n_11876),
.B(n_11942),
.Y(n_13554)
);

OAI21xp5_ASAP7_75t_L g13555 ( 
.A1(n_12916),
.A2(n_11951),
.B(n_12288),
.Y(n_13555)
);

OAI21x1_ASAP7_75t_L g13556 ( 
.A1(n_12709),
.A2(n_12323),
.B(n_12149),
.Y(n_13556)
);

OR3x4_ASAP7_75t_SL g13557 ( 
.A(n_13439),
.B(n_12511),
.C(n_11966),
.Y(n_13557)
);

INVx1_ASAP7_75t_L g13558 ( 
.A(n_12991),
.Y(n_13558)
);

INVx1_ASAP7_75t_L g13559 ( 
.A(n_12857),
.Y(n_13559)
);

AOI22x1_ASAP7_75t_L g13560 ( 
.A1(n_12909),
.A2(n_12229),
.B1(n_11826),
.B2(n_11851),
.Y(n_13560)
);

OAI21x1_ASAP7_75t_L g13561 ( 
.A1(n_12702),
.A2(n_12285),
.B(n_12103),
.Y(n_13561)
);

INVx1_ASAP7_75t_L g13562 ( 
.A(n_12863),
.Y(n_13562)
);

AND2x4_ASAP7_75t_L g13563 ( 
.A(n_13249),
.B(n_13083),
.Y(n_13563)
);

BUFx6f_ASAP7_75t_L g13564 ( 
.A(n_13378),
.Y(n_13564)
);

OA21x2_ASAP7_75t_L g13565 ( 
.A1(n_12877),
.A2(n_12286),
.B(n_12418),
.Y(n_13565)
);

INVx2_ASAP7_75t_SL g13566 ( 
.A(n_12740),
.Y(n_13566)
);

OAI21x1_ASAP7_75t_L g13567 ( 
.A1(n_12797),
.A2(n_12307),
.B(n_12280),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_12895),
.Y(n_13568)
);

OAI21x1_ASAP7_75t_L g13569 ( 
.A1(n_12750),
.A2(n_12197),
.B(n_12183),
.Y(n_13569)
);

AO21x2_ASAP7_75t_L g13570 ( 
.A1(n_12769),
.A2(n_12131),
.B(n_12555),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_12791),
.Y(n_13571)
);

OAI21x1_ASAP7_75t_L g13572 ( 
.A1(n_12779),
.A2(n_12172),
.B(n_12554),
.Y(n_13572)
);

INVx1_ASAP7_75t_L g13573 ( 
.A(n_12828),
.Y(n_13573)
);

CKINVDCx6p67_ASAP7_75t_R g13574 ( 
.A(n_13141),
.Y(n_13574)
);

INVx1_ASAP7_75t_L g13575 ( 
.A(n_12837),
.Y(n_13575)
);

NAND2x1p5_ASAP7_75t_L g13576 ( 
.A(n_12770),
.B(n_11805),
.Y(n_13576)
);

OAI21x1_ASAP7_75t_SL g13577 ( 
.A1(n_13426),
.A2(n_12622),
.B(n_11886),
.Y(n_13577)
);

AND2x4_ASAP7_75t_L g13578 ( 
.A(n_12958),
.B(n_11860),
.Y(n_13578)
);

BUFx4f_ASAP7_75t_SL g13579 ( 
.A(n_13454),
.Y(n_13579)
);

BUFx3_ASAP7_75t_L g13580 ( 
.A(n_13248),
.Y(n_13580)
);

AND2x2_ASAP7_75t_L g13581 ( 
.A(n_13204),
.B(n_13464),
.Y(n_13581)
);

OAI21x1_ASAP7_75t_L g13582 ( 
.A1(n_12783),
.A2(n_12679),
.B(n_12350),
.Y(n_13582)
);

AOI21xp5_ASAP7_75t_L g13583 ( 
.A1(n_12817),
.A2(n_12426),
.B(n_12462),
.Y(n_13583)
);

NAND2x1p5_ASAP7_75t_L g13584 ( 
.A(n_13048),
.B(n_11860),
.Y(n_13584)
);

BUFx3_ASAP7_75t_L g13585 ( 
.A(n_13459),
.Y(n_13585)
);

CKINVDCx16_ASAP7_75t_R g13586 ( 
.A(n_12912),
.Y(n_13586)
);

BUFx6f_ASAP7_75t_L g13587 ( 
.A(n_12752),
.Y(n_13587)
);

INVx2_ASAP7_75t_L g13588 ( 
.A(n_12694),
.Y(n_13588)
);

BUFx2_ASAP7_75t_L g13589 ( 
.A(n_13333),
.Y(n_13589)
);

INVx2_ASAP7_75t_L g13590 ( 
.A(n_12742),
.Y(n_13590)
);

BUFx3_ASAP7_75t_L g13591 ( 
.A(n_12896),
.Y(n_13591)
);

HB1xp67_ASAP7_75t_L g13592 ( 
.A(n_13108),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_12840),
.Y(n_13593)
);

AO21x2_ASAP7_75t_L g13594 ( 
.A1(n_12775),
.A2(n_12667),
.B(n_12630),
.Y(n_13594)
);

OR2x2_ASAP7_75t_L g13595 ( 
.A(n_12842),
.B(n_12332),
.Y(n_13595)
);

NOR2xp33_ASAP7_75t_L g13596 ( 
.A(n_13440),
.B(n_11872),
.Y(n_13596)
);

OAI21x1_ASAP7_75t_L g13597 ( 
.A1(n_12761),
.A2(n_12289),
.B(n_12025),
.Y(n_13597)
);

OAI21xp5_ASAP7_75t_L g13598 ( 
.A1(n_12923),
.A2(n_12454),
.B(n_12227),
.Y(n_13598)
);

AND2x2_ASAP7_75t_L g13599 ( 
.A(n_13156),
.B(n_11872),
.Y(n_13599)
);

CKINVDCx5p33_ASAP7_75t_R g13600 ( 
.A(n_12826),
.Y(n_13600)
);

INVx5_ASAP7_75t_L g13601 ( 
.A(n_13098),
.Y(n_13601)
);

OAI21x1_ASAP7_75t_L g13602 ( 
.A1(n_12755),
.A2(n_12227),
.B(n_12292),
.Y(n_13602)
);

AO21x1_ASAP7_75t_L g13603 ( 
.A1(n_12854),
.A2(n_13092),
.B(n_12973),
.Y(n_13603)
);

AOI22x1_ASAP7_75t_L g13604 ( 
.A1(n_12757),
.A2(n_11880),
.B1(n_12530),
.B2(n_11830),
.Y(n_13604)
);

NAND2x1p5_ASAP7_75t_L g13605 ( 
.A(n_13169),
.B(n_11880),
.Y(n_13605)
);

INVx1_ASAP7_75t_L g13606 ( 
.A(n_12843),
.Y(n_13606)
);

HB1xp67_ASAP7_75t_L g13607 ( 
.A(n_12751),
.Y(n_13607)
);

CKINVDCx6p67_ASAP7_75t_R g13608 ( 
.A(n_13284),
.Y(n_13608)
);

BUFx3_ASAP7_75t_L g13609 ( 
.A(n_13196),
.Y(n_13609)
);

AO21x2_ASAP7_75t_L g13610 ( 
.A1(n_12816),
.A2(n_12530),
.B(n_1721),
.Y(n_13610)
);

INVx6_ASAP7_75t_L g13611 ( 
.A(n_12752),
.Y(n_13611)
);

BUFx2_ASAP7_75t_SL g13612 ( 
.A(n_13284),
.Y(n_13612)
);

AND2x4_ASAP7_75t_L g13613 ( 
.A(n_12780),
.B(n_1724),
.Y(n_13613)
);

INVx1_ASAP7_75t_L g13614 ( 
.A(n_12850),
.Y(n_13614)
);

AO21x2_ASAP7_75t_L g13615 ( 
.A1(n_12844),
.A2(n_1725),
.B(n_1726),
.Y(n_13615)
);

INVx1_ASAP7_75t_SL g13616 ( 
.A(n_13290),
.Y(n_13616)
);

INVx2_ASAP7_75t_L g13617 ( 
.A(n_12789),
.Y(n_13617)
);

NOR2xp33_ASAP7_75t_L g13618 ( 
.A(n_13239),
.B(n_1727),
.Y(n_13618)
);

BUFx6f_ASAP7_75t_L g13619 ( 
.A(n_12771),
.Y(n_13619)
);

INVx3_ASAP7_75t_L g13620 ( 
.A(n_13113),
.Y(n_13620)
);

OAI21x1_ASAP7_75t_L g13621 ( 
.A1(n_12759),
.A2(n_1727),
.B(n_1728),
.Y(n_13621)
);

NAND2xp5_ASAP7_75t_L g13622 ( 
.A(n_13117),
.B(n_1728),
.Y(n_13622)
);

INVx8_ASAP7_75t_L g13623 ( 
.A(n_13365),
.Y(n_13623)
);

CKINVDCx5p33_ASAP7_75t_R g13624 ( 
.A(n_12995),
.Y(n_13624)
);

BUFx3_ASAP7_75t_L g13625 ( 
.A(n_13210),
.Y(n_13625)
);

BUFx2_ASAP7_75t_L g13626 ( 
.A(n_13191),
.Y(n_13626)
);

NAND2x1p5_ASAP7_75t_L g13627 ( 
.A(n_13315),
.B(n_1729),
.Y(n_13627)
);

NOR2xp33_ASAP7_75t_L g13628 ( 
.A(n_13247),
.B(n_1729),
.Y(n_13628)
);

INVx1_ASAP7_75t_L g13629 ( 
.A(n_12851),
.Y(n_13629)
);

INVx2_ASAP7_75t_L g13630 ( 
.A(n_12803),
.Y(n_13630)
);

OAI21x1_ASAP7_75t_L g13631 ( 
.A1(n_12838),
.A2(n_12830),
.B(n_12829),
.Y(n_13631)
);

AO21x2_ASAP7_75t_L g13632 ( 
.A1(n_12846),
.A2(n_1730),
.B(n_1731),
.Y(n_13632)
);

CKINVDCx5p33_ASAP7_75t_R g13633 ( 
.A(n_13262),
.Y(n_13633)
);

BUFx6f_ASAP7_75t_L g13634 ( 
.A(n_12771),
.Y(n_13634)
);

HB1xp67_ASAP7_75t_L g13635 ( 
.A(n_12833),
.Y(n_13635)
);

OAI21xp5_ASAP7_75t_L g13636 ( 
.A1(n_12725),
.A2(n_1730),
.B(n_1731),
.Y(n_13636)
);

INVx8_ASAP7_75t_L g13637 ( 
.A(n_13365),
.Y(n_13637)
);

INVx2_ASAP7_75t_SL g13638 ( 
.A(n_12982),
.Y(n_13638)
);

BUFx3_ASAP7_75t_L g13639 ( 
.A(n_12867),
.Y(n_13639)
);

AO21x2_ASAP7_75t_L g13640 ( 
.A1(n_12864),
.A2(n_1732),
.B(n_1733),
.Y(n_13640)
);

OR2x6_ASAP7_75t_L g13641 ( 
.A(n_13126),
.B(n_1732),
.Y(n_13641)
);

CKINVDCx20_ASAP7_75t_R g13642 ( 
.A(n_13416),
.Y(n_13642)
);

INVx3_ASAP7_75t_L g13643 ( 
.A(n_13149),
.Y(n_13643)
);

INVx1_ASAP7_75t_L g13644 ( 
.A(n_12924),
.Y(n_13644)
);

AOI22xp5_ASAP7_75t_L g13645 ( 
.A1(n_13385),
.A2(n_1735),
.B1(n_1733),
.B2(n_1734),
.Y(n_13645)
);

AO21x2_ASAP7_75t_L g13646 ( 
.A1(n_12865),
.A2(n_1734),
.B(n_1735),
.Y(n_13646)
);

INVx2_ASAP7_75t_L g13647 ( 
.A(n_12934),
.Y(n_13647)
);

INVx3_ASAP7_75t_L g13648 ( 
.A(n_13259),
.Y(n_13648)
);

AND2x2_ASAP7_75t_L g13649 ( 
.A(n_13303),
.B(n_1736),
.Y(n_13649)
);

OAI21x1_ASAP7_75t_L g13650 ( 
.A1(n_12836),
.A2(n_1736),
.B(n_1737),
.Y(n_13650)
);

INVx2_ASAP7_75t_SL g13651 ( 
.A(n_13062),
.Y(n_13651)
);

NAND2x1p5_ASAP7_75t_L g13652 ( 
.A(n_13088),
.B(n_1737),
.Y(n_13652)
);

OAI21x1_ASAP7_75t_L g13653 ( 
.A1(n_12810),
.A2(n_1738),
.B(n_1739),
.Y(n_13653)
);

BUFx2_ASAP7_75t_SL g13654 ( 
.A(n_12790),
.Y(n_13654)
);

BUFx2_ASAP7_75t_SL g13655 ( 
.A(n_12914),
.Y(n_13655)
);

AO21x2_ASAP7_75t_L g13656 ( 
.A1(n_12876),
.A2(n_1738),
.B(n_1740),
.Y(n_13656)
);

NAND2xp5_ASAP7_75t_L g13657 ( 
.A(n_13189),
.B(n_12727),
.Y(n_13657)
);

INVx2_ASAP7_75t_SL g13658 ( 
.A(n_12911),
.Y(n_13658)
);

INVxp67_ASAP7_75t_SL g13659 ( 
.A(n_13093),
.Y(n_13659)
);

NAND2xp5_ASAP7_75t_L g13660 ( 
.A(n_13202),
.B(n_1740),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_12933),
.Y(n_13661)
);

INVx5_ASAP7_75t_SL g13662 ( 
.A(n_12867),
.Y(n_13662)
);

INVx2_ASAP7_75t_L g13663 ( 
.A(n_12978),
.Y(n_13663)
);

AND2x2_ASAP7_75t_L g13664 ( 
.A(n_13452),
.B(n_1741),
.Y(n_13664)
);

HB1xp67_ASAP7_75t_L g13665 ( 
.A(n_12979),
.Y(n_13665)
);

OAI21x1_ASAP7_75t_L g13666 ( 
.A1(n_12861),
.A2(n_1741),
.B(n_1742),
.Y(n_13666)
);

BUFx2_ASAP7_75t_L g13667 ( 
.A(n_13208),
.Y(n_13667)
);

AND2x4_ASAP7_75t_L g13668 ( 
.A(n_13199),
.B(n_1742),
.Y(n_13668)
);

BUFx12f_ASAP7_75t_L g13669 ( 
.A(n_12891),
.Y(n_13669)
);

AO21x2_ASAP7_75t_L g13670 ( 
.A1(n_12878),
.A2(n_1743),
.B(n_1744),
.Y(n_13670)
);

INVx4_ASAP7_75t_L g13671 ( 
.A(n_13024),
.Y(n_13671)
);

BUFx2_ASAP7_75t_L g13672 ( 
.A(n_13458),
.Y(n_13672)
);

BUFx12f_ASAP7_75t_L g13673 ( 
.A(n_12891),
.Y(n_13673)
);

OAI21x1_ASAP7_75t_L g13674 ( 
.A1(n_12764),
.A2(n_1743),
.B(n_1744),
.Y(n_13674)
);

BUFx2_ASAP7_75t_L g13675 ( 
.A(n_13420),
.Y(n_13675)
);

INVx3_ASAP7_75t_L g13676 ( 
.A(n_13339),
.Y(n_13676)
);

INVx3_ASAP7_75t_SL g13677 ( 
.A(n_13098),
.Y(n_13677)
);

HB1xp67_ASAP7_75t_L g13678 ( 
.A(n_13041),
.Y(n_13678)
);

OA21x2_ASAP7_75t_L g13679 ( 
.A1(n_12946),
.A2(n_1745),
.B(n_1746),
.Y(n_13679)
);

INVx2_ASAP7_75t_L g13680 ( 
.A(n_13111),
.Y(n_13680)
);

AO21x2_ASAP7_75t_L g13681 ( 
.A1(n_12879),
.A2(n_1747),
.B(n_1748),
.Y(n_13681)
);

INVx1_ASAP7_75t_L g13682 ( 
.A(n_12948),
.Y(n_13682)
);

NAND2xp5_ASAP7_75t_L g13683 ( 
.A(n_13311),
.B(n_1747),
.Y(n_13683)
);

NAND2xp5_ASAP7_75t_SL g13684 ( 
.A(n_13183),
.B(n_1748),
.Y(n_13684)
);

BUFx8_ASAP7_75t_L g13685 ( 
.A(n_13432),
.Y(n_13685)
);

INVx1_ASAP7_75t_L g13686 ( 
.A(n_12977),
.Y(n_13686)
);

AND2x4_ASAP7_75t_L g13687 ( 
.A(n_12997),
.B(n_1749),
.Y(n_13687)
);

BUFx6f_ASAP7_75t_L g13688 ( 
.A(n_12929),
.Y(n_13688)
);

OAI21xp5_ASAP7_75t_L g13689 ( 
.A1(n_12772),
.A2(n_1749),
.B(n_1750),
.Y(n_13689)
);

INVx1_ASAP7_75t_L g13690 ( 
.A(n_12990),
.Y(n_13690)
);

INVx2_ASAP7_75t_L g13691 ( 
.A(n_13178),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_13029),
.Y(n_13692)
);

INVx2_ASAP7_75t_SL g13693 ( 
.A(n_13462),
.Y(n_13693)
);

OAI21xp5_ASAP7_75t_L g13694 ( 
.A1(n_13192),
.A2(n_1750),
.B(n_1751),
.Y(n_13694)
);

INVx3_ASAP7_75t_L g13695 ( 
.A(n_12918),
.Y(n_13695)
);

INVx2_ASAP7_75t_L g13696 ( 
.A(n_13178),
.Y(n_13696)
);

AO21x2_ASAP7_75t_L g13697 ( 
.A1(n_12882),
.A2(n_1751),
.B(n_1752),
.Y(n_13697)
);

AO21x2_ASAP7_75t_L g13698 ( 
.A1(n_12893),
.A2(n_1753),
.B(n_1754),
.Y(n_13698)
);

NAND2x1p5_ASAP7_75t_L g13699 ( 
.A(n_13388),
.B(n_1753),
.Y(n_13699)
);

CKINVDCx20_ASAP7_75t_R g13700 ( 
.A(n_13425),
.Y(n_13700)
);

OR2x2_ASAP7_75t_L g13701 ( 
.A(n_13031),
.B(n_1754),
.Y(n_13701)
);

NOR2xp33_ASAP7_75t_L g13702 ( 
.A(n_13467),
.B(n_1755),
.Y(n_13702)
);

INVx6_ASAP7_75t_L g13703 ( 
.A(n_12974),
.Y(n_13703)
);

BUFx2_ASAP7_75t_SL g13704 ( 
.A(n_13068),
.Y(n_13704)
);

AND2x2_ASAP7_75t_L g13705 ( 
.A(n_13261),
.B(n_1755),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13040),
.Y(n_13706)
);

INVx2_ASAP7_75t_L g13707 ( 
.A(n_13178),
.Y(n_13707)
);

NAND2x1p5_ASAP7_75t_L g13708 ( 
.A(n_13355),
.B(n_1756),
.Y(n_13708)
);

OAI21x1_ASAP7_75t_L g13709 ( 
.A1(n_12806),
.A2(n_1756),
.B(n_1757),
.Y(n_13709)
);

BUFx3_ASAP7_75t_L g13710 ( 
.A(n_13433),
.Y(n_13710)
);

INVxp67_ASAP7_75t_SL g13711 ( 
.A(n_12952),
.Y(n_13711)
);

INVx1_ASAP7_75t_SL g13712 ( 
.A(n_13234),
.Y(n_13712)
);

BUFx12f_ASAP7_75t_L g13713 ( 
.A(n_13112),
.Y(n_13713)
);

OAI21x1_ASAP7_75t_L g13714 ( 
.A1(n_12855),
.A2(n_1758),
.B(n_1759),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_13066),
.Y(n_13715)
);

HB1xp67_ASAP7_75t_L g13716 ( 
.A(n_13078),
.Y(n_13716)
);

AO21x2_ASAP7_75t_L g13717 ( 
.A1(n_12900),
.A2(n_1759),
.B(n_1760),
.Y(n_13717)
);

INVx3_ASAP7_75t_L g13718 ( 
.A(n_12961),
.Y(n_13718)
);

INVx8_ASAP7_75t_L g13719 ( 
.A(n_13272),
.Y(n_13719)
);

OAI21x1_ASAP7_75t_L g13720 ( 
.A1(n_12856),
.A2(n_1760),
.B(n_1761),
.Y(n_13720)
);

AND2x4_ASAP7_75t_L g13721 ( 
.A(n_13101),
.B(n_1761),
.Y(n_13721)
);

INVx1_ASAP7_75t_L g13722 ( 
.A(n_13114),
.Y(n_13722)
);

BUFx3_ASAP7_75t_L g13723 ( 
.A(n_13244),
.Y(n_13723)
);

HB1xp67_ASAP7_75t_L g13724 ( 
.A(n_13218),
.Y(n_13724)
);

BUFx2_ASAP7_75t_L g13725 ( 
.A(n_13254),
.Y(n_13725)
);

OAI21x1_ASAP7_75t_L g13726 ( 
.A1(n_13106),
.A2(n_1762),
.B(n_1763),
.Y(n_13726)
);

OAI21x1_ASAP7_75t_L g13727 ( 
.A1(n_12753),
.A2(n_12827),
.B(n_12747),
.Y(n_13727)
);

OAI21x1_ASAP7_75t_L g13728 ( 
.A1(n_12969),
.A2(n_1762),
.B(n_1763),
.Y(n_13728)
);

NAND2xp5_ASAP7_75t_SL g13729 ( 
.A(n_12807),
.B(n_1764),
.Y(n_13729)
);

INVx1_ASAP7_75t_SL g13730 ( 
.A(n_13278),
.Y(n_13730)
);

NAND2x1_ASAP7_75t_L g13731 ( 
.A(n_13264),
.B(n_1764),
.Y(n_13731)
);

INVx1_ASAP7_75t_L g13732 ( 
.A(n_13178),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_13282),
.Y(n_13733)
);

AO21x2_ASAP7_75t_L g13734 ( 
.A1(n_12903),
.A2(n_1765),
.B(n_1766),
.Y(n_13734)
);

OAI21x1_ASAP7_75t_L g13735 ( 
.A1(n_13137),
.A2(n_1765),
.B(n_1766),
.Y(n_13735)
);

AO21x2_ASAP7_75t_L g13736 ( 
.A1(n_12904),
.A2(n_1767),
.B(n_1768),
.Y(n_13736)
);

INVx4_ASAP7_75t_L g13737 ( 
.A(n_12705),
.Y(n_13737)
);

INVx2_ASAP7_75t_SL g13738 ( 
.A(n_13380),
.Y(n_13738)
);

AO21x2_ASAP7_75t_L g13739 ( 
.A1(n_12739),
.A2(n_1767),
.B(n_1768),
.Y(n_13739)
);

INVx1_ASAP7_75t_L g13740 ( 
.A(n_13287),
.Y(n_13740)
);

AOI21xp5_ASAP7_75t_L g13741 ( 
.A1(n_13160),
.A2(n_1769),
.B(n_1770),
.Y(n_13741)
);

INVx5_ASAP7_75t_L g13742 ( 
.A(n_12862),
.Y(n_13742)
);

INVx3_ASAP7_75t_SL g13743 ( 
.A(n_13400),
.Y(n_13743)
);

INVx1_ASAP7_75t_L g13744 ( 
.A(n_13179),
.Y(n_13744)
);

OAI21x1_ASAP7_75t_L g13745 ( 
.A1(n_13060),
.A2(n_1769),
.B(n_1770),
.Y(n_13745)
);

AND2x4_ASAP7_75t_L g13746 ( 
.A(n_13255),
.B(n_1771),
.Y(n_13746)
);

OAI21x1_ASAP7_75t_L g13747 ( 
.A1(n_12732),
.A2(n_1771),
.B(n_1772),
.Y(n_13747)
);

INVxp33_ASAP7_75t_L g13748 ( 
.A(n_12921),
.Y(n_13748)
);

NAND2x1p5_ASAP7_75t_L g13749 ( 
.A(n_13100),
.B(n_1772),
.Y(n_13749)
);

NAND2xp5_ASAP7_75t_SL g13750 ( 
.A(n_12839),
.B(n_1773),
.Y(n_13750)
);

BUFx5_ASAP7_75t_L g13751 ( 
.A(n_13474),
.Y(n_13751)
);

INVx1_ASAP7_75t_L g13752 ( 
.A(n_12868),
.Y(n_13752)
);

AOI21x1_ASAP7_75t_L g13753 ( 
.A1(n_12959),
.A2(n_12712),
.B(n_12697),
.Y(n_13753)
);

INVx1_ASAP7_75t_L g13754 ( 
.A(n_12907),
.Y(n_13754)
);

INVx3_ASAP7_75t_L g13755 ( 
.A(n_13273),
.Y(n_13755)
);

BUFx12f_ASAP7_75t_L g13756 ( 
.A(n_13320),
.Y(n_13756)
);

INVx1_ASAP7_75t_L g13757 ( 
.A(n_13326),
.Y(n_13757)
);

AOI22x1_ASAP7_75t_L g13758 ( 
.A1(n_12823),
.A2(n_1775),
.B1(n_1773),
.B2(n_1774),
.Y(n_13758)
);

AO21x2_ASAP7_75t_L g13759 ( 
.A1(n_13422),
.A2(n_1774),
.B(n_1775),
.Y(n_13759)
);

NOR2x1_ASAP7_75t_R g13760 ( 
.A(n_12719),
.B(n_1776),
.Y(n_13760)
);

OAI21x1_ASAP7_75t_L g13761 ( 
.A1(n_12866),
.A2(n_1776),
.B(n_1777),
.Y(n_13761)
);

NAND2x1_ASAP7_75t_L g13762 ( 
.A(n_13146),
.B(n_1777),
.Y(n_13762)
);

INVx3_ASAP7_75t_L g13763 ( 
.A(n_13463),
.Y(n_13763)
);

INVx1_ASAP7_75t_L g13764 ( 
.A(n_13151),
.Y(n_13764)
);

OAI21x1_ASAP7_75t_L g13765 ( 
.A1(n_12871),
.A2(n_1778),
.B(n_1779),
.Y(n_13765)
);

AO21x2_ASAP7_75t_L g13766 ( 
.A1(n_13105),
.A2(n_1778),
.B(n_1779),
.Y(n_13766)
);

OAI21x1_ASAP7_75t_L g13767 ( 
.A1(n_12874),
.A2(n_1780),
.B(n_1781),
.Y(n_13767)
);

HB1xp67_ASAP7_75t_L g13768 ( 
.A(n_13371),
.Y(n_13768)
);

INVxp67_ASAP7_75t_SL g13769 ( 
.A(n_13319),
.Y(n_13769)
);

INVx3_ASAP7_75t_SL g13770 ( 
.A(n_12804),
.Y(n_13770)
);

INVx2_ASAP7_75t_L g13771 ( 
.A(n_13384),
.Y(n_13771)
);

INVx1_ASAP7_75t_L g13772 ( 
.A(n_12735),
.Y(n_13772)
);

OAI21x1_ASAP7_75t_L g13773 ( 
.A1(n_12884),
.A2(n_1780),
.B(n_1781),
.Y(n_13773)
);

OAI21x1_ASAP7_75t_L g13774 ( 
.A1(n_12889),
.A2(n_1782),
.B(n_1783),
.Y(n_13774)
);

AO21x2_ASAP7_75t_L g13775 ( 
.A1(n_12704),
.A2(n_1782),
.B(n_1783),
.Y(n_13775)
);

INVx1_ASAP7_75t_L g13776 ( 
.A(n_12737),
.Y(n_13776)
);

AO21x2_ASAP7_75t_L g13777 ( 
.A1(n_12721),
.A2(n_1784),
.B(n_1785),
.Y(n_13777)
);

AND2x4_ASAP7_75t_L g13778 ( 
.A(n_13377),
.B(n_1785),
.Y(n_13778)
);

INVx3_ASAP7_75t_L g13779 ( 
.A(n_13429),
.Y(n_13779)
);

OA21x2_ASAP7_75t_L g13780 ( 
.A1(n_12722),
.A2(n_1786),
.B(n_1787),
.Y(n_13780)
);

INVx1_ASAP7_75t_SL g13781 ( 
.A(n_13064),
.Y(n_13781)
);

BUFx8_ASAP7_75t_L g13782 ( 
.A(n_12860),
.Y(n_13782)
);

OAI21x1_ASAP7_75t_L g13783 ( 
.A1(n_12899),
.A2(n_1786),
.B(n_1788),
.Y(n_13783)
);

OAI21x1_ASAP7_75t_L g13784 ( 
.A1(n_13289),
.A2(n_1789),
.B(n_1790),
.Y(n_13784)
);

BUFx6f_ASAP7_75t_L g13785 ( 
.A(n_13225),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_12741),
.Y(n_13786)
);

NAND2x1p5_ASAP7_75t_L g13787 ( 
.A(n_13147),
.B(n_1789),
.Y(n_13787)
);

OAI21x1_ASAP7_75t_L g13788 ( 
.A1(n_13001),
.A2(n_1790),
.B(n_1791),
.Y(n_13788)
);

AND2x4_ASAP7_75t_L g13789 ( 
.A(n_13389),
.B(n_1791),
.Y(n_13789)
);

AND2x2_ASAP7_75t_L g13790 ( 
.A(n_13403),
.B(n_1792),
.Y(n_13790)
);

HB1xp67_ASAP7_75t_L g13791 ( 
.A(n_13324),
.Y(n_13791)
);

OAI21x1_ASAP7_75t_L g13792 ( 
.A1(n_13010),
.A2(n_1792),
.B(n_1793),
.Y(n_13792)
);

OAI21x1_ASAP7_75t_SL g13793 ( 
.A1(n_12733),
.A2(n_1793),
.B(n_1794),
.Y(n_13793)
);

OR2x2_ASAP7_75t_L g13794 ( 
.A(n_13406),
.B(n_13316),
.Y(n_13794)
);

INVx1_ASAP7_75t_L g13795 ( 
.A(n_12960),
.Y(n_13795)
);

NAND2x1p5_ASAP7_75t_L g13796 ( 
.A(n_13252),
.B(n_1794),
.Y(n_13796)
);

AND2x2_ASAP7_75t_L g13797 ( 
.A(n_13470),
.B(n_13468),
.Y(n_13797)
);

INVx4_ASAP7_75t_L g13798 ( 
.A(n_13306),
.Y(n_13798)
);

BUFx2_ASAP7_75t_L g13799 ( 
.A(n_13469),
.Y(n_13799)
);

AO21x2_ASAP7_75t_L g13800 ( 
.A1(n_13354),
.A2(n_1795),
.B(n_1796),
.Y(n_13800)
);

INVx6_ASAP7_75t_SL g13801 ( 
.A(n_12825),
.Y(n_13801)
);

CKINVDCx11_ASAP7_75t_R g13802 ( 
.A(n_12908),
.Y(n_13802)
);

OAI21x1_ASAP7_75t_SL g13803 ( 
.A1(n_12970),
.A2(n_1795),
.B(n_1796),
.Y(n_13803)
);

BUFx2_ASAP7_75t_L g13804 ( 
.A(n_13045),
.Y(n_13804)
);

OA21x2_ASAP7_75t_L g13805 ( 
.A1(n_12703),
.A2(n_1797),
.B(n_1798),
.Y(n_13805)
);

BUFx4_ASAP7_75t_SL g13806 ( 
.A(n_13277),
.Y(n_13806)
);

BUFx2_ASAP7_75t_L g13807 ( 
.A(n_13019),
.Y(n_13807)
);

BUFx3_ASAP7_75t_L g13808 ( 
.A(n_13076),
.Y(n_13808)
);

BUFx3_ASAP7_75t_L g13809 ( 
.A(n_13143),
.Y(n_13809)
);

BUFx2_ASAP7_75t_L g13810 ( 
.A(n_13052),
.Y(n_13810)
);

NAND2xp5_ASAP7_75t_L g13811 ( 
.A(n_12748),
.B(n_1797),
.Y(n_13811)
);

AND2x4_ASAP7_75t_L g13812 ( 
.A(n_13056),
.B(n_1798),
.Y(n_13812)
);

BUFx3_ASAP7_75t_L g13813 ( 
.A(n_13211),
.Y(n_13813)
);

BUFx6f_ASAP7_75t_L g13814 ( 
.A(n_13267),
.Y(n_13814)
);

INVx5_ASAP7_75t_L g13815 ( 
.A(n_13186),
.Y(n_13815)
);

INVx3_ASAP7_75t_L g13816 ( 
.A(n_13050),
.Y(n_13816)
);

INVx2_ASAP7_75t_SL g13817 ( 
.A(n_13063),
.Y(n_13817)
);

AOI22x1_ASAP7_75t_L g13818 ( 
.A1(n_12823),
.A2(n_1801),
.B1(n_1799),
.B2(n_1800),
.Y(n_13818)
);

INVx6_ASAP7_75t_L g13819 ( 
.A(n_13285),
.Y(n_13819)
);

NAND2x1p5_ASAP7_75t_L g13820 ( 
.A(n_13266),
.B(n_1799),
.Y(n_13820)
);

AND2x4_ASAP7_75t_L g13821 ( 
.A(n_13291),
.B(n_1800),
.Y(n_13821)
);

NAND2xp5_ASAP7_75t_L g13822 ( 
.A(n_13376),
.B(n_1801),
.Y(n_13822)
);

BUFx2_ASAP7_75t_L g13823 ( 
.A(n_12743),
.Y(n_13823)
);

INVx1_ASAP7_75t_L g13824 ( 
.A(n_12690),
.Y(n_13824)
);

INVx4_ASAP7_75t_L g13825 ( 
.A(n_13235),
.Y(n_13825)
);

BUFx2_ASAP7_75t_L g13826 ( 
.A(n_12744),
.Y(n_13826)
);

OAI21xp5_ASAP7_75t_L g13827 ( 
.A1(n_12898),
.A2(n_1802),
.B(n_1803),
.Y(n_13827)
);

BUFx2_ASAP7_75t_SL g13828 ( 
.A(n_12700),
.Y(n_13828)
);

CKINVDCx20_ASAP7_75t_R g13829 ( 
.A(n_13009),
.Y(n_13829)
);

INVx1_ASAP7_75t_L g13830 ( 
.A(n_12690),
.Y(n_13830)
);

INVx6_ASAP7_75t_L g13831 ( 
.A(n_12716),
.Y(n_13831)
);

OR2x6_ASAP7_75t_L g13832 ( 
.A(n_13447),
.B(n_1802),
.Y(n_13832)
);

AND2x6_ASAP7_75t_L g13833 ( 
.A(n_12793),
.B(n_1803),
.Y(n_13833)
);

INVx1_ASAP7_75t_L g13834 ( 
.A(n_12698),
.Y(n_13834)
);

NAND2x1p5_ASAP7_75t_L g13835 ( 
.A(n_12781),
.B(n_1804),
.Y(n_13835)
);

BUFx6f_ASAP7_75t_L g13836 ( 
.A(n_13465),
.Y(n_13836)
);

INVx1_ASAP7_75t_L g13837 ( 
.A(n_12698),
.Y(n_13837)
);

AO21x2_ASAP7_75t_L g13838 ( 
.A1(n_13361),
.A2(n_1804),
.B(n_1805),
.Y(n_13838)
);

AO21x2_ASAP7_75t_L g13839 ( 
.A1(n_13364),
.A2(n_1805),
.B(n_1806),
.Y(n_13839)
);

INVx3_ASAP7_75t_L g13840 ( 
.A(n_12717),
.Y(n_13840)
);

OAI21x1_ASAP7_75t_L g13841 ( 
.A1(n_13061),
.A2(n_13079),
.B(n_13067),
.Y(n_13841)
);

INVx1_ASAP7_75t_L g13842 ( 
.A(n_12887),
.Y(n_13842)
);

NOR2xp33_ASAP7_75t_L g13843 ( 
.A(n_13345),
.B(n_1807),
.Y(n_13843)
);

AND2x4_ASAP7_75t_L g13844 ( 
.A(n_13390),
.B(n_13236),
.Y(n_13844)
);

INVx3_ASAP7_75t_L g13845 ( 
.A(n_13336),
.Y(n_13845)
);

BUFx6f_ASAP7_75t_L g13846 ( 
.A(n_12943),
.Y(n_13846)
);

BUFx3_ASAP7_75t_L g13847 ( 
.A(n_12936),
.Y(n_13847)
);

OAI21x1_ASAP7_75t_SL g13848 ( 
.A1(n_13435),
.A2(n_1807),
.B(n_1808),
.Y(n_13848)
);

INVx2_ASAP7_75t_SL g13849 ( 
.A(n_12963),
.Y(n_13849)
);

NAND2x1p5_ASAP7_75t_L g13850 ( 
.A(n_12849),
.B(n_1808),
.Y(n_13850)
);

BUFx6f_ASAP7_75t_L g13851 ( 
.A(n_12711),
.Y(n_13851)
);

OAI21x1_ASAP7_75t_L g13852 ( 
.A1(n_13081),
.A2(n_13089),
.B(n_13082),
.Y(n_13852)
);

OAI21x1_ASAP7_75t_L g13853 ( 
.A1(n_13091),
.A2(n_1809),
.B(n_1810),
.Y(n_13853)
);

BUFx6f_ASAP7_75t_L g13854 ( 
.A(n_12812),
.Y(n_13854)
);

CKINVDCx16_ASAP7_75t_R g13855 ( 
.A(n_13123),
.Y(n_13855)
);

CKINVDCx20_ASAP7_75t_R g13856 ( 
.A(n_13398),
.Y(n_13856)
);

NAND2x1p5_ASAP7_75t_L g13857 ( 
.A(n_12835),
.B(n_1809),
.Y(n_13857)
);

OAI21x1_ASAP7_75t_L g13858 ( 
.A1(n_13099),
.A2(n_1810),
.B(n_1811),
.Y(n_13858)
);

INVx1_ASAP7_75t_L g13859 ( 
.A(n_12852),
.Y(n_13859)
);

AOI22x1_ASAP7_75t_L g13860 ( 
.A1(n_13073),
.A2(n_1813),
.B1(n_1811),
.B2(n_1812),
.Y(n_13860)
);

NAND2x1p5_ASAP7_75t_L g13861 ( 
.A(n_12994),
.B(n_1812),
.Y(n_13861)
);

INVx2_ASAP7_75t_SL g13862 ( 
.A(n_12693),
.Y(n_13862)
);

CKINVDCx16_ASAP7_75t_R g13863 ( 
.A(n_13443),
.Y(n_13863)
);

INVx1_ASAP7_75t_SL g13864 ( 
.A(n_13150),
.Y(n_13864)
);

BUFx12f_ASAP7_75t_L g13865 ( 
.A(n_13343),
.Y(n_13865)
);

AO21x2_ASAP7_75t_L g13866 ( 
.A1(n_13393),
.A2(n_1813),
.B(n_1814),
.Y(n_13866)
);

NAND2x1p5_ASAP7_75t_L g13867 ( 
.A(n_12953),
.B(n_13102),
.Y(n_13867)
);

BUFx2_ASAP7_75t_SL g13868 ( 
.A(n_13283),
.Y(n_13868)
);

BUFx2_ASAP7_75t_R g13869 ( 
.A(n_13203),
.Y(n_13869)
);

OAI21x1_ASAP7_75t_L g13870 ( 
.A1(n_12940),
.A2(n_1814),
.B(n_1815),
.Y(n_13870)
);

INVx1_ASAP7_75t_SL g13871 ( 
.A(n_13084),
.Y(n_13871)
);

BUFx12f_ASAP7_75t_L g13872 ( 
.A(n_13450),
.Y(n_13872)
);

BUFx3_ASAP7_75t_L g13873 ( 
.A(n_12763),
.Y(n_13873)
);

OAI21x1_ASAP7_75t_L g13874 ( 
.A1(n_12987),
.A2(n_1815),
.B(n_1816),
.Y(n_13874)
);

BUFx3_ASAP7_75t_L g13875 ( 
.A(n_12782),
.Y(n_13875)
);

INVx1_ASAP7_75t_L g13876 ( 
.A(n_12951),
.Y(n_13876)
);

OAI21x1_ASAP7_75t_SL g13877 ( 
.A1(n_13383),
.A2(n_13188),
.B(n_13124),
.Y(n_13877)
);

BUFx6f_ASAP7_75t_L g13878 ( 
.A(n_13086),
.Y(n_13878)
);

NAND2x1_ASAP7_75t_L g13879 ( 
.A(n_13185),
.B(n_12745),
.Y(n_13879)
);

AO21x2_ASAP7_75t_L g13880 ( 
.A1(n_13404),
.A2(n_1816),
.B(n_1817),
.Y(n_13880)
);

INVx1_ASAP7_75t_SL g13881 ( 
.A(n_13090),
.Y(n_13881)
);

AND2x4_ASAP7_75t_L g13882 ( 
.A(n_13231),
.B(n_1817),
.Y(n_13882)
);

INVx2_ASAP7_75t_L g13883 ( 
.A(n_12701),
.Y(n_13883)
);

OAI21xp5_ASAP7_75t_L g13884 ( 
.A1(n_12901),
.A2(n_1818),
.B(n_1819),
.Y(n_13884)
);

NAND2xp5_ASAP7_75t_L g13885 ( 
.A(n_13047),
.B(n_1818),
.Y(n_13885)
);

CKINVDCx8_ASAP7_75t_R g13886 ( 
.A(n_13215),
.Y(n_13886)
);

BUFx6f_ASAP7_75t_L g13887 ( 
.A(n_13049),
.Y(n_13887)
);

AND2x4_ASAP7_75t_L g13888 ( 
.A(n_13232),
.B(n_1820),
.Y(n_13888)
);

OAI21x1_ASAP7_75t_L g13889 ( 
.A1(n_13016),
.A2(n_1820),
.B(n_1821),
.Y(n_13889)
);

NAND2x1p5_ASAP7_75t_L g13890 ( 
.A(n_13166),
.B(n_13071),
.Y(n_13890)
);

INVx1_ASAP7_75t_L g13891 ( 
.A(n_12955),
.Y(n_13891)
);

AND2x2_ASAP7_75t_L g13892 ( 
.A(n_13457),
.B(n_1821),
.Y(n_13892)
);

INVx2_ASAP7_75t_SL g13893 ( 
.A(n_12734),
.Y(n_13893)
);

CKINVDCx5p33_ASAP7_75t_R g13894 ( 
.A(n_12966),
.Y(n_13894)
);

BUFx2_ASAP7_75t_L g13895 ( 
.A(n_13104),
.Y(n_13895)
);

NAND2xp5_ASAP7_75t_L g13896 ( 
.A(n_13057),
.B(n_1822),
.Y(n_13896)
);

INVx2_ASAP7_75t_L g13897 ( 
.A(n_12984),
.Y(n_13897)
);

INVx1_ASAP7_75t_L g13898 ( 
.A(n_12957),
.Y(n_13898)
);

BUFx3_ASAP7_75t_L g13899 ( 
.A(n_13158),
.Y(n_13899)
);

OAI21x1_ASAP7_75t_L g13900 ( 
.A1(n_13021),
.A2(n_1822),
.B(n_1823),
.Y(n_13900)
);

AND2x6_ASAP7_75t_L g13901 ( 
.A(n_13163),
.B(n_1824),
.Y(n_13901)
);

AO21x2_ASAP7_75t_L g13902 ( 
.A1(n_12787),
.A2(n_1825),
.B(n_1826),
.Y(n_13902)
);

AOI21x1_ASAP7_75t_L g13903 ( 
.A1(n_13338),
.A2(n_1825),
.B(n_1826),
.Y(n_13903)
);

BUFx4f_ASAP7_75t_L g13904 ( 
.A(n_13325),
.Y(n_13904)
);

INVx1_ASAP7_75t_L g13905 ( 
.A(n_12968),
.Y(n_13905)
);

INVx1_ASAP7_75t_SL g13906 ( 
.A(n_13394),
.Y(n_13906)
);

AO21x2_ASAP7_75t_L g13907 ( 
.A1(n_12805),
.A2(n_1827),
.B(n_1828),
.Y(n_13907)
);

INVx1_ASAP7_75t_L g13908 ( 
.A(n_12972),
.Y(n_13908)
);

INVx2_ASAP7_75t_L g13909 ( 
.A(n_12988),
.Y(n_13909)
);

OAI21x1_ASAP7_75t_L g13910 ( 
.A1(n_13030),
.A2(n_1828),
.B(n_1829),
.Y(n_13910)
);

INVx1_ASAP7_75t_L g13911 ( 
.A(n_13007),
.Y(n_13911)
);

BUFx3_ASAP7_75t_L g13912 ( 
.A(n_13395),
.Y(n_13912)
);

NAND2xp5_ASAP7_75t_L g13913 ( 
.A(n_13116),
.B(n_1829),
.Y(n_13913)
);

AO21x2_ASAP7_75t_L g13914 ( 
.A1(n_12897),
.A2(n_12999),
.B(n_12996),
.Y(n_13914)
);

BUFx3_ASAP7_75t_L g13915 ( 
.A(n_13399),
.Y(n_13915)
);

OAI21xp5_ASAP7_75t_L g13916 ( 
.A1(n_12881),
.A2(n_1830),
.B(n_1831),
.Y(n_13916)
);

OAI21x1_ASAP7_75t_L g13917 ( 
.A1(n_12947),
.A2(n_1830),
.B(n_1831),
.Y(n_13917)
);

INVx1_ASAP7_75t_L g13918 ( 
.A(n_13025),
.Y(n_13918)
);

OAI21x1_ASAP7_75t_L g13919 ( 
.A1(n_12981),
.A2(n_1832),
.B(n_1833),
.Y(n_13919)
);

BUFx6f_ASAP7_75t_SL g13920 ( 
.A(n_13205),
.Y(n_13920)
);

OA21x2_ASAP7_75t_L g13921 ( 
.A1(n_13181),
.A2(n_1833),
.B(n_1834),
.Y(n_13921)
);

INVx6_ASAP7_75t_L g13922 ( 
.A(n_13332),
.Y(n_13922)
);

AO21x2_ASAP7_75t_L g13923 ( 
.A1(n_13000),
.A2(n_1834),
.B(n_1835),
.Y(n_13923)
);

NOR2xp33_ASAP7_75t_L g13924 ( 
.A(n_13334),
.B(n_1835),
.Y(n_13924)
);

INVx1_ASAP7_75t_L g13925 ( 
.A(n_12913),
.Y(n_13925)
);

AND2x2_ASAP7_75t_L g13926 ( 
.A(n_13175),
.B(n_1836),
.Y(n_13926)
);

OAI21x1_ASAP7_75t_L g13927 ( 
.A1(n_12986),
.A2(n_1837),
.B(n_1838),
.Y(n_13927)
);

NAND2xp5_ASAP7_75t_L g13928 ( 
.A(n_13168),
.B(n_1837),
.Y(n_13928)
);

HB1xp67_ASAP7_75t_L g13929 ( 
.A(n_12917),
.Y(n_13929)
);

BUFx6f_ASAP7_75t_L g13930 ( 
.A(n_13201),
.Y(n_13930)
);

BUFx6f_ASAP7_75t_L g13931 ( 
.A(n_13417),
.Y(n_13931)
);

OA21x2_ASAP7_75t_L g13932 ( 
.A1(n_12932),
.A2(n_1839),
.B(n_1840),
.Y(n_13932)
);

AO21x2_ASAP7_75t_L g13933 ( 
.A1(n_13005),
.A2(n_1839),
.B(n_1840),
.Y(n_13933)
);

INVx1_ASAP7_75t_L g13934 ( 
.A(n_12925),
.Y(n_13934)
);

NAND2xp5_ASAP7_75t_L g13935 ( 
.A(n_12935),
.B(n_1841),
.Y(n_13935)
);

INVxp67_ASAP7_75t_SL g13936 ( 
.A(n_12941),
.Y(n_13936)
);

BUFx3_ASAP7_75t_L g13937 ( 
.A(n_13421),
.Y(n_13937)
);

INVx1_ASAP7_75t_L g13938 ( 
.A(n_13034),
.Y(n_13938)
);

NAND2xp5_ASAP7_75t_L g13939 ( 
.A(n_12945),
.B(n_1841),
.Y(n_13939)
);

CKINVDCx20_ASAP7_75t_R g13940 ( 
.A(n_13387),
.Y(n_13940)
);

NOR2xp33_ASAP7_75t_L g13941 ( 
.A(n_13342),
.B(n_1842),
.Y(n_13941)
);

INVx1_ASAP7_75t_L g13942 ( 
.A(n_13036),
.Y(n_13942)
);

INVx1_ASAP7_75t_L g13943 ( 
.A(n_13037),
.Y(n_13943)
);

NOR2xp33_ASAP7_75t_L g13944 ( 
.A(n_13349),
.B(n_1843),
.Y(n_13944)
);

INVx1_ASAP7_75t_L g13945 ( 
.A(n_13039),
.Y(n_13945)
);

OAI21x1_ASAP7_75t_L g13946 ( 
.A1(n_13120),
.A2(n_13131),
.B(n_13121),
.Y(n_13946)
);

AO21x2_ASAP7_75t_L g13947 ( 
.A1(n_12798),
.A2(n_1843),
.B(n_1844),
.Y(n_13947)
);

AND2x4_ASAP7_75t_L g13948 ( 
.A(n_13258),
.B(n_1844),
.Y(n_13948)
);

CKINVDCx11_ASAP7_75t_R g13949 ( 
.A(n_13341),
.Y(n_13949)
);

OAI21x1_ASAP7_75t_L g13950 ( 
.A1(n_12993),
.A2(n_1845),
.B(n_1846),
.Y(n_13950)
);

AO21x2_ASAP7_75t_L g13951 ( 
.A1(n_12848),
.A2(n_1845),
.B(n_1846),
.Y(n_13951)
);

NOR2xp33_ASAP7_75t_L g13952 ( 
.A(n_13352),
.B(n_1847),
.Y(n_13952)
);

BUFx2_ASAP7_75t_SL g13953 ( 
.A(n_13242),
.Y(n_13953)
);

NAND2x1p5_ASAP7_75t_L g13954 ( 
.A(n_12919),
.B(n_1847),
.Y(n_13954)
);

AND2x4_ASAP7_75t_L g13955 ( 
.A(n_13269),
.B(n_13276),
.Y(n_13955)
);

INVx1_ASAP7_75t_L g13956 ( 
.A(n_13044),
.Y(n_13956)
);

AND2x2_ASAP7_75t_L g13957 ( 
.A(n_13409),
.B(n_1848),
.Y(n_13957)
);

CKINVDCx6p67_ASAP7_75t_R g13958 ( 
.A(n_13442),
.Y(n_13958)
);

AO21x2_ASAP7_75t_L g13959 ( 
.A1(n_12853),
.A2(n_1848),
.B(n_1849),
.Y(n_13959)
);

AO21x2_ASAP7_75t_L g13960 ( 
.A1(n_12858),
.A2(n_1849),
.B(n_1850),
.Y(n_13960)
);

BUFx2_ASAP7_75t_R g13961 ( 
.A(n_13357),
.Y(n_13961)
);

NAND2x1p5_ASAP7_75t_L g13962 ( 
.A(n_13302),
.B(n_1850),
.Y(n_13962)
);

OAI21x1_ASAP7_75t_L g13963 ( 
.A1(n_12992),
.A2(n_1851),
.B(n_1852),
.Y(n_13963)
);

CKINVDCx11_ASAP7_75t_R g13964 ( 
.A(n_13405),
.Y(n_13964)
);

INVxp67_ASAP7_75t_SL g13965 ( 
.A(n_13054),
.Y(n_13965)
);

INVx6_ASAP7_75t_L g13966 ( 
.A(n_13471),
.Y(n_13966)
);

AO21x2_ASAP7_75t_L g13967 ( 
.A1(n_12869),
.A2(n_1852),
.B(n_1853),
.Y(n_13967)
);

BUFx2_ASAP7_75t_SL g13968 ( 
.A(n_12949),
.Y(n_13968)
);

INVx1_ASAP7_75t_L g13969 ( 
.A(n_13055),
.Y(n_13969)
);

BUFx2_ASAP7_75t_L g13970 ( 
.A(n_13359),
.Y(n_13970)
);

INVx1_ASAP7_75t_L g13971 ( 
.A(n_13065),
.Y(n_13971)
);

OAI21xp5_ASAP7_75t_L g13972 ( 
.A1(n_13184),
.A2(n_1853),
.B(n_1854),
.Y(n_13972)
);

AOI22x1_ASAP7_75t_L g13973 ( 
.A1(n_13256),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.Y(n_13973)
);

INVx4_ASAP7_75t_SL g13974 ( 
.A(n_13453),
.Y(n_13974)
);

BUFx3_ASAP7_75t_L g13975 ( 
.A(n_13446),
.Y(n_13975)
);

NAND2x1p5_ASAP7_75t_L g13976 ( 
.A(n_13344),
.B(n_1855),
.Y(n_13976)
);

INVxp67_ASAP7_75t_SL g13977 ( 
.A(n_13070),
.Y(n_13977)
);

INVx1_ASAP7_75t_SL g13978 ( 
.A(n_13455),
.Y(n_13978)
);

INVx3_ASAP7_75t_SL g13979 ( 
.A(n_13379),
.Y(n_13979)
);

INVx2_ASAP7_75t_SL g13980 ( 
.A(n_13077),
.Y(n_13980)
);

AOI22x1_ASAP7_75t_L g13981 ( 
.A1(n_13268),
.A2(n_1859),
.B1(n_1857),
.B2(n_1858),
.Y(n_13981)
);

BUFx2_ASAP7_75t_SL g13982 ( 
.A(n_13022),
.Y(n_13982)
);

OAI21x1_ASAP7_75t_L g13983 ( 
.A1(n_12820),
.A2(n_1857),
.B(n_1859),
.Y(n_13983)
);

BUFx3_ASAP7_75t_L g13984 ( 
.A(n_13373),
.Y(n_13984)
);

CKINVDCx20_ASAP7_75t_R g13985 ( 
.A(n_13360),
.Y(n_13985)
);

OAI21x1_ASAP7_75t_L g13986 ( 
.A1(n_13053),
.A2(n_1860),
.B(n_1861),
.Y(n_13986)
);

INVx1_ASAP7_75t_L g13987 ( 
.A(n_13122),
.Y(n_13987)
);

BUFx2_ASAP7_75t_L g13988 ( 
.A(n_13366),
.Y(n_13988)
);

INVx1_ASAP7_75t_L g13989 ( 
.A(n_13125),
.Y(n_13989)
);

BUFx12f_ASAP7_75t_L g13990 ( 
.A(n_13279),
.Y(n_13990)
);

AOI22xp33_ASAP7_75t_L g13991 ( 
.A1(n_12800),
.A2(n_1863),
.B1(n_1860),
.B2(n_1862),
.Y(n_13991)
);

BUFx6f_ASAP7_75t_L g13992 ( 
.A(n_13134),
.Y(n_13992)
);

INVx2_ASAP7_75t_L g13993 ( 
.A(n_13148),
.Y(n_13993)
);

INVx2_ASAP7_75t_L g13994 ( 
.A(n_13410),
.Y(n_13994)
);

INVx1_ASAP7_75t_L g13995 ( 
.A(n_12731),
.Y(n_13995)
);

BUFx10_ASAP7_75t_L g13996 ( 
.A(n_13314),
.Y(n_13996)
);

OAI21xp5_ASAP7_75t_L g13997 ( 
.A1(n_13253),
.A2(n_1863),
.B(n_1864),
.Y(n_13997)
);

INVx1_ASAP7_75t_L g13998 ( 
.A(n_12731),
.Y(n_13998)
);

INVx1_ASAP7_75t_SL g13999 ( 
.A(n_13187),
.Y(n_13999)
);

INVx1_ASAP7_75t_L g14000 ( 
.A(n_12720),
.Y(n_14000)
);

OAI21xp5_ASAP7_75t_L g14001 ( 
.A1(n_12754),
.A2(n_1864),
.B(n_1865),
.Y(n_14001)
);

NOR2xp33_ASAP7_75t_L g14002 ( 
.A(n_13362),
.B(n_13367),
.Y(n_14002)
);

AOI21xp5_ASAP7_75t_L g14003 ( 
.A1(n_12811),
.A2(n_1866),
.B(n_1867),
.Y(n_14003)
);

BUFx2_ASAP7_75t_L g14004 ( 
.A(n_13415),
.Y(n_14004)
);

INVx3_ASAP7_75t_L g14005 ( 
.A(n_13419),
.Y(n_14005)
);

INVx1_ASAP7_75t_L g14006 ( 
.A(n_12720),
.Y(n_14006)
);

INVx4_ASAP7_75t_L g14007 ( 
.A(n_12920),
.Y(n_14007)
);

CKINVDCx6p67_ASAP7_75t_R g14008 ( 
.A(n_13369),
.Y(n_14008)
);

OAI21x1_ASAP7_75t_L g14009 ( 
.A1(n_12756),
.A2(n_1866),
.B(n_1867),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_13423),
.Y(n_14010)
);

AOI22x1_ASAP7_75t_L g14011 ( 
.A1(n_13271),
.A2(n_1870),
.B1(n_1868),
.B2(n_1869),
.Y(n_14011)
);

AND2x2_ASAP7_75t_L g14012 ( 
.A(n_13438),
.B(n_1868),
.Y(n_14012)
);

INVx1_ASAP7_75t_SL g14013 ( 
.A(n_13190),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_13448),
.Y(n_14014)
);

BUFx2_ASAP7_75t_L g14015 ( 
.A(n_13460),
.Y(n_14015)
);

BUFx3_ASAP7_75t_L g14016 ( 
.A(n_13206),
.Y(n_14016)
);

BUFx5_ASAP7_75t_L g14017 ( 
.A(n_12819),
.Y(n_14017)
);

INVx4_ASAP7_75t_L g14018 ( 
.A(n_12920),
.Y(n_14018)
);

NOR2xp67_ASAP7_75t_L g14019 ( 
.A(n_13214),
.B(n_1869),
.Y(n_14019)
);

INVx3_ASAP7_75t_L g14020 ( 
.A(n_13466),
.Y(n_14020)
);

INVx2_ASAP7_75t_L g14021 ( 
.A(n_13171),
.Y(n_14021)
);

OAI21x1_ASAP7_75t_L g14022 ( 
.A1(n_13133),
.A2(n_1871),
.B(n_1872),
.Y(n_14022)
);

OAI21x1_ASAP7_75t_L g14023 ( 
.A1(n_13241),
.A2(n_1871),
.B(n_1872),
.Y(n_14023)
);

NOR2x1_ASAP7_75t_R g14024 ( 
.A(n_13182),
.B(n_1873),
.Y(n_14024)
);

OAI21x1_ASAP7_75t_L g14025 ( 
.A1(n_13297),
.A2(n_1873),
.B(n_1875),
.Y(n_14025)
);

AO21x2_ASAP7_75t_L g14026 ( 
.A1(n_13428),
.A2(n_1875),
.B(n_1876),
.Y(n_14026)
);

NAND2x1p5_ASAP7_75t_L g14027 ( 
.A(n_13176),
.B(n_1876),
.Y(n_14027)
);

INVx1_ASAP7_75t_L g14028 ( 
.A(n_12699),
.Y(n_14028)
);

BUFx5_ASAP7_75t_L g14029 ( 
.A(n_13265),
.Y(n_14029)
);

INVx3_ASAP7_75t_L g14030 ( 
.A(n_13340),
.Y(n_14030)
);

BUFx6f_ASAP7_75t_L g14031 ( 
.A(n_13217),
.Y(n_14031)
);

BUFx6f_ASAP7_75t_L g14032 ( 
.A(n_13223),
.Y(n_14032)
);

INVx3_ASAP7_75t_L g14033 ( 
.A(n_13353),
.Y(n_14033)
);

OAI21x1_ASAP7_75t_L g14034 ( 
.A1(n_13391),
.A2(n_1877),
.B(n_1878),
.Y(n_14034)
);

BUFx3_ASAP7_75t_L g14035 ( 
.A(n_13228),
.Y(n_14035)
);

INVxp67_ASAP7_75t_SL g14036 ( 
.A(n_13318),
.Y(n_14036)
);

INVx1_ASAP7_75t_L g14037 ( 
.A(n_12738),
.Y(n_14037)
);

INVx3_ASAP7_75t_L g14038 ( 
.A(n_13328),
.Y(n_14038)
);

HB1xp67_ASAP7_75t_L g14039 ( 
.A(n_12767),
.Y(n_14039)
);

INVx2_ASAP7_75t_SL g14040 ( 
.A(n_13233),
.Y(n_14040)
);

NAND2xp5_ASAP7_75t_L g14041 ( 
.A(n_13237),
.B(n_1877),
.Y(n_14041)
);

BUFx2_ASAP7_75t_L g14042 ( 
.A(n_12767),
.Y(n_14042)
);

AOI22xp33_ASAP7_75t_L g14043 ( 
.A1(n_13441),
.A2(n_1880),
.B1(n_1878),
.B2(n_1879),
.Y(n_14043)
);

AO21x2_ASAP7_75t_L g14044 ( 
.A1(n_13431),
.A2(n_1879),
.B(n_1881),
.Y(n_14044)
);

INVx3_ASAP7_75t_L g14045 ( 
.A(n_13002),
.Y(n_14045)
);

INVx1_ASAP7_75t_L g14046 ( 
.A(n_12738),
.Y(n_14046)
);

INVx1_ASAP7_75t_L g14047 ( 
.A(n_13154),
.Y(n_14047)
);

OAI21x1_ASAP7_75t_L g14048 ( 
.A1(n_13216),
.A2(n_13145),
.B(n_13144),
.Y(n_14048)
);

NAND2xp5_ASAP7_75t_L g14049 ( 
.A(n_13240),
.B(n_1881),
.Y(n_14049)
);

INVxp67_ASAP7_75t_SL g14050 ( 
.A(n_13170),
.Y(n_14050)
);

INVx4_ASAP7_75t_L g14051 ( 
.A(n_13418),
.Y(n_14051)
);

AOI22xp5_ASAP7_75t_SL g14052 ( 
.A1(n_13968),
.A2(n_13351),
.B1(n_13329),
.B2(n_13473),
.Y(n_14052)
);

INVx2_ASAP7_75t_L g14053 ( 
.A(n_13751),
.Y(n_14053)
);

AOI22xp33_ASAP7_75t_L g14054 ( 
.A1(n_13964),
.A2(n_12875),
.B1(n_12892),
.B2(n_13198),
.Y(n_14054)
);

BUFx6f_ASAP7_75t_L g14055 ( 
.A(n_13492),
.Y(n_14055)
);

NOR2xp67_ASAP7_75t_SL g14056 ( 
.A(n_13601),
.B(n_13307),
.Y(n_14056)
);

AND2x2_ASAP7_75t_L g14057 ( 
.A(n_13581),
.B(n_12922),
.Y(n_14057)
);

NAND2xp5_ASAP7_75t_SL g14058 ( 
.A(n_13603),
.B(n_12928),
.Y(n_14058)
);

INVx3_ASAP7_75t_L g14059 ( 
.A(n_13502),
.Y(n_14059)
);

AO21x2_ASAP7_75t_L g14060 ( 
.A1(n_14039),
.A2(n_12841),
.B(n_12822),
.Y(n_14060)
);

OAI21x1_ASAP7_75t_L g14061 ( 
.A1(n_13524),
.A2(n_12724),
.B(n_13356),
.Y(n_14061)
);

OAI21x1_ASAP7_75t_L g14062 ( 
.A1(n_13691),
.A2(n_13411),
.B(n_13226),
.Y(n_14062)
);

INVx1_ASAP7_75t_L g14063 ( 
.A(n_13716),
.Y(n_14063)
);

NOR2xp33_ASAP7_75t_SL g14064 ( 
.A(n_13547),
.B(n_13414),
.Y(n_14064)
);

INVx1_ASAP7_75t_L g14065 ( 
.A(n_13488),
.Y(n_14065)
);

INVx1_ASAP7_75t_L g14066 ( 
.A(n_13500),
.Y(n_14066)
);

AOI22xp5_ASAP7_75t_L g14067 ( 
.A1(n_13729),
.A2(n_13136),
.B1(n_13219),
.B2(n_13445),
.Y(n_14067)
);

OAI221xp5_ASAP7_75t_L g14068 ( 
.A1(n_13694),
.A2(n_12956),
.B1(n_13227),
.B2(n_13221),
.C(n_12883),
.Y(n_14068)
);

OAI21x1_ASAP7_75t_L g14069 ( 
.A1(n_13696),
.A2(n_13229),
.B(n_13224),
.Y(n_14069)
);

NOR2x1_ASAP7_75t_R g14070 ( 
.A(n_13703),
.B(n_13246),
.Y(n_14070)
);

NAND2x1p5_ASAP7_75t_L g14071 ( 
.A(n_13484),
.B(n_13172),
.Y(n_14071)
);

OAI22xp33_ASAP7_75t_L g14072 ( 
.A1(n_14007),
.A2(n_12715),
.B1(n_13127),
.B2(n_13094),
.Y(n_14072)
);

NAND2xp5_ASAP7_75t_L g14073 ( 
.A(n_13659),
.B(n_13257),
.Y(n_14073)
);

OAI21x1_ASAP7_75t_L g14074 ( 
.A1(n_13707),
.A2(n_13230),
.B(n_12964),
.Y(n_14074)
);

INVx1_ASAP7_75t_L g14075 ( 
.A(n_13508),
.Y(n_14075)
);

NAND2xp5_ASAP7_75t_L g14076 ( 
.A(n_13711),
.B(n_13280),
.Y(n_14076)
);

INVx2_ASAP7_75t_L g14077 ( 
.A(n_13751),
.Y(n_14077)
);

BUFx6f_ASAP7_75t_L g14078 ( 
.A(n_13494),
.Y(n_14078)
);

OAI21x1_ASAP7_75t_L g14079 ( 
.A1(n_13879),
.A2(n_13159),
.B(n_13220),
.Y(n_14079)
);

AO31x2_ASAP7_75t_L g14080 ( 
.A1(n_14042),
.A2(n_12888),
.A3(n_13347),
.B(n_12894),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13936),
.B(n_13286),
.Y(n_14081)
);

OAI21x1_ASAP7_75t_L g14082 ( 
.A1(n_13732),
.A2(n_13020),
.B(n_13288),
.Y(n_14082)
);

OAI21xp5_ASAP7_75t_L g14083 ( 
.A1(n_13741),
.A2(n_13028),
.B(n_12746),
.Y(n_14083)
);

AOI22xp33_ASAP7_75t_L g14084 ( 
.A1(n_13901),
.A2(n_13392),
.B1(n_13375),
.B2(n_13132),
.Y(n_14084)
);

NAND2xp5_ASAP7_75t_L g14085 ( 
.A(n_13965),
.B(n_13293),
.Y(n_14085)
);

AND2x2_ASAP7_75t_L g14086 ( 
.A(n_13730),
.B(n_12922),
.Y(n_14086)
);

OAI21x1_ASAP7_75t_L g14087 ( 
.A1(n_13824),
.A2(n_13834),
.B(n_13830),
.Y(n_14087)
);

OAI21x1_ASAP7_75t_L g14088 ( 
.A1(n_13837),
.A2(n_13370),
.B(n_13381),
.Y(n_14088)
);

NAND2xp5_ASAP7_75t_L g14089 ( 
.A(n_13977),
.B(n_13296),
.Y(n_14089)
);

INVxp67_ASAP7_75t_L g14090 ( 
.A(n_13596),
.Y(n_14090)
);

O2A1O1Ixp33_ASAP7_75t_L g14091 ( 
.A1(n_13750),
.A2(n_13684),
.B(n_13877),
.C(n_13598),
.Y(n_14091)
);

BUFx3_ASAP7_75t_L g14092 ( 
.A(n_13700),
.Y(n_14092)
);

CKINVDCx11_ASAP7_75t_R g14093 ( 
.A(n_13557),
.Y(n_14093)
);

BUFx4f_ASAP7_75t_L g14094 ( 
.A(n_13608),
.Y(n_14094)
);

NOR2xp67_ASAP7_75t_L g14095 ( 
.A(n_13601),
.B(n_13304),
.Y(n_14095)
);

INVx2_ASAP7_75t_L g14096 ( 
.A(n_13751),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_13511),
.Y(n_14097)
);

AOI221xp5_ASAP7_75t_L g14098 ( 
.A1(n_13555),
.A2(n_12718),
.B1(n_12729),
.B2(n_13436),
.C(n_13401),
.Y(n_14098)
);

AND2x2_ASAP7_75t_L g14099 ( 
.A(n_13589),
.B(n_13308),
.Y(n_14099)
);

BUFx3_ASAP7_75t_L g14100 ( 
.A(n_13478),
.Y(n_14100)
);

OAI21xp5_ASAP7_75t_L g14101 ( 
.A1(n_13499),
.A2(n_13023),
.B(n_12976),
.Y(n_14101)
);

AO21x2_ASAP7_75t_L g14102 ( 
.A1(n_13859),
.A2(n_12902),
.B(n_13222),
.Y(n_14102)
);

OR2x2_ASAP7_75t_L g14103 ( 
.A(n_13493),
.B(n_13327),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13520),
.Y(n_14104)
);

BUFx12f_ASAP7_75t_L g14105 ( 
.A(n_13534),
.Y(n_14105)
);

AND2x4_ASAP7_75t_L g14106 ( 
.A(n_13546),
.B(n_13358),
.Y(n_14106)
);

OAI21x1_ASAP7_75t_L g14107 ( 
.A1(n_13753),
.A2(n_13386),
.B(n_13014),
.Y(n_14107)
);

AOI21xp5_ASAP7_75t_L g14108 ( 
.A1(n_13523),
.A2(n_13074),
.B(n_13059),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_13528),
.Y(n_14109)
);

NAND2xp5_ASAP7_75t_L g14110 ( 
.A(n_13876),
.B(n_13891),
.Y(n_14110)
);

NAND2xp5_ASAP7_75t_L g14111 ( 
.A(n_13898),
.B(n_13115),
.Y(n_14111)
);

OA21x2_ASAP7_75t_L g14112 ( 
.A1(n_13501),
.A2(n_13335),
.B(n_13140),
.Y(n_14112)
);

NAND2xp5_ASAP7_75t_SL g14113 ( 
.A(n_13742),
.B(n_13174),
.Y(n_14113)
);

INVx2_ASAP7_75t_L g14114 ( 
.A(n_13531),
.Y(n_14114)
);

NAND2xp33_ASAP7_75t_L g14115 ( 
.A(n_13600),
.B(n_13624),
.Y(n_14115)
);

O2A1O1Ixp33_ASAP7_75t_L g14116 ( 
.A1(n_13972),
.A2(n_12774),
.B(n_13195),
.C(n_12954),
.Y(n_14116)
);

OAI21x1_ASAP7_75t_L g14117 ( 
.A1(n_14005),
.A2(n_13003),
.B(n_12778),
.Y(n_14117)
);

AND2x4_ASAP7_75t_L g14118 ( 
.A(n_13580),
.B(n_13072),
.Y(n_14118)
);

AND2x2_ASAP7_75t_L g14119 ( 
.A(n_13563),
.B(n_13397),
.Y(n_14119)
);

INVx1_ASAP7_75t_L g14120 ( 
.A(n_13559),
.Y(n_14120)
);

INVx2_ASAP7_75t_L g14121 ( 
.A(n_13539),
.Y(n_14121)
);

OAI21x1_ASAP7_75t_L g14122 ( 
.A1(n_14020),
.A2(n_12784),
.B(n_12776),
.Y(n_14122)
);

NAND2xp5_ASAP7_75t_L g14123 ( 
.A(n_13905),
.B(n_13908),
.Y(n_14123)
);

AND2x4_ASAP7_75t_L g14124 ( 
.A(n_13485),
.B(n_13521),
.Y(n_14124)
);

OR2x2_ASAP7_75t_L g14125 ( 
.A(n_13675),
.B(n_13072),
.Y(n_14125)
);

INVx2_ASAP7_75t_SL g14126 ( 
.A(n_13495),
.Y(n_14126)
);

OAI21xp5_ASAP7_75t_L g14127 ( 
.A1(n_13811),
.A2(n_13046),
.B(n_13035),
.Y(n_14127)
);

AOI22xp5_ASAP7_75t_L g14128 ( 
.A1(n_13901),
.A2(n_13165),
.B1(n_13424),
.B2(n_12692),
.Y(n_14128)
);

AOI21xp5_ASAP7_75t_L g14129 ( 
.A1(n_13583),
.A2(n_13110),
.B(n_13080),
.Y(n_14129)
);

NAND2x1_ASAP7_75t_L g14130 ( 
.A(n_13577),
.B(n_12975),
.Y(n_14130)
);

OAI21x1_ASAP7_75t_L g14131 ( 
.A1(n_14047),
.A2(n_12786),
.B(n_12785),
.Y(n_14131)
);

NAND2xp5_ASAP7_75t_L g14132 ( 
.A(n_13911),
.B(n_12799),
.Y(n_14132)
);

AOI22xp33_ASAP7_75t_L g14133 ( 
.A1(n_13949),
.A2(n_13152),
.B1(n_13155),
.B2(n_13069),
.Y(n_14133)
);

AO22x2_ASAP7_75t_L g14134 ( 
.A1(n_14018),
.A2(n_14051),
.B1(n_13982),
.B2(n_13868),
.Y(n_14134)
);

BUFx8_ASAP7_75t_L g14135 ( 
.A(n_13920),
.Y(n_14135)
);

OAI21x1_ASAP7_75t_L g14136 ( 
.A1(n_13631),
.A2(n_12808),
.B(n_12788),
.Y(n_14136)
);

AND2x4_ASAP7_75t_L g14137 ( 
.A(n_13676),
.B(n_12799),
.Y(n_14137)
);

NAND2xp5_ASAP7_75t_L g14138 ( 
.A(n_13918),
.B(n_12824),
.Y(n_14138)
);

NAND2x1_ASAP7_75t_L g14139 ( 
.A(n_13725),
.B(n_13434),
.Y(n_14139)
);

NAND2xp5_ASAP7_75t_L g14140 ( 
.A(n_13925),
.B(n_12824),
.Y(n_14140)
);

A2O1A1Ixp33_ASAP7_75t_L g14141 ( 
.A1(n_13529),
.A2(n_12937),
.B(n_12983),
.C(n_12915),
.Y(n_14141)
);

OR2x6_ASAP7_75t_L g14142 ( 
.A(n_13526),
.B(n_13346),
.Y(n_14142)
);

OR2x2_ASAP7_75t_L g14143 ( 
.A(n_13672),
.B(n_12870),
.Y(n_14143)
);

INVx1_ASAP7_75t_L g14144 ( 
.A(n_13562),
.Y(n_14144)
);

BUFx2_ASAP7_75t_L g14145 ( 
.A(n_13574),
.Y(n_14145)
);

AND2x4_ASAP7_75t_L g14146 ( 
.A(n_13514),
.B(n_12870),
.Y(n_14146)
);

AND2x2_ASAP7_75t_L g14147 ( 
.A(n_13626),
.B(n_13397),
.Y(n_14147)
);

BUFx4f_ASAP7_75t_SL g14148 ( 
.A(n_13642),
.Y(n_14148)
);

INVx2_ASAP7_75t_L g14149 ( 
.A(n_13545),
.Y(n_14149)
);

OAI21xp33_ASAP7_75t_L g14150 ( 
.A1(n_13645),
.A2(n_12886),
.B(n_13043),
.Y(n_14150)
);

AND2x2_ASAP7_75t_L g14151 ( 
.A(n_13667),
.B(n_13453),
.Y(n_14151)
);

AND2x4_ASAP7_75t_L g14152 ( 
.A(n_13638),
.B(n_12906),
.Y(n_14152)
);

AOI22xp33_ASAP7_75t_L g14153 ( 
.A1(n_13530),
.A2(n_13118),
.B1(n_13058),
.B2(n_13119),
.Y(n_14153)
);

CKINVDCx20_ASAP7_75t_R g14154 ( 
.A(n_13586),
.Y(n_14154)
);

INVxp67_ASAP7_75t_L g14155 ( 
.A(n_13510),
.Y(n_14155)
);

AO32x2_ASAP7_75t_L g14156 ( 
.A1(n_13862),
.A2(n_12845),
.A3(n_12794),
.B1(n_13103),
.B2(n_13331),
.Y(n_14156)
);

INVx1_ASAP7_75t_SL g14157 ( 
.A(n_13496),
.Y(n_14157)
);

A2O1A1Ixp33_ASAP7_75t_L g14158 ( 
.A1(n_13636),
.A2(n_13292),
.B(n_13412),
.C(n_13408),
.Y(n_14158)
);

INVx8_ASAP7_75t_L g14159 ( 
.A(n_13623),
.Y(n_14159)
);

OAI21x1_ASAP7_75t_L g14160 ( 
.A1(n_14021),
.A2(n_12813),
.B(n_12809),
.Y(n_14160)
);

OAI21x1_ASAP7_75t_L g14161 ( 
.A1(n_13995),
.A2(n_12818),
.B(n_12815),
.Y(n_14161)
);

BUFx6f_ASAP7_75t_L g14162 ( 
.A(n_13505),
.Y(n_14162)
);

AND2x6_ASAP7_75t_L g14163 ( 
.A(n_13836),
.B(n_13161),
.Y(n_14163)
);

AOI22xp5_ASAP7_75t_L g14164 ( 
.A1(n_13489),
.A2(n_13274),
.B1(n_13418),
.B2(n_13275),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_13568),
.Y(n_14165)
);

OAI21x1_ASAP7_75t_SL g14166 ( 
.A1(n_13803),
.A2(n_13449),
.B(n_12834),
.Y(n_14166)
);

OAI21x1_ASAP7_75t_SL g14167 ( 
.A1(n_13793),
.A2(n_13177),
.B(n_13138),
.Y(n_14167)
);

OAI21x1_ASAP7_75t_L g14168 ( 
.A1(n_13998),
.A2(n_12821),
.B(n_13368),
.Y(n_14168)
);

AOI21xp5_ASAP7_75t_L g14169 ( 
.A1(n_14003),
.A2(n_13245),
.B(n_13033),
.Y(n_14169)
);

INVx2_ASAP7_75t_L g14170 ( 
.A(n_13558),
.Y(n_14170)
);

OAI21x1_ASAP7_75t_L g14171 ( 
.A1(n_14000),
.A2(n_13374),
.B(n_13337),
.Y(n_14171)
);

AOI21xp5_ASAP7_75t_L g14172 ( 
.A1(n_13689),
.A2(n_13051),
.B(n_13006),
.Y(n_14172)
);

NAND2xp5_ASAP7_75t_L g14173 ( 
.A(n_13934),
.B(n_12906),
.Y(n_14173)
);

OAI21x1_ASAP7_75t_L g14174 ( 
.A1(n_14006),
.A2(n_13042),
.B(n_13038),
.Y(n_14174)
);

AO21x2_ASAP7_75t_L g14175 ( 
.A1(n_14050),
.A2(n_13194),
.B(n_13164),
.Y(n_14175)
);

NAND2xp5_ASAP7_75t_L g14176 ( 
.A(n_13769),
.B(n_12927),
.Y(n_14176)
);

OAI21x1_ASAP7_75t_L g14177 ( 
.A1(n_13727),
.A2(n_13096),
.B(n_13095),
.Y(n_14177)
);

OAI21x1_ASAP7_75t_L g14178 ( 
.A1(n_13994),
.A2(n_13109),
.B(n_13097),
.Y(n_14178)
);

INVx1_ASAP7_75t_L g14179 ( 
.A(n_13644),
.Y(n_14179)
);

AO21x1_ASAP7_75t_L g14180 ( 
.A1(n_14027),
.A2(n_12872),
.B(n_13243),
.Y(n_14180)
);

BUFx2_ASAP7_75t_L g14181 ( 
.A(n_13509),
.Y(n_14181)
);

INVx1_ASAP7_75t_L g14182 ( 
.A(n_13661),
.Y(n_14182)
);

OAI21x1_ASAP7_75t_L g14183 ( 
.A1(n_14037),
.A2(n_13157),
.B(n_13135),
.Y(n_14183)
);

INVx1_ASAP7_75t_L g14184 ( 
.A(n_13682),
.Y(n_14184)
);

INVxp33_ASAP7_75t_L g14185 ( 
.A(n_13498),
.Y(n_14185)
);

OAI22xp5_ASAP7_75t_L g14186 ( 
.A1(n_13958),
.A2(n_13153),
.B1(n_13075),
.B2(n_12926),
.Y(n_14186)
);

INVx1_ASAP7_75t_L g14187 ( 
.A(n_13686),
.Y(n_14187)
);

INVx2_ASAP7_75t_SL g14188 ( 
.A(n_13481),
.Y(n_14188)
);

OR2x6_ASAP7_75t_L g14189 ( 
.A(n_13612),
.B(n_13309),
.Y(n_14189)
);

OAI21x1_ASAP7_75t_L g14190 ( 
.A1(n_14046),
.A2(n_13193),
.B(n_13167),
.Y(n_14190)
);

OAI21x1_ASAP7_75t_L g14191 ( 
.A1(n_14030),
.A2(n_12773),
.B(n_13197),
.Y(n_14191)
);

OAI21x1_ASAP7_75t_L g14192 ( 
.A1(n_14033),
.A2(n_13212),
.B(n_13209),
.Y(n_14192)
);

BUFx12f_ASAP7_75t_L g14193 ( 
.A(n_13641),
.Y(n_14193)
);

NAND2xp5_ASAP7_75t_L g14194 ( 
.A(n_13772),
.B(n_12927),
.Y(n_14194)
);

AOI21xp5_ASAP7_75t_L g14195 ( 
.A1(n_13916),
.A2(n_13139),
.B(n_13281),
.Y(n_14195)
);

NOR2x1_ASAP7_75t_R g14196 ( 
.A(n_13713),
.B(n_13475),
.Y(n_14196)
);

BUFx2_ASAP7_75t_SL g14197 ( 
.A(n_13815),
.Y(n_14197)
);

OA21x2_ASAP7_75t_L g14198 ( 
.A1(n_13550),
.A2(n_13294),
.B(n_13427),
.Y(n_14198)
);

INVx1_ASAP7_75t_L g14199 ( 
.A(n_13690),
.Y(n_14199)
);

NAND2xp5_ASAP7_75t_L g14200 ( 
.A(n_13776),
.B(n_12930),
.Y(n_14200)
);

OAI21x1_ASAP7_75t_L g14201 ( 
.A1(n_14038),
.A2(n_13301),
.B(n_13298),
.Y(n_14201)
);

OAI22xp33_ASAP7_75t_SL g14202 ( 
.A1(n_13743),
.A2(n_13162),
.B1(n_13413),
.B2(n_13444),
.Y(n_14202)
);

INVx2_ASAP7_75t_L g14203 ( 
.A(n_13525),
.Y(n_14203)
);

INVx1_ASAP7_75t_L g14204 ( 
.A(n_13571),
.Y(n_14204)
);

AO21x2_ASAP7_75t_L g14205 ( 
.A1(n_14010),
.A2(n_13323),
.B(n_13312),
.Y(n_14205)
);

OR2x2_ASAP7_75t_L g14206 ( 
.A(n_13477),
.B(n_13491),
.Y(n_14206)
);

NOR2xp67_ASAP7_75t_L g14207 ( 
.A(n_13742),
.B(n_13295),
.Y(n_14207)
);

OAI22xp5_ASAP7_75t_SL g14208 ( 
.A1(n_13538),
.A2(n_13382),
.B1(n_12985),
.B2(n_13263),
.Y(n_14208)
);

AOI21xp5_ASAP7_75t_L g14209 ( 
.A1(n_14001),
.A2(n_13330),
.B(n_13313),
.Y(n_14209)
);

OA21x2_ASAP7_75t_L g14210 ( 
.A1(n_13970),
.A2(n_13200),
.B(n_12859),
.Y(n_14210)
);

NAND2x1p5_ASAP7_75t_L g14211 ( 
.A(n_13541),
.B(n_13407),
.Y(n_14211)
);

OAI21x1_ASAP7_75t_L g14212 ( 
.A1(n_13841),
.A2(n_13260),
.B(n_13472),
.Y(n_14212)
);

NAND2xp5_ASAP7_75t_SL g14213 ( 
.A(n_13509),
.B(n_12796),
.Y(n_14213)
);

OA21x2_ASAP7_75t_L g14214 ( 
.A1(n_13988),
.A2(n_13430),
.B(n_13142),
.Y(n_14214)
);

OAI21x1_ASAP7_75t_L g14215 ( 
.A1(n_13852),
.A2(n_13299),
.B(n_13008),
.Y(n_14215)
);

CKINVDCx5p33_ASAP7_75t_R g14216 ( 
.A(n_13480),
.Y(n_14216)
);

AND2x4_ASAP7_75t_L g14217 ( 
.A(n_13651),
.B(n_12930),
.Y(n_14217)
);

O2A1O1Ixp33_ASAP7_75t_L g14218 ( 
.A1(n_13832),
.A2(n_13997),
.B(n_13848),
.C(n_13884),
.Y(n_14218)
);

OAI21x1_ASAP7_75t_L g14219 ( 
.A1(n_13946),
.A2(n_13011),
.B(n_12980),
.Y(n_14219)
);

OAI21xp5_ASAP7_75t_L g14220 ( 
.A1(n_13479),
.A2(n_13533),
.B(n_13597),
.Y(n_14220)
);

OAI21x1_ASAP7_75t_L g14221 ( 
.A1(n_14014),
.A2(n_12872),
.B(n_13475),
.Y(n_14221)
);

BUFx2_ASAP7_75t_L g14222 ( 
.A(n_13509),
.Y(n_14222)
);

OA21x2_ASAP7_75t_L g14223 ( 
.A1(n_14004),
.A2(n_14015),
.B(n_13575),
.Y(n_14223)
);

OAI21x1_ASAP7_75t_L g14224 ( 
.A1(n_14045),
.A2(n_12950),
.B(n_12938),
.Y(n_14224)
);

A2O1A1Ixp33_ASAP7_75t_L g14225 ( 
.A1(n_13904),
.A2(n_13213),
.B(n_13310),
.C(n_13305),
.Y(n_14225)
);

AO21x2_ASAP7_75t_L g14226 ( 
.A1(n_13504),
.A2(n_13310),
.B(n_13305),
.Y(n_14226)
);

INVx2_ASAP7_75t_L g14227 ( 
.A(n_13573),
.Y(n_14227)
);

AOI22xp5_ASAP7_75t_L g14228 ( 
.A1(n_14026),
.A2(n_13213),
.B1(n_12950),
.B2(n_12962),
.Y(n_14228)
);

NOR2x1_ASAP7_75t_R g14229 ( 
.A(n_13654),
.B(n_13402),
.Y(n_14229)
);

AO21x2_ASAP7_75t_L g14230 ( 
.A1(n_14028),
.A2(n_13396),
.B(n_13363),
.Y(n_14230)
);

INVx1_ASAP7_75t_L g14231 ( 
.A(n_13593),
.Y(n_14231)
);

OA21x2_ASAP7_75t_L g14232 ( 
.A1(n_13606),
.A2(n_12962),
.B(n_12938),
.Y(n_14232)
);

AOI21xp33_ASAP7_75t_L g14233 ( 
.A1(n_13565),
.A2(n_1882),
.B(n_1883),
.Y(n_14233)
);

AND2x4_ASAP7_75t_L g14234 ( 
.A(n_13616),
.B(n_12971),
.Y(n_14234)
);

OAI21x1_ASAP7_75t_L g14235 ( 
.A1(n_13602),
.A2(n_13018),
.B(n_12971),
.Y(n_14235)
);

NOR2xp67_ASAP7_75t_L g14236 ( 
.A(n_13815),
.B(n_1882),
.Y(n_14236)
);

BUFx8_ASAP7_75t_L g14237 ( 
.A(n_13833),
.Y(n_14237)
);

INVx2_ASAP7_75t_SL g14238 ( 
.A(n_13486),
.Y(n_14238)
);

OAI21x1_ASAP7_75t_L g14239 ( 
.A1(n_14048),
.A2(n_13018),
.B(n_13363),
.Y(n_14239)
);

AND2x4_ASAP7_75t_L g14240 ( 
.A(n_13503),
.B(n_13396),
.Y(n_14240)
);

NAND2xp5_ASAP7_75t_L g14241 ( 
.A(n_13786),
.B(n_13402),
.Y(n_14241)
);

INVx1_ASAP7_75t_L g14242 ( 
.A(n_13614),
.Y(n_14242)
);

INVx3_ASAP7_75t_L g14243 ( 
.A(n_13507),
.Y(n_14243)
);

INVx2_ASAP7_75t_SL g14244 ( 
.A(n_13490),
.Y(n_14244)
);

OAI21x1_ASAP7_75t_L g14245 ( 
.A1(n_14036),
.A2(n_13461),
.B(n_1883),
.Y(n_14245)
);

INVx1_ASAP7_75t_L g14246 ( 
.A(n_13629),
.Y(n_14246)
);

NOR2xp33_ASAP7_75t_L g14247 ( 
.A(n_13671),
.B(n_13748),
.Y(n_14247)
);

NOR2xp33_ASAP7_75t_L g14248 ( 
.A(n_13712),
.B(n_1884),
.Y(n_14248)
);

BUFx3_ASAP7_75t_L g14249 ( 
.A(n_13543),
.Y(n_14249)
);

OAI22xp5_ASAP7_75t_SL g14250 ( 
.A1(n_13855),
.A2(n_13461),
.B1(n_1886),
.B2(n_1884),
.Y(n_14250)
);

OAI21x1_ASAP7_75t_L g14251 ( 
.A1(n_13506),
.A2(n_1885),
.B(n_1886),
.Y(n_14251)
);

AOI21xp5_ASAP7_75t_L g14252 ( 
.A1(n_13827),
.A2(n_1885),
.B(n_1887),
.Y(n_14252)
);

NAND2xp5_ASAP7_75t_L g14253 ( 
.A(n_13929),
.B(n_1887),
.Y(n_14253)
);

OAI21x1_ASAP7_75t_L g14254 ( 
.A1(n_13582),
.A2(n_1888),
.B(n_1889),
.Y(n_14254)
);

OAI21x1_ASAP7_75t_L g14255 ( 
.A1(n_13522),
.A2(n_13745),
.B(n_13549),
.Y(n_14255)
);

INVx2_ASAP7_75t_SL g14256 ( 
.A(n_13518),
.Y(n_14256)
);

NOR2xp67_ASAP7_75t_L g14257 ( 
.A(n_13519),
.B(n_1889),
.Y(n_14257)
);

AOI22xp33_ASAP7_75t_L g14258 ( 
.A1(n_13973),
.A2(n_1892),
.B1(n_1890),
.B2(n_1891),
.Y(n_14258)
);

INVx1_ASAP7_75t_L g14259 ( 
.A(n_13724),
.Y(n_14259)
);

OAI221xp5_ASAP7_75t_SL g14260 ( 
.A1(n_14043),
.A2(n_1892),
.B1(n_1890),
.B2(n_1891),
.C(n_1893),
.Y(n_14260)
);

OAI21x1_ASAP7_75t_L g14261 ( 
.A1(n_13512),
.A2(n_1893),
.B(n_1894),
.Y(n_14261)
);

AND2x4_ASAP7_75t_L g14262 ( 
.A(n_13517),
.B(n_1894),
.Y(n_14262)
);

OAI21x1_ASAP7_75t_L g14263 ( 
.A1(n_13692),
.A2(n_1895),
.B(n_1896),
.Y(n_14263)
);

OAI21xp5_ASAP7_75t_L g14264 ( 
.A1(n_13548),
.A2(n_13843),
.B(n_13552),
.Y(n_14264)
);

NOR2xp67_ASAP7_75t_SL g14265 ( 
.A(n_13655),
.B(n_1895),
.Y(n_14265)
);

INVx1_ASAP7_75t_L g14266 ( 
.A(n_13706),
.Y(n_14266)
);

INVx2_ASAP7_75t_L g14267 ( 
.A(n_13715),
.Y(n_14267)
);

AOI22xp33_ASAP7_75t_L g14268 ( 
.A1(n_13981),
.A2(n_1898),
.B1(n_1896),
.B2(n_1897),
.Y(n_14268)
);

OAI22xp5_ASAP7_75t_SL g14269 ( 
.A1(n_13846),
.A2(n_1900),
.B1(n_1897),
.B2(n_1899),
.Y(n_14269)
);

INVx2_ASAP7_75t_L g14270 ( 
.A(n_13722),
.Y(n_14270)
);

CKINVDCx5p33_ASAP7_75t_R g14271 ( 
.A(n_13633),
.Y(n_14271)
);

OAI21x1_ASAP7_75t_L g14272 ( 
.A1(n_13733),
.A2(n_1899),
.B(n_1900),
.Y(n_14272)
);

AND2x4_ASAP7_75t_L g14273 ( 
.A(n_13537),
.B(n_1901),
.Y(n_14273)
);

OAI21x1_ASAP7_75t_L g14274 ( 
.A1(n_13740),
.A2(n_1902),
.B(n_1903),
.Y(n_14274)
);

OAI21x1_ASAP7_75t_L g14275 ( 
.A1(n_13757),
.A2(n_1902),
.B(n_1904),
.Y(n_14275)
);

OR2x2_ASAP7_75t_L g14276 ( 
.A(n_13483),
.B(n_1904),
.Y(n_14276)
);

INVx2_ASAP7_75t_L g14277 ( 
.A(n_13588),
.Y(n_14277)
);

OAI21x1_ASAP7_75t_L g14278 ( 
.A1(n_13744),
.A2(n_1905),
.B(n_1906),
.Y(n_14278)
);

INVx1_ASAP7_75t_L g14279 ( 
.A(n_13791),
.Y(n_14279)
);

AND2x2_ASAP7_75t_L g14280 ( 
.A(n_13592),
.B(n_1905),
.Y(n_14280)
);

O2A1O1Ixp33_ASAP7_75t_L g14281 ( 
.A1(n_13979),
.A2(n_1908),
.B(n_1906),
.C(n_1907),
.Y(n_14281)
);

INVx2_ASAP7_75t_L g14282 ( 
.A(n_13590),
.Y(n_14282)
);

OAI21x1_ASAP7_75t_L g14283 ( 
.A1(n_13764),
.A2(n_1908),
.B(n_1909),
.Y(n_14283)
);

INVx3_ASAP7_75t_L g14284 ( 
.A(n_13532),
.Y(n_14284)
);

A2O1A1Ixp33_ASAP7_75t_L g14285 ( 
.A1(n_13536),
.A2(n_1911),
.B(n_1909),
.C(n_1910),
.Y(n_14285)
);

INVx1_ASAP7_75t_SL g14286 ( 
.A(n_13677),
.Y(n_14286)
);

NAND2x1p5_ASAP7_75t_L g14287 ( 
.A(n_13799),
.B(n_1911),
.Y(n_14287)
);

CKINVDCx5p33_ASAP7_75t_R g14288 ( 
.A(n_13591),
.Y(n_14288)
);

INVx2_ASAP7_75t_L g14289 ( 
.A(n_13617),
.Y(n_14289)
);

AND2x4_ASAP7_75t_L g14290 ( 
.A(n_13551),
.B(n_1912),
.Y(n_14290)
);

OAI21x1_ASAP7_75t_SL g14291 ( 
.A1(n_13758),
.A2(n_13818),
.B(n_13693),
.Y(n_14291)
);

OAI21x1_ASAP7_75t_L g14292 ( 
.A1(n_13576),
.A2(n_1912),
.B(n_1913),
.Y(n_14292)
);

CKINVDCx5p33_ASAP7_75t_R g14293 ( 
.A(n_13609),
.Y(n_14293)
);

NOR2x1_ASAP7_75t_L g14294 ( 
.A(n_13540),
.B(n_1913),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_13768),
.Y(n_14295)
);

OAI22xp5_ASAP7_75t_L g14296 ( 
.A1(n_13869),
.A2(n_1916),
.B1(n_1914),
.B2(n_1915),
.Y(n_14296)
);

AOI21xp5_ASAP7_75t_L g14297 ( 
.A1(n_13739),
.A2(n_1914),
.B(n_1915),
.Y(n_14297)
);

OAI21x1_ASAP7_75t_SL g14298 ( 
.A1(n_13738),
.A2(n_1916),
.B(n_1917),
.Y(n_14298)
);

AND2x2_ASAP7_75t_L g14299 ( 
.A(n_13845),
.B(n_1917),
.Y(n_14299)
);

AOI21xp33_ASAP7_75t_SL g14300 ( 
.A1(n_13542),
.A2(n_1918),
.B(n_1919),
.Y(n_14300)
);

INVx2_ASAP7_75t_L g14301 ( 
.A(n_13630),
.Y(n_14301)
);

BUFx3_ASAP7_75t_L g14302 ( 
.A(n_13487),
.Y(n_14302)
);

OAI22xp33_ASAP7_75t_L g14303 ( 
.A1(n_13846),
.A2(n_1920),
.B1(n_1918),
.B2(n_1919),
.Y(n_14303)
);

OA21x2_ASAP7_75t_L g14304 ( 
.A1(n_13657),
.A2(n_1920),
.B(n_1921),
.Y(n_14304)
);

CKINVDCx5p33_ASAP7_75t_R g14305 ( 
.A(n_13625),
.Y(n_14305)
);

INVx2_ASAP7_75t_L g14306 ( 
.A(n_13647),
.Y(n_14306)
);

OAI21x1_ASAP7_75t_L g14307 ( 
.A1(n_13569),
.A2(n_1922),
.B(n_1923),
.Y(n_14307)
);

BUFx6f_ASAP7_75t_L g14308 ( 
.A(n_13476),
.Y(n_14308)
);

OAI21x1_ASAP7_75t_L g14309 ( 
.A1(n_13567),
.A2(n_1923),
.B(n_1924),
.Y(n_14309)
);

AOI22xp33_ASAP7_75t_SL g14310 ( 
.A1(n_13604),
.A2(n_1926),
.B1(n_1924),
.B2(n_1925),
.Y(n_14310)
);

AO31x2_ASAP7_75t_L g14311 ( 
.A1(n_13938),
.A2(n_1927),
.A3(n_1925),
.B(n_1926),
.Y(n_14311)
);

AO21x2_ASAP7_75t_L g14312 ( 
.A1(n_13660),
.A2(n_1927),
.B(n_1928),
.Y(n_14312)
);

INVx2_ASAP7_75t_L g14313 ( 
.A(n_13663),
.Y(n_14313)
);

OAI21xp5_ASAP7_75t_L g14314 ( 
.A1(n_13618),
.A2(n_1928),
.B(n_1929),
.Y(n_14314)
);

HB1xp67_ASAP7_75t_L g14315 ( 
.A(n_13607),
.Y(n_14315)
);

AOI22xp33_ASAP7_75t_L g14316 ( 
.A1(n_14011),
.A2(n_1931),
.B1(n_1929),
.B2(n_1930),
.Y(n_14316)
);

NAND2x1p5_ASAP7_75t_L g14317 ( 
.A(n_13566),
.B(n_1931),
.Y(n_14317)
);

NOR2xp33_ASAP7_75t_SL g14318 ( 
.A(n_13961),
.B(n_1932),
.Y(n_14318)
);

NOR2xp33_ASAP7_75t_L g14319 ( 
.A(n_13942),
.B(n_1932),
.Y(n_14319)
);

AO21x2_ASAP7_75t_L g14320 ( 
.A1(n_13622),
.A2(n_1933),
.B(n_1934),
.Y(n_14320)
);

OAI22xp33_ASAP7_75t_L g14321 ( 
.A1(n_13863),
.A2(n_1935),
.B1(n_1933),
.B2(n_1934),
.Y(n_14321)
);

NAND2xp33_ASAP7_75t_SL g14322 ( 
.A(n_13836),
.B(n_1935),
.Y(n_14322)
);

O2A1O1Ixp5_ASAP7_75t_L g14323 ( 
.A1(n_13955),
.A2(n_13844),
.B(n_13731),
.C(n_13762),
.Y(n_14323)
);

AND2x2_ASAP7_75t_L g14324 ( 
.A(n_13816),
.B(n_1936),
.Y(n_14324)
);

OAI21xp5_ASAP7_75t_L g14325 ( 
.A1(n_13628),
.A2(n_1936),
.B(n_1937),
.Y(n_14325)
);

OAI21x1_ASAP7_75t_L g14326 ( 
.A1(n_13794),
.A2(n_1937),
.B(n_1938),
.Y(n_14326)
);

AND2x4_ASAP7_75t_L g14327 ( 
.A(n_13797),
.B(n_1939),
.Y(n_14327)
);

O2A1O1Ixp33_ASAP7_75t_L g14328 ( 
.A1(n_13890),
.A2(n_1941),
.B(n_1939),
.C(n_1940),
.Y(n_14328)
);

BUFx2_ASAP7_75t_L g14329 ( 
.A(n_13895),
.Y(n_14329)
);

INVx2_ASAP7_75t_L g14330 ( 
.A(n_13680),
.Y(n_14330)
);

OAI21x1_ASAP7_75t_L g14331 ( 
.A1(n_13560),
.A2(n_1940),
.B(n_1942),
.Y(n_14331)
);

NAND2xp5_ASAP7_75t_L g14332 ( 
.A(n_13943),
.B(n_1942),
.Y(n_14332)
);

NAND2xp5_ASAP7_75t_L g14333 ( 
.A(n_13945),
.B(n_1943),
.Y(n_14333)
);

OAI21x1_ASAP7_75t_L g14334 ( 
.A1(n_13572),
.A2(n_13909),
.B(n_13897),
.Y(n_14334)
);

INVx1_ASAP7_75t_L g14335 ( 
.A(n_13635),
.Y(n_14335)
);

OA21x2_ASAP7_75t_L g14336 ( 
.A1(n_13956),
.A2(n_1943),
.B(n_1944),
.Y(n_14336)
);

OAI21x1_ASAP7_75t_L g14337 ( 
.A1(n_13993),
.A2(n_13595),
.B(n_13735),
.Y(n_14337)
);

AOI21xp5_ASAP7_75t_L g14338 ( 
.A1(n_13947),
.A2(n_13959),
.B(n_13951),
.Y(n_14338)
);

INVx3_ASAP7_75t_L g14339 ( 
.A(n_13620),
.Y(n_14339)
);

OAI21x1_ASAP7_75t_L g14340 ( 
.A1(n_13554),
.A2(n_1944),
.B(n_1945),
.Y(n_14340)
);

BUFx4_ASAP7_75t_R g14341 ( 
.A(n_13996),
.Y(n_14341)
);

BUFx2_ASAP7_75t_L g14342 ( 
.A(n_13515),
.Y(n_14342)
);

BUFx2_ASAP7_75t_R g14343 ( 
.A(n_13886),
.Y(n_14343)
);

NAND2xp5_ASAP7_75t_L g14344 ( 
.A(n_13969),
.B(n_1945),
.Y(n_14344)
);

OAI21x1_ASAP7_75t_L g14345 ( 
.A1(n_13621),
.A2(n_1946),
.B(n_1947),
.Y(n_14345)
);

OAI22xp5_ASAP7_75t_L g14346 ( 
.A1(n_13991),
.A2(n_1948),
.B1(n_1946),
.B2(n_1947),
.Y(n_14346)
);

OAI21x1_ASAP7_75t_L g14347 ( 
.A1(n_13650),
.A2(n_1948),
.B(n_1949),
.Y(n_14347)
);

BUFx2_ASAP7_75t_L g14348 ( 
.A(n_13515),
.Y(n_14348)
);

NAND2xp5_ASAP7_75t_L g14349 ( 
.A(n_13971),
.B(n_1950),
.Y(n_14349)
);

OAI21x1_ASAP7_75t_L g14350 ( 
.A1(n_13883),
.A2(n_13718),
.B(n_13695),
.Y(n_14350)
);

OAI21x1_ASAP7_75t_SL g14351 ( 
.A1(n_13658),
.A2(n_1951),
.B(n_1952),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_13665),
.Y(n_14352)
);

INVx1_ASAP7_75t_L g14353 ( 
.A(n_13678),
.Y(n_14353)
);

INVx3_ASAP7_75t_L g14354 ( 
.A(n_13643),
.Y(n_14354)
);

NOR2x1_ASAP7_75t_SL g14355 ( 
.A(n_13828),
.B(n_1951),
.Y(n_14355)
);

INVx3_ASAP7_75t_L g14356 ( 
.A(n_13648),
.Y(n_14356)
);

INVx3_ASAP7_75t_L g14357 ( 
.A(n_13688),
.Y(n_14357)
);

OR3x4_ASAP7_75t_SL g14358 ( 
.A(n_13806),
.B(n_13579),
.C(n_13760),
.Y(n_14358)
);

O2A1O1Ixp5_ASAP7_75t_L g14359 ( 
.A1(n_13987),
.A2(n_1954),
.B(n_1952),
.C(n_1953),
.Y(n_14359)
);

OR2x2_ASAP7_75t_L g14360 ( 
.A(n_13752),
.B(n_1953),
.Y(n_14360)
);

INVxp67_ASAP7_75t_SL g14361 ( 
.A(n_14031),
.Y(n_14361)
);

AOI22xp33_ASAP7_75t_L g14362 ( 
.A1(n_14044),
.A2(n_1957),
.B1(n_1955),
.B2(n_1956),
.Y(n_14362)
);

OAI21x1_ASAP7_75t_L g14363 ( 
.A1(n_13989),
.A2(n_1955),
.B(n_1956),
.Y(n_14363)
);

HB1xp67_ASAP7_75t_L g14364 ( 
.A(n_13781),
.Y(n_14364)
);

INVx1_ASAP7_75t_L g14365 ( 
.A(n_13754),
.Y(n_14365)
);

OAI22xp5_ASAP7_75t_L g14366 ( 
.A1(n_13922),
.A2(n_13953),
.B1(n_13544),
.B2(n_13857),
.Y(n_14366)
);

OAI21x1_ASAP7_75t_L g14367 ( 
.A1(n_13709),
.A2(n_1958),
.B(n_1959),
.Y(n_14367)
);

INVx1_ASAP7_75t_L g14368 ( 
.A(n_13795),
.Y(n_14368)
);

AOI21xp5_ASAP7_75t_L g14369 ( 
.A1(n_13960),
.A2(n_1958),
.B(n_1959),
.Y(n_14369)
);

AO21x2_ASAP7_75t_L g14370 ( 
.A1(n_14019),
.A2(n_1960),
.B(n_1961),
.Y(n_14370)
);

OA21x2_ASAP7_75t_L g14371 ( 
.A1(n_13807),
.A2(n_1960),
.B(n_1962),
.Y(n_14371)
);

INVx3_ASAP7_75t_L g14372 ( 
.A(n_13688),
.Y(n_14372)
);

AOI21xp33_ASAP7_75t_L g14373 ( 
.A1(n_14024),
.A2(n_1962),
.B(n_1963),
.Y(n_14373)
);

OAI21xp33_ASAP7_75t_SL g14374 ( 
.A1(n_13893),
.A2(n_1963),
.B(n_1965),
.Y(n_14374)
);

NOR2xp67_ASAP7_75t_L g14375 ( 
.A(n_13980),
.B(n_1965),
.Y(n_14375)
);

OR2x2_ASAP7_75t_L g14376 ( 
.A(n_13771),
.B(n_1966),
.Y(n_14376)
);

BUFx3_ASAP7_75t_L g14377 ( 
.A(n_13669),
.Y(n_14377)
);

INVx1_ASAP7_75t_SL g14378 ( 
.A(n_13770),
.Y(n_14378)
);

OAI21x1_ASAP7_75t_L g14379 ( 
.A1(n_13784),
.A2(n_1966),
.B(n_1967),
.Y(n_14379)
);

OAI21x1_ASAP7_75t_L g14380 ( 
.A1(n_13653),
.A2(n_1967),
.B(n_1969),
.Y(n_14380)
);

AND2x4_ASAP7_75t_L g14381 ( 
.A(n_13763),
.B(n_1969),
.Y(n_14381)
);

AOI22xp33_ASAP7_75t_L g14382 ( 
.A1(n_13967),
.A2(n_1972),
.B1(n_1970),
.B2(n_1971),
.Y(n_14382)
);

INVx1_ASAP7_75t_L g14383 ( 
.A(n_13842),
.Y(n_14383)
);

BUFx3_ASAP7_75t_L g14384 ( 
.A(n_13673),
.Y(n_14384)
);

INVx2_ASAP7_75t_L g14385 ( 
.A(n_13779),
.Y(n_14385)
);

CKINVDCx5p33_ASAP7_75t_R g14386 ( 
.A(n_13553),
.Y(n_14386)
);

OAI21x1_ASAP7_75t_L g14387 ( 
.A1(n_13666),
.A2(n_1970),
.B(n_1971),
.Y(n_14387)
);

INVx2_ASAP7_75t_SL g14388 ( 
.A(n_13611),
.Y(n_14388)
);

INVx1_ASAP7_75t_L g14389 ( 
.A(n_13701),
.Y(n_14389)
);

NAND2xp5_ASAP7_75t_L g14390 ( 
.A(n_13864),
.B(n_1972),
.Y(n_14390)
);

BUFx3_ASAP7_75t_L g14391 ( 
.A(n_13585),
.Y(n_14391)
);

INVx1_ASAP7_75t_L g14392 ( 
.A(n_13679),
.Y(n_14392)
);

INVxp67_ASAP7_75t_L g14393 ( 
.A(n_13516),
.Y(n_14393)
);

O2A1O1Ixp33_ASAP7_75t_SL g14394 ( 
.A1(n_13885),
.A2(n_1975),
.B(n_1973),
.C(n_1974),
.Y(n_14394)
);

AO21x1_ASAP7_75t_L g14395 ( 
.A1(n_13708),
.A2(n_14002),
.B(n_13825),
.Y(n_14395)
);

AND2x4_ASAP7_75t_L g14396 ( 
.A(n_13723),
.B(n_1974),
.Y(n_14396)
);

OAI21x1_ASAP7_75t_L g14397 ( 
.A1(n_13674),
.A2(n_1975),
.B(n_1976),
.Y(n_14397)
);

CKINVDCx6p67_ASAP7_75t_R g14398 ( 
.A(n_13833),
.Y(n_14398)
);

INVx2_ASAP7_75t_L g14399 ( 
.A(n_13515),
.Y(n_14399)
);

INVx2_ASAP7_75t_L g14400 ( 
.A(n_13804),
.Y(n_14400)
);

BUFx2_ASAP7_75t_L g14401 ( 
.A(n_13584),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_13823),
.Y(n_14402)
);

BUFx2_ASAP7_75t_L g14403 ( 
.A(n_13605),
.Y(n_14403)
);

INVx1_ASAP7_75t_L g14404 ( 
.A(n_13826),
.Y(n_14404)
);

AOI22xp33_ASAP7_75t_L g14405 ( 
.A1(n_13800),
.A2(n_13839),
.B1(n_13866),
.B2(n_13838),
.Y(n_14405)
);

INVx2_ASAP7_75t_L g14406 ( 
.A(n_13808),
.Y(n_14406)
);

OR2x2_ASAP7_75t_L g14407 ( 
.A(n_13871),
.B(n_1977),
.Y(n_14407)
);

BUFx2_ASAP7_75t_L g14408 ( 
.A(n_13810),
.Y(n_14408)
);

OAI21x1_ASAP7_75t_SL g14409 ( 
.A1(n_13849),
.A2(n_1977),
.B(n_1978),
.Y(n_14409)
);

OAI21x1_ASAP7_75t_L g14410 ( 
.A1(n_13714),
.A2(n_1979),
.B(n_1980),
.Y(n_14410)
);

AOI21x1_ASAP7_75t_L g14411 ( 
.A1(n_13683),
.A2(n_1979),
.B(n_1980),
.Y(n_14411)
);

OAI221xp5_ASAP7_75t_SL g14412 ( 
.A1(n_13896),
.A2(n_1983),
.B1(n_1981),
.B2(n_1982),
.C(n_1984),
.Y(n_14412)
);

OAI21x1_ASAP7_75t_L g14413 ( 
.A1(n_13720),
.A2(n_1981),
.B(n_1982),
.Y(n_14413)
);

OR3x4_ASAP7_75t_SL g14414 ( 
.A(n_14008),
.B(n_1983),
.C(n_1984),
.Y(n_14414)
);

HB1xp67_ASAP7_75t_L g14415 ( 
.A(n_14040),
.Y(n_14415)
);

OAI21x1_ASAP7_75t_SL g14416 ( 
.A1(n_13527),
.A2(n_1985),
.B(n_1986),
.Y(n_14416)
);

AND2x2_ASAP7_75t_L g14417 ( 
.A(n_13599),
.B(n_1987),
.Y(n_14417)
);

BUFx2_ASAP7_75t_L g14418 ( 
.A(n_13756),
.Y(n_14418)
);

AOI21xp5_ASAP7_75t_L g14419 ( 
.A1(n_13759),
.A2(n_1988),
.B(n_1989),
.Y(n_14419)
);

OA21x2_ASAP7_75t_L g14420 ( 
.A1(n_14025),
.A2(n_1988),
.B(n_1990),
.Y(n_14420)
);

HB1xp67_ASAP7_75t_L g14421 ( 
.A(n_13881),
.Y(n_14421)
);

NAND2xp33_ASAP7_75t_SL g14422 ( 
.A(n_13887),
.B(n_1990),
.Y(n_14422)
);

OAI21x1_ASAP7_75t_L g14423 ( 
.A1(n_13728),
.A2(n_1991),
.B(n_1992),
.Y(n_14423)
);

OAI21x1_ASAP7_75t_L g14424 ( 
.A1(n_13726),
.A2(n_13747),
.B(n_14034),
.Y(n_14424)
);

OAI21x1_ASAP7_75t_L g14425 ( 
.A1(n_14022),
.A2(n_1991),
.B(n_1992),
.Y(n_14425)
);

OR2x2_ASAP7_75t_L g14426 ( 
.A(n_13906),
.B(n_1993),
.Y(n_14426)
);

OAI21x1_ASAP7_75t_L g14427 ( 
.A1(n_13761),
.A2(n_1993),
.B(n_1994),
.Y(n_14427)
);

NOR2x1p5_ASAP7_75t_L g14428 ( 
.A(n_13851),
.B(n_1995),
.Y(n_14428)
);

NOR2x1_ASAP7_75t_L g14429 ( 
.A(n_13899),
.B(n_1996),
.Y(n_14429)
);

AOI22xp33_ASAP7_75t_L g14430 ( 
.A1(n_13990),
.A2(n_1998),
.B1(n_1996),
.B2(n_1997),
.Y(n_14430)
);

OAI22xp5_ASAP7_75t_L g14431 ( 
.A1(n_13867),
.A2(n_1999),
.B1(n_1997),
.B2(n_1998),
.Y(n_14431)
);

INVx2_ASAP7_75t_L g14432 ( 
.A(n_13809),
.Y(n_14432)
);

OAI21x1_ASAP7_75t_L g14433 ( 
.A1(n_13765),
.A2(n_1999),
.B(n_2001),
.Y(n_14433)
);

AND2x2_ASAP7_75t_L g14434 ( 
.A(n_13840),
.B(n_2001),
.Y(n_14434)
);

OR2x2_ASAP7_75t_L g14435 ( 
.A(n_13978),
.B(n_2002),
.Y(n_14435)
);

INVx5_ASAP7_75t_L g14436 ( 
.A(n_13930),
.Y(n_14436)
);

BUFx2_ASAP7_75t_R g14437 ( 
.A(n_13704),
.Y(n_14437)
);

OA21x2_ASAP7_75t_L g14438 ( 
.A1(n_13822),
.A2(n_2003),
.B(n_2004),
.Y(n_14438)
);

INVx1_ASAP7_75t_L g14439 ( 
.A(n_13974),
.Y(n_14439)
);

OAI21x1_ASAP7_75t_L g14440 ( 
.A1(n_13767),
.A2(n_2003),
.B(n_2004),
.Y(n_14440)
);

NAND2x1p5_ASAP7_75t_L g14441 ( 
.A(n_13737),
.B(n_2005),
.Y(n_14441)
);

AO21x2_ASAP7_75t_L g14442 ( 
.A1(n_13907),
.A2(n_2005),
.B(n_2006),
.Y(n_14442)
);

AO21x1_ASAP7_75t_L g14443 ( 
.A1(n_13702),
.A2(n_2006),
.B(n_2007),
.Y(n_14443)
);

AOI21xp5_ASAP7_75t_L g14444 ( 
.A1(n_13914),
.A2(n_13556),
.B(n_13880),
.Y(n_14444)
);

AO21x2_ASAP7_75t_L g14445 ( 
.A1(n_13664),
.A2(n_2007),
.B(n_2008),
.Y(n_14445)
);

INVx2_ASAP7_75t_L g14446 ( 
.A(n_13813),
.Y(n_14446)
);

OAI21x1_ASAP7_75t_L g14447 ( 
.A1(n_13773),
.A2(n_2008),
.B(n_2009),
.Y(n_14447)
);

BUFx6f_ASAP7_75t_L g14448 ( 
.A(n_13482),
.Y(n_14448)
);

OAI21x1_ASAP7_75t_L g14449 ( 
.A1(n_13774),
.A2(n_2010),
.B(n_2011),
.Y(n_14449)
);

INVx1_ASAP7_75t_L g14450 ( 
.A(n_13649),
.Y(n_14450)
);

BUFx2_ASAP7_75t_L g14451 ( 
.A(n_13847),
.Y(n_14451)
);

OAI221xp5_ASAP7_75t_L g14452 ( 
.A1(n_13850),
.A2(n_2012),
.B1(n_2010),
.B2(n_2011),
.C(n_2013),
.Y(n_14452)
);

OAI22xp33_ASAP7_75t_SL g14453 ( 
.A1(n_13831),
.A2(n_2014),
.B1(n_2012),
.B2(n_2013),
.Y(n_14453)
);

OAI21x1_ASAP7_75t_L g14454 ( 
.A1(n_13783),
.A2(n_2014),
.B(n_2015),
.Y(n_14454)
);

INVx6_ASAP7_75t_L g14455 ( 
.A(n_13685),
.Y(n_14455)
);

INVx1_ASAP7_75t_L g14456 ( 
.A(n_13780),
.Y(n_14456)
);

OAI221xp5_ASAP7_75t_L g14457 ( 
.A1(n_13924),
.A2(n_2017),
.B1(n_2015),
.B2(n_2016),
.C(n_2018),
.Y(n_14457)
);

NAND2xp5_ASAP7_75t_L g14458 ( 
.A(n_13999),
.B(n_14013),
.Y(n_14458)
);

OAI21x1_ASAP7_75t_L g14459 ( 
.A1(n_13788),
.A2(n_2016),
.B(n_2017),
.Y(n_14459)
);

AND2x2_ASAP7_75t_L g14460 ( 
.A(n_13578),
.B(n_2018),
.Y(n_14460)
);

OAI21x1_ASAP7_75t_L g14461 ( 
.A1(n_13792),
.A2(n_2019),
.B(n_2020),
.Y(n_14461)
);

AOI22xp33_ASAP7_75t_L g14462 ( 
.A1(n_14031),
.A2(n_2021),
.B1(n_2019),
.B2(n_2020),
.Y(n_14462)
);

INVx1_ASAP7_75t_L g14463 ( 
.A(n_13805),
.Y(n_14463)
);

AOI22xp5_ASAP7_75t_L g14464 ( 
.A1(n_13594),
.A2(n_2024),
.B1(n_2022),
.B2(n_2023),
.Y(n_14464)
);

INVxp67_ASAP7_75t_L g14465 ( 
.A(n_13610),
.Y(n_14465)
);

INVx1_ASAP7_75t_L g14466 ( 
.A(n_13932),
.Y(n_14466)
);

OR2x2_ASAP7_75t_SL g14467 ( 
.A(n_13930),
.B(n_2023),
.Y(n_14467)
);

AO21x1_ASAP7_75t_L g14468 ( 
.A1(n_13535),
.A2(n_2025),
.B(n_2026),
.Y(n_14468)
);

INVx2_ASAP7_75t_L g14469 ( 
.A(n_13817),
.Y(n_14469)
);

OR2x6_ASAP7_75t_L g14470 ( 
.A(n_13637),
.B(n_2026),
.Y(n_14470)
);

INVx1_ASAP7_75t_L g14471 ( 
.A(n_13790),
.Y(n_14471)
);

INVx8_ASAP7_75t_L g14472 ( 
.A(n_13587),
.Y(n_14472)
);

AOI21x1_ASAP7_75t_L g14473 ( 
.A1(n_13935),
.A2(n_2027),
.B(n_2028),
.Y(n_14473)
);

HB1xp67_ASAP7_75t_L g14474 ( 
.A(n_13992),
.Y(n_14474)
);

OAI22xp5_ASAP7_75t_L g14475 ( 
.A1(n_13749),
.A2(n_2029),
.B1(n_2027),
.B2(n_2028),
.Y(n_14475)
);

NAND2x1p5_ASAP7_75t_L g14476 ( 
.A(n_13710),
.B(n_2029),
.Y(n_14476)
);

OA21x2_ASAP7_75t_L g14477 ( 
.A1(n_13939),
.A2(n_2030),
.B(n_2031),
.Y(n_14477)
);

OAI21x1_ASAP7_75t_L g14478 ( 
.A1(n_13853),
.A2(n_2030),
.B(n_2031),
.Y(n_14478)
);

CKINVDCx20_ASAP7_75t_R g14479 ( 
.A(n_13856),
.Y(n_14479)
);

OAI21x1_ASAP7_75t_L g14480 ( 
.A1(n_13858),
.A2(n_2032),
.B(n_2033),
.Y(n_14480)
);

OAI22xp5_ASAP7_75t_L g14481 ( 
.A1(n_13787),
.A2(n_2034),
.B1(n_2032),
.B2(n_2033),
.Y(n_14481)
);

AND2x4_ASAP7_75t_L g14482 ( 
.A(n_13755),
.B(n_2035),
.Y(n_14482)
);

CKINVDCx16_ASAP7_75t_R g14483 ( 
.A(n_13865),
.Y(n_14483)
);

OA21x2_ASAP7_75t_L g14484 ( 
.A1(n_13913),
.A2(n_2035),
.B(n_2036),
.Y(n_14484)
);

OAI22xp33_ASAP7_75t_L g14485 ( 
.A1(n_13887),
.A2(n_2038),
.B1(n_2036),
.B2(n_2037),
.Y(n_14485)
);

AO22x2_ASAP7_75t_L g14486 ( 
.A1(n_13798),
.A2(n_2039),
.B1(n_2037),
.B2(n_2038),
.Y(n_14486)
);

INVx2_ASAP7_75t_L g14487 ( 
.A(n_14032),
.Y(n_14487)
);

OA21x2_ASAP7_75t_L g14488 ( 
.A1(n_14041),
.A2(n_2040),
.B(n_2041),
.Y(n_14488)
);

NAND2x1p5_ASAP7_75t_L g14489 ( 
.A(n_13851),
.B(n_2041),
.Y(n_14489)
);

AO21x2_ASAP7_75t_L g14490 ( 
.A1(n_13928),
.A2(n_2042),
.B(n_2043),
.Y(n_14490)
);

OAI21x1_ASAP7_75t_L g14491 ( 
.A1(n_13870),
.A2(n_2042),
.B(n_2043),
.Y(n_14491)
);

OR2x2_ASAP7_75t_L g14492 ( 
.A(n_13912),
.B(n_2044),
.Y(n_14492)
);

OR2x2_ASAP7_75t_L g14493 ( 
.A(n_13915),
.B(n_2045),
.Y(n_14493)
);

AOI22xp33_ASAP7_75t_L g14494 ( 
.A1(n_14032),
.A2(n_2047),
.B1(n_2045),
.B2(n_2046),
.Y(n_14494)
);

AOI22xp33_ASAP7_75t_L g14495 ( 
.A1(n_14017),
.A2(n_2048),
.B1(n_2046),
.B2(n_2047),
.Y(n_14495)
);

NAND2xp5_ASAP7_75t_L g14496 ( 
.A(n_13992),
.B(n_2048),
.Y(n_14496)
);

BUFx4_ASAP7_75t_SL g14497 ( 
.A(n_13639),
.Y(n_14497)
);

NAND2xp5_ASAP7_75t_L g14498 ( 
.A(n_13937),
.B(n_2050),
.Y(n_14498)
);

INVx1_ASAP7_75t_L g14499 ( 
.A(n_14204),
.Y(n_14499)
);

OR2x2_ASAP7_75t_L g14500 ( 
.A(n_14206),
.B(n_13975),
.Y(n_14500)
);

INVx2_ASAP7_75t_L g14501 ( 
.A(n_14408),
.Y(n_14501)
);

A2O1A1Ixp33_ASAP7_75t_L g14502 ( 
.A1(n_14091),
.A2(n_13944),
.B(n_13952),
.C(n_13941),
.Y(n_14502)
);

OA21x2_ASAP7_75t_L g14503 ( 
.A1(n_14393),
.A2(n_13894),
.B(n_14049),
.Y(n_14503)
);

NAND2x1p5_ASAP7_75t_L g14504 ( 
.A(n_14451),
.B(n_13854),
.Y(n_14504)
);

HB1xp67_ASAP7_75t_L g14505 ( 
.A(n_14315),
.Y(n_14505)
);

INVx2_ASAP7_75t_SL g14506 ( 
.A(n_14497),
.Y(n_14506)
);

AND2x4_ASAP7_75t_L g14507 ( 
.A(n_14145),
.B(n_13687),
.Y(n_14507)
);

INVx1_ASAP7_75t_SL g14508 ( 
.A(n_14437),
.Y(n_14508)
);

AOI21xp5_ASAP7_75t_L g14509 ( 
.A1(n_14108),
.A2(n_13902),
.B(n_13766),
.Y(n_14509)
);

NAND3xp33_ASAP7_75t_L g14510 ( 
.A(n_14444),
.B(n_13860),
.C(n_13921),
.Y(n_14510)
);

AND2x4_ASAP7_75t_L g14511 ( 
.A(n_14256),
.B(n_13721),
.Y(n_14511)
);

NAND2xp5_ASAP7_75t_L g14512 ( 
.A(n_14086),
.B(n_14016),
.Y(n_14512)
);

AOI21xp5_ASAP7_75t_L g14513 ( 
.A1(n_14129),
.A2(n_13777),
.B(n_13775),
.Y(n_14513)
);

INVx1_ASAP7_75t_L g14514 ( 
.A(n_14231),
.Y(n_14514)
);

NAND2xp5_ASAP7_75t_L g14515 ( 
.A(n_14057),
.B(n_14035),
.Y(n_14515)
);

AO21x2_ASAP7_75t_L g14516 ( 
.A1(n_14155),
.A2(n_13632),
.B(n_13615),
.Y(n_14516)
);

INVx2_ASAP7_75t_L g14517 ( 
.A(n_14329),
.Y(n_14517)
);

NAND2x1p5_ASAP7_75t_L g14518 ( 
.A(n_14181),
.B(n_13854),
.Y(n_14518)
);

OAI21x1_ASAP7_75t_L g14519 ( 
.A1(n_14087),
.A2(n_13889),
.B(n_13874),
.Y(n_14519)
);

INVx1_ASAP7_75t_L g14520 ( 
.A(n_14242),
.Y(n_14520)
);

OA21x2_ASAP7_75t_L g14521 ( 
.A1(n_14395),
.A2(n_13910),
.B(n_13900),
.Y(n_14521)
);

NAND2xp5_ASAP7_75t_L g14522 ( 
.A(n_14147),
.B(n_13984),
.Y(n_14522)
);

BUFx2_ASAP7_75t_L g14523 ( 
.A(n_14154),
.Y(n_14523)
);

INVx1_ASAP7_75t_L g14524 ( 
.A(n_14246),
.Y(n_14524)
);

INVx1_ASAP7_75t_L g14525 ( 
.A(n_14266),
.Y(n_14525)
);

OAI21x1_ASAP7_75t_L g14526 ( 
.A1(n_14334),
.A2(n_13919),
.B(n_13917),
.Y(n_14526)
);

AOI21x1_ASAP7_75t_L g14527 ( 
.A1(n_14294),
.A2(n_13903),
.B(n_13957),
.Y(n_14527)
);

AO21x2_ASAP7_75t_L g14528 ( 
.A1(n_14220),
.A2(n_13646),
.B(n_13640),
.Y(n_14528)
);

INVx2_ASAP7_75t_L g14529 ( 
.A(n_14399),
.Y(n_14529)
);

OR2x2_ASAP7_75t_L g14530 ( 
.A(n_14364),
.B(n_13656),
.Y(n_14530)
);

OAI21x1_ASAP7_75t_L g14531 ( 
.A1(n_14350),
.A2(n_13950),
.B(n_13927),
.Y(n_14531)
);

NAND2xp5_ASAP7_75t_SL g14532 ( 
.A(n_14436),
.B(n_13878),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_14065),
.Y(n_14533)
);

INVx1_ASAP7_75t_L g14534 ( 
.A(n_14066),
.Y(n_14534)
);

AND2x4_ASAP7_75t_L g14535 ( 
.A(n_14286),
.B(n_13882),
.Y(n_14535)
);

AND2x2_ASAP7_75t_L g14536 ( 
.A(n_14197),
.B(n_13814),
.Y(n_14536)
);

AOI21xp5_ASAP7_75t_L g14537 ( 
.A1(n_14101),
.A2(n_14058),
.B(n_14158),
.Y(n_14537)
);

INVx1_ASAP7_75t_L g14538 ( 
.A(n_14075),
.Y(n_14538)
);

HB1xp67_ASAP7_75t_L g14539 ( 
.A(n_14421),
.Y(n_14539)
);

AOI21xp5_ASAP7_75t_L g14540 ( 
.A1(n_14172),
.A2(n_13570),
.B(n_13670),
.Y(n_14540)
);

NAND2xp5_ASAP7_75t_L g14541 ( 
.A(n_14234),
.B(n_13888),
.Y(n_14541)
);

INVx5_ASAP7_75t_SL g14542 ( 
.A(n_14470),
.Y(n_14542)
);

HB1xp67_ASAP7_75t_L g14543 ( 
.A(n_14463),
.Y(n_14543)
);

INVx1_ASAP7_75t_L g14544 ( 
.A(n_14097),
.Y(n_14544)
);

INVx2_ASAP7_75t_L g14545 ( 
.A(n_14400),
.Y(n_14545)
);

AO21x2_ASAP7_75t_L g14546 ( 
.A1(n_14456),
.A2(n_13697),
.B(n_13681),
.Y(n_14546)
);

INVxp67_ASAP7_75t_L g14547 ( 
.A(n_14070),
.Y(n_14547)
);

AO21x2_ASAP7_75t_L g14548 ( 
.A1(n_14466),
.A2(n_13717),
.B(n_13698),
.Y(n_14548)
);

OAI21x1_ASAP7_75t_L g14549 ( 
.A1(n_14323),
.A2(n_13983),
.B(n_13963),
.Y(n_14549)
);

CKINVDCx20_ASAP7_75t_R g14550 ( 
.A(n_14148),
.Y(n_14550)
);

NOR2xp33_ASAP7_75t_L g14551 ( 
.A(n_14185),
.B(n_13966),
.Y(n_14551)
);

INVx1_ASAP7_75t_L g14552 ( 
.A(n_14104),
.Y(n_14552)
);

AND2x2_ASAP7_75t_L g14553 ( 
.A(n_14134),
.B(n_13814),
.Y(n_14553)
);

INVx4_ASAP7_75t_L g14554 ( 
.A(n_14105),
.Y(n_14554)
);

OAI21x1_ASAP7_75t_L g14555 ( 
.A1(n_14337),
.A2(n_13986),
.B(n_14023),
.Y(n_14555)
);

AND2x2_ASAP7_75t_L g14556 ( 
.A(n_14119),
.B(n_13931),
.Y(n_14556)
);

A2O1A1Ixp33_ASAP7_75t_L g14557 ( 
.A1(n_14052),
.A2(n_14012),
.B(n_14009),
.C(n_13948),
.Y(n_14557)
);

OAI21x1_ASAP7_75t_SL g14558 ( 
.A1(n_14355),
.A2(n_13782),
.B(n_13802),
.Y(n_14558)
);

OAI21x1_ASAP7_75t_L g14559 ( 
.A1(n_14255),
.A2(n_13627),
.B(n_13652),
.Y(n_14559)
);

AOI21xp5_ASAP7_75t_L g14560 ( 
.A1(n_14209),
.A2(n_14195),
.B(n_14083),
.Y(n_14560)
);

INVx3_ASAP7_75t_L g14561 ( 
.A(n_14055),
.Y(n_14561)
);

HB1xp67_ASAP7_75t_L g14562 ( 
.A(n_14465),
.Y(n_14562)
);

NAND2xp5_ASAP7_75t_L g14563 ( 
.A(n_14151),
.B(n_14402),
.Y(n_14563)
);

INVx3_ASAP7_75t_L g14564 ( 
.A(n_14055),
.Y(n_14564)
);

AND2x6_ASAP7_75t_L g14565 ( 
.A(n_14429),
.B(n_13662),
.Y(n_14565)
);

OAI21xp5_ASAP7_75t_L g14566 ( 
.A1(n_14338),
.A2(n_14169),
.B(n_14233),
.Y(n_14566)
);

INVx2_ASAP7_75t_L g14567 ( 
.A(n_14053),
.Y(n_14567)
);

INVx1_ASAP7_75t_L g14568 ( 
.A(n_14109),
.Y(n_14568)
);

INVx1_ASAP7_75t_L g14569 ( 
.A(n_14120),
.Y(n_14569)
);

AND2x2_ASAP7_75t_L g14570 ( 
.A(n_14243),
.B(n_13873),
.Y(n_14570)
);

NOR2xp33_ASAP7_75t_L g14571 ( 
.A(n_14093),
.B(n_13875),
.Y(n_14571)
);

NAND2xp5_ASAP7_75t_L g14572 ( 
.A(n_14404),
.B(n_13734),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_14144),
.Y(n_14573)
);

INVxp67_ASAP7_75t_L g14574 ( 
.A(n_14229),
.Y(n_14574)
);

AOI21xp5_ASAP7_75t_L g14575 ( 
.A1(n_14127),
.A2(n_13736),
.B(n_13923),
.Y(n_14575)
);

AOI21xp5_ASAP7_75t_L g14576 ( 
.A1(n_14186),
.A2(n_13933),
.B(n_13835),
.Y(n_14576)
);

INVx1_ASAP7_75t_L g14577 ( 
.A(n_14165),
.Y(n_14577)
);

INVx1_ASAP7_75t_L g14578 ( 
.A(n_14179),
.Y(n_14578)
);

OAI21x1_ASAP7_75t_L g14579 ( 
.A1(n_14239),
.A2(n_13699),
.B(n_13820),
.Y(n_14579)
);

AOI21xp5_ASAP7_75t_L g14580 ( 
.A1(n_14252),
.A2(n_14218),
.B(n_14072),
.Y(n_14580)
);

OR2x6_ASAP7_75t_L g14581 ( 
.A(n_14236),
.B(n_13878),
.Y(n_14581)
);

CKINVDCx6p67_ASAP7_75t_R g14582 ( 
.A(n_14470),
.Y(n_14582)
);

AO31x2_ASAP7_75t_L g14583 ( 
.A1(n_14392),
.A2(n_14029),
.A3(n_14017),
.B(n_13954),
.Y(n_14583)
);

OR2x2_ASAP7_75t_L g14584 ( 
.A(n_14226),
.B(n_14103),
.Y(n_14584)
);

NAND2xp5_ASAP7_75t_L g14585 ( 
.A(n_14241),
.B(n_13705),
.Y(n_14585)
);

AND2x4_ASAP7_75t_L g14586 ( 
.A(n_14378),
.B(n_13668),
.Y(n_14586)
);

AOI21xp5_ASAP7_75t_L g14587 ( 
.A1(n_14141),
.A2(n_13861),
.B(n_13796),
.Y(n_14587)
);

OR2x6_ASAP7_75t_L g14588 ( 
.A(n_14095),
.B(n_13719),
.Y(n_14588)
);

OAI21x1_ASAP7_75t_L g14589 ( 
.A1(n_14223),
.A2(n_13561),
.B(n_13962),
.Y(n_14589)
);

INVx1_ASAP7_75t_SL g14590 ( 
.A(n_14343),
.Y(n_14590)
);

NAND2x1p5_ASAP7_75t_L g14591 ( 
.A(n_14222),
.B(n_13613),
.Y(n_14591)
);

AOI222xp33_ASAP7_75t_L g14592 ( 
.A1(n_14208),
.A2(n_13926),
.B1(n_13892),
.B2(n_13985),
.C1(n_13940),
.C2(n_13812),
.Y(n_14592)
);

NAND2xp5_ASAP7_75t_L g14593 ( 
.A(n_14132),
.B(n_14017),
.Y(n_14593)
);

AOI21xp5_ASAP7_75t_L g14594 ( 
.A1(n_14153),
.A2(n_14068),
.B(n_14328),
.Y(n_14594)
);

AOI21xp5_ASAP7_75t_L g14595 ( 
.A1(n_14116),
.A2(n_13976),
.B(n_13778),
.Y(n_14595)
);

BUFx3_ASAP7_75t_L g14596 ( 
.A(n_14238),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_14182),
.Y(n_14597)
);

OA21x2_ASAP7_75t_L g14598 ( 
.A1(n_14090),
.A2(n_13789),
.B(n_13746),
.Y(n_14598)
);

OAI21x1_ASAP7_75t_L g14599 ( 
.A1(n_14224),
.A2(n_13801),
.B(n_13819),
.Y(n_14599)
);

AO21x2_ASAP7_75t_L g14600 ( 
.A1(n_14439),
.A2(n_13821),
.B(n_13872),
.Y(n_14600)
);

INVx2_ASAP7_75t_L g14601 ( 
.A(n_14077),
.Y(n_14601)
);

INVx2_ASAP7_75t_SL g14602 ( 
.A(n_14094),
.Y(n_14602)
);

NAND2x1p5_ASAP7_75t_L g14603 ( 
.A(n_14436),
.B(n_13785),
.Y(n_14603)
);

INVx2_ASAP7_75t_L g14604 ( 
.A(n_14096),
.Y(n_14604)
);

INVx1_ASAP7_75t_L g14605 ( 
.A(n_14184),
.Y(n_14605)
);

OAI21x1_ASAP7_75t_L g14606 ( 
.A1(n_14176),
.A2(n_13829),
.B(n_14029),
.Y(n_14606)
);

OAI21x1_ASAP7_75t_L g14607 ( 
.A1(n_14171),
.A2(n_14029),
.B(n_13497),
.Y(n_14607)
);

NAND2xp5_ASAP7_75t_L g14608 ( 
.A(n_14138),
.B(n_13785),
.Y(n_14608)
);

INVx1_ASAP7_75t_SL g14609 ( 
.A(n_14341),
.Y(n_14609)
);

INVx2_ASAP7_75t_L g14610 ( 
.A(n_14342),
.Y(n_14610)
);

INVx5_ASAP7_75t_L g14611 ( 
.A(n_14455),
.Y(n_14611)
);

NAND2xp5_ASAP7_75t_L g14612 ( 
.A(n_14140),
.B(n_13482),
.Y(n_14612)
);

AOI21xp5_ASAP7_75t_L g14613 ( 
.A1(n_14202),
.A2(n_13619),
.B(n_13587),
.Y(n_14613)
);

INVx2_ASAP7_75t_L g14614 ( 
.A(n_14348),
.Y(n_14614)
);

OAI21x1_ASAP7_75t_L g14615 ( 
.A1(n_14173),
.A2(n_14200),
.B(n_14194),
.Y(n_14615)
);

INVx3_ASAP7_75t_L g14616 ( 
.A(n_14078),
.Y(n_14616)
);

AND2x4_ASAP7_75t_L g14617 ( 
.A(n_14418),
.B(n_13497),
.Y(n_14617)
);

OAI21x1_ASAP7_75t_L g14618 ( 
.A1(n_14143),
.A2(n_13564),
.B(n_13513),
.Y(n_14618)
);

INVx1_ASAP7_75t_L g14619 ( 
.A(n_14187),
.Y(n_14619)
);

NAND2xp5_ASAP7_75t_L g14620 ( 
.A(n_14146),
.B(n_13513),
.Y(n_14620)
);

OAI22xp33_ASAP7_75t_SL g14621 ( 
.A1(n_14139),
.A2(n_13564),
.B1(n_13634),
.B2(n_13619),
.Y(n_14621)
);

OA21x2_ASAP7_75t_L g14622 ( 
.A1(n_14264),
.A2(n_14221),
.B(n_14111),
.Y(n_14622)
);

AOI21xp5_ASAP7_75t_L g14623 ( 
.A1(n_14297),
.A2(n_13634),
.B(n_2050),
.Y(n_14623)
);

AND2x4_ASAP7_75t_L g14624 ( 
.A(n_14284),
.B(n_14124),
.Y(n_14624)
);

OA21x2_ASAP7_75t_L g14625 ( 
.A1(n_14063),
.A2(n_2051),
.B(n_2052),
.Y(n_14625)
);

OAI21x1_ASAP7_75t_L g14626 ( 
.A1(n_14125),
.A2(n_2051),
.B(n_2052),
.Y(n_14626)
);

OAI21x1_ASAP7_75t_L g14627 ( 
.A1(n_14088),
.A2(n_2053),
.B(n_2054),
.Y(n_14627)
);

AND2x4_ASAP7_75t_L g14628 ( 
.A(n_14361),
.B(n_2053),
.Y(n_14628)
);

AO21x2_ASAP7_75t_L g14629 ( 
.A1(n_14300),
.A2(n_2054),
.B(n_2055),
.Y(n_14629)
);

INVx1_ASAP7_75t_L g14630 ( 
.A(n_14199),
.Y(n_14630)
);

AO21x2_ASAP7_75t_L g14631 ( 
.A1(n_14253),
.A2(n_2055),
.B(n_2056),
.Y(n_14631)
);

AO21x2_ASAP7_75t_L g14632 ( 
.A1(n_14332),
.A2(n_2056),
.B(n_2057),
.Y(n_14632)
);

AO31x2_ASAP7_75t_L g14633 ( 
.A1(n_14180),
.A2(n_2059),
.A3(n_2057),
.B(n_2058),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_14227),
.Y(n_14634)
);

AOI21xp5_ASAP7_75t_L g14635 ( 
.A1(n_14113),
.A2(n_14084),
.B(n_14196),
.Y(n_14635)
);

INVx2_ASAP7_75t_L g14636 ( 
.A(n_14277),
.Y(n_14636)
);

INVx1_ASAP7_75t_L g14637 ( 
.A(n_14267),
.Y(n_14637)
);

CKINVDCx5p33_ASAP7_75t_R g14638 ( 
.A(n_14216),
.Y(n_14638)
);

AND2x2_ASAP7_75t_L g14639 ( 
.A(n_14401),
.B(n_2058),
.Y(n_14639)
);

BUFx3_ASAP7_75t_L g14640 ( 
.A(n_14100),
.Y(n_14640)
);

OAI21x1_ASAP7_75t_L g14641 ( 
.A1(n_14069),
.A2(n_2059),
.B(n_2060),
.Y(n_14641)
);

OR2x2_ASAP7_75t_L g14642 ( 
.A(n_14076),
.B(n_2060),
.Y(n_14642)
);

NOR2xp33_ASAP7_75t_SL g14643 ( 
.A(n_14318),
.B(n_2061),
.Y(n_14643)
);

NAND2xp5_ASAP7_75t_L g14644 ( 
.A(n_14415),
.B(n_2061),
.Y(n_14644)
);

BUFx10_ASAP7_75t_L g14645 ( 
.A(n_14248),
.Y(n_14645)
);

OAI21x1_ASAP7_75t_L g14646 ( 
.A1(n_14235),
.A2(n_2063),
.B(n_2064),
.Y(n_14646)
);

BUFx2_ASAP7_75t_L g14647 ( 
.A(n_14135),
.Y(n_14647)
);

NAND2xp5_ASAP7_75t_SL g14648 ( 
.A(n_14366),
.B(n_2065),
.Y(n_14648)
);

INVx1_ASAP7_75t_L g14649 ( 
.A(n_14270),
.Y(n_14649)
);

OAI21xp5_ASAP7_75t_L g14650 ( 
.A1(n_14215),
.A2(n_2065),
.B(n_2066),
.Y(n_14650)
);

OAI21x1_ASAP7_75t_L g14651 ( 
.A1(n_14079),
.A2(n_2066),
.B(n_2067),
.Y(n_14651)
);

INVx2_ASAP7_75t_L g14652 ( 
.A(n_14282),
.Y(n_14652)
);

INVx1_ASAP7_75t_L g14653 ( 
.A(n_14365),
.Y(n_14653)
);

AO31x2_ASAP7_75t_L g14654 ( 
.A1(n_14468),
.A2(n_2069),
.A3(n_2067),
.B(n_2068),
.Y(n_14654)
);

INVxp67_ASAP7_75t_SL g14655 ( 
.A(n_14207),
.Y(n_14655)
);

OAI21xp5_ASAP7_75t_L g14656 ( 
.A1(n_14219),
.A2(n_2068),
.B(n_2069),
.Y(n_14656)
);

INVx2_ASAP7_75t_L g14657 ( 
.A(n_14289),
.Y(n_14657)
);

NAND2xp5_ASAP7_75t_L g14658 ( 
.A(n_14110),
.B(n_2070),
.Y(n_14658)
);

OAI21x1_ASAP7_75t_L g14659 ( 
.A1(n_14130),
.A2(n_2070),
.B(n_2071),
.Y(n_14659)
);

INVx3_ASAP7_75t_L g14660 ( 
.A(n_14078),
.Y(n_14660)
);

BUFx3_ASAP7_75t_L g14661 ( 
.A(n_14092),
.Y(n_14661)
);

NAND2xp5_ASAP7_75t_L g14662 ( 
.A(n_14123),
.B(n_14259),
.Y(n_14662)
);

AO21x2_ASAP7_75t_L g14663 ( 
.A1(n_14333),
.A2(n_2071),
.B(n_2072),
.Y(n_14663)
);

OAI21xp5_ASAP7_75t_L g14664 ( 
.A1(n_14067),
.A2(n_2072),
.B(n_2073),
.Y(n_14664)
);

O2A1O1Ixp33_ASAP7_75t_L g14665 ( 
.A1(n_14189),
.A2(n_2075),
.B(n_2073),
.C(n_2074),
.Y(n_14665)
);

OAI221xp5_ASAP7_75t_L g14666 ( 
.A1(n_14054),
.A2(n_2076),
.B1(n_2074),
.B2(n_2075),
.C(n_2077),
.Y(n_14666)
);

AOI21xp5_ASAP7_75t_L g14667 ( 
.A1(n_14214),
.A2(n_2076),
.B(n_2077),
.Y(n_14667)
);

A2O1A1Ixp33_ASAP7_75t_L g14668 ( 
.A1(n_14281),
.A2(n_2080),
.B(n_2078),
.C(n_2079),
.Y(n_14668)
);

INVx2_ASAP7_75t_SL g14669 ( 
.A(n_14159),
.Y(n_14669)
);

INVx2_ASAP7_75t_L g14670 ( 
.A(n_14301),
.Y(n_14670)
);

INVx1_ASAP7_75t_L g14671 ( 
.A(n_14368),
.Y(n_14671)
);

INVx1_ASAP7_75t_L g14672 ( 
.A(n_14279),
.Y(n_14672)
);

INVx3_ASAP7_75t_L g14673 ( 
.A(n_14308),
.Y(n_14673)
);

OA21x2_ASAP7_75t_L g14674 ( 
.A1(n_14295),
.A2(n_2078),
.B(n_2080),
.Y(n_14674)
);

INVx1_ASAP7_75t_L g14675 ( 
.A(n_14383),
.Y(n_14675)
);

BUFx3_ASAP7_75t_L g14676 ( 
.A(n_14302),
.Y(n_14676)
);

AND2x2_ASAP7_75t_L g14677 ( 
.A(n_14403),
.B(n_2081),
.Y(n_14677)
);

AND3x1_ASAP7_75t_L g14678 ( 
.A(n_14064),
.B(n_2082),
.C(n_2083),
.Y(n_14678)
);

BUFx8_ASAP7_75t_L g14679 ( 
.A(n_14308),
.Y(n_14679)
);

OR2x2_ASAP7_75t_L g14680 ( 
.A(n_14073),
.B(n_2082),
.Y(n_14680)
);

INVx3_ASAP7_75t_L g14681 ( 
.A(n_14377),
.Y(n_14681)
);

OAI21x1_ASAP7_75t_L g14682 ( 
.A1(n_14061),
.A2(n_2083),
.B(n_2084),
.Y(n_14682)
);

HB1xp67_ASAP7_75t_L g14683 ( 
.A(n_14152),
.Y(n_14683)
);

HB1xp67_ASAP7_75t_L g14684 ( 
.A(n_14217),
.Y(n_14684)
);

INVx1_ASAP7_75t_L g14685 ( 
.A(n_14114),
.Y(n_14685)
);

NOR2xp33_ASAP7_75t_L g14686 ( 
.A(n_14483),
.B(n_2085),
.Y(n_14686)
);

NOR4xp25_ASAP7_75t_L g14687 ( 
.A(n_14412),
.B(n_2087),
.C(n_2085),
.D(n_2086),
.Y(n_14687)
);

A2O1A1Ixp33_ASAP7_75t_L g14688 ( 
.A1(n_14150),
.A2(n_2088),
.B(n_2086),
.C(n_2087),
.Y(n_14688)
);

OAI21x1_ASAP7_75t_L g14689 ( 
.A1(n_14168),
.A2(n_2089),
.B(n_2090),
.Y(n_14689)
);

OR2x6_ASAP7_75t_L g14690 ( 
.A(n_14142),
.B(n_2089),
.Y(n_14690)
);

AO21x2_ASAP7_75t_L g14691 ( 
.A1(n_14344),
.A2(n_2091),
.B(n_2092),
.Y(n_14691)
);

INVx1_ASAP7_75t_L g14692 ( 
.A(n_14121),
.Y(n_14692)
);

OAI21x1_ASAP7_75t_L g14693 ( 
.A1(n_14074),
.A2(n_14354),
.B(n_14339),
.Y(n_14693)
);

OAI21x1_ASAP7_75t_L g14694 ( 
.A1(n_14356),
.A2(n_2093),
.B(n_2094),
.Y(n_14694)
);

INVx3_ASAP7_75t_L g14695 ( 
.A(n_14384),
.Y(n_14695)
);

AOI21xp5_ASAP7_75t_L g14696 ( 
.A1(n_14419),
.A2(n_2095),
.B(n_2096),
.Y(n_14696)
);

AOI21xp33_ASAP7_75t_L g14697 ( 
.A1(n_14112),
.A2(n_2096),
.B(n_2097),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_14149),
.Y(n_14698)
);

AOI22xp5_ASAP7_75t_L g14699 ( 
.A1(n_14056),
.A2(n_2100),
.B1(n_2097),
.B2(n_2099),
.Y(n_14699)
);

NAND2x1p5_ASAP7_75t_L g14700 ( 
.A(n_14375),
.B(n_2099),
.Y(n_14700)
);

AND2x2_ASAP7_75t_L g14701 ( 
.A(n_14474),
.B(n_2100),
.Y(n_14701)
);

AOI21xp33_ASAP7_75t_SL g14702 ( 
.A1(n_14296),
.A2(n_14189),
.B(n_14213),
.Y(n_14702)
);

OAI21x1_ASAP7_75t_L g14703 ( 
.A1(n_14071),
.A2(n_14203),
.B(n_14170),
.Y(n_14703)
);

BUFx8_ASAP7_75t_SL g14704 ( 
.A(n_14162),
.Y(n_14704)
);

NAND2xp5_ASAP7_75t_L g14705 ( 
.A(n_14081),
.B(n_14085),
.Y(n_14705)
);

OA21x2_ASAP7_75t_L g14706 ( 
.A1(n_14335),
.A2(n_2101),
.B(n_2102),
.Y(n_14706)
);

A2O1A1Ixp33_ASAP7_75t_L g14707 ( 
.A1(n_14098),
.A2(n_2104),
.B(n_2101),
.C(n_2103),
.Y(n_14707)
);

INVx1_ASAP7_75t_L g14708 ( 
.A(n_14389),
.Y(n_14708)
);

CKINVDCx16_ASAP7_75t_R g14709 ( 
.A(n_14358),
.Y(n_14709)
);

OR2x2_ASAP7_75t_L g14710 ( 
.A(n_14089),
.B(n_2103),
.Y(n_14710)
);

AO21x2_ASAP7_75t_L g14711 ( 
.A1(n_14349),
.A2(n_2104),
.B(n_2105),
.Y(n_14711)
);

INVx1_ASAP7_75t_L g14712 ( 
.A(n_14352),
.Y(n_14712)
);

OR2x2_ASAP7_75t_L g14713 ( 
.A(n_14458),
.B(n_2105),
.Y(n_14713)
);

BUFx6f_ASAP7_75t_L g14714 ( 
.A(n_14162),
.Y(n_14714)
);

INVx1_ASAP7_75t_L g14715 ( 
.A(n_14353),
.Y(n_14715)
);

OAI21x1_ASAP7_75t_SL g14716 ( 
.A1(n_14291),
.A2(n_2106),
.B(n_2107),
.Y(n_14716)
);

NOR2xp33_ASAP7_75t_L g14717 ( 
.A(n_14157),
.B(n_2107),
.Y(n_14717)
);

NAND2x1p5_ASAP7_75t_L g14718 ( 
.A(n_14257),
.B(n_2108),
.Y(n_14718)
);

INVx4_ASAP7_75t_L g14719 ( 
.A(n_14159),
.Y(n_14719)
);

OAI21xp5_ASAP7_75t_L g14720 ( 
.A1(n_14225),
.A2(n_14405),
.B(n_14201),
.Y(n_14720)
);

A2O1A1Ixp33_ASAP7_75t_L g14721 ( 
.A1(n_14464),
.A2(n_2110),
.B(n_2108),
.C(n_2109),
.Y(n_14721)
);

AND2x4_ASAP7_75t_L g14722 ( 
.A(n_14244),
.B(n_2109),
.Y(n_14722)
);

NAND2xp5_ASAP7_75t_L g14723 ( 
.A(n_14240),
.B(n_2110),
.Y(n_14723)
);

INVx1_ASAP7_75t_SL g14724 ( 
.A(n_14398),
.Y(n_14724)
);

OAI21x1_ASAP7_75t_L g14725 ( 
.A1(n_14306),
.A2(n_2111),
.B(n_2112),
.Y(n_14725)
);

AND2x2_ASAP7_75t_L g14726 ( 
.A(n_14106),
.B(n_2111),
.Y(n_14726)
);

OAI21x1_ASAP7_75t_L g14727 ( 
.A1(n_14313),
.A2(n_2112),
.B(n_2113),
.Y(n_14727)
);

BUFx3_ASAP7_75t_L g14728 ( 
.A(n_14237),
.Y(n_14728)
);

AO21x2_ASAP7_75t_L g14729 ( 
.A1(n_14390),
.A2(n_2113),
.B(n_2114),
.Y(n_14729)
);

CKINVDCx14_ASAP7_75t_R g14730 ( 
.A(n_14479),
.Y(n_14730)
);

NAND2xp5_ASAP7_75t_L g14731 ( 
.A(n_14228),
.B(n_2114),
.Y(n_14731)
);

INVx2_ASAP7_75t_L g14732 ( 
.A(n_14330),
.Y(n_14732)
);

NAND2xp5_ASAP7_75t_L g14733 ( 
.A(n_14099),
.B(n_2115),
.Y(n_14733)
);

INVx1_ASAP7_75t_L g14734 ( 
.A(n_14232),
.Y(n_14734)
);

AND2x4_ASAP7_75t_L g14735 ( 
.A(n_14487),
.B(n_14126),
.Y(n_14735)
);

INVx2_ASAP7_75t_SL g14736 ( 
.A(n_14472),
.Y(n_14736)
);

BUFx2_ASAP7_75t_L g14737 ( 
.A(n_14059),
.Y(n_14737)
);

OA21x2_ASAP7_75t_L g14738 ( 
.A1(n_14247),
.A2(n_2115),
.B(n_2116),
.Y(n_14738)
);

INVx1_ASAP7_75t_L g14739 ( 
.A(n_14137),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_14376),
.Y(n_14740)
);

INVx2_ASAP7_75t_SL g14741 ( 
.A(n_14472),
.Y(n_14741)
);

INVx1_ASAP7_75t_L g14742 ( 
.A(n_14336),
.Y(n_14742)
);

AO31x2_ASAP7_75t_L g14743 ( 
.A1(n_14443),
.A2(n_2118),
.A3(n_2116),
.B(n_2117),
.Y(n_14743)
);

AOI21xp5_ASAP7_75t_L g14744 ( 
.A1(n_14369),
.A2(n_2117),
.B(n_2118),
.Y(n_14744)
);

AND2x2_ASAP7_75t_L g14745 ( 
.A(n_14469),
.B(n_2119),
.Y(n_14745)
);

CKINVDCx11_ASAP7_75t_R g14746 ( 
.A(n_14414),
.Y(n_14746)
);

INVx1_ASAP7_75t_L g14747 ( 
.A(n_14450),
.Y(n_14747)
);

AND2x2_ASAP7_75t_L g14748 ( 
.A(n_14385),
.B(n_2119),
.Y(n_14748)
);

OA21x2_ASAP7_75t_L g14749 ( 
.A1(n_14107),
.A2(n_2120),
.B(n_2121),
.Y(n_14749)
);

AO31x2_ASAP7_75t_L g14750 ( 
.A1(n_14319),
.A2(n_2122),
.A3(n_2120),
.B(n_2121),
.Y(n_14750)
);

INVx1_ASAP7_75t_L g14751 ( 
.A(n_14471),
.Y(n_14751)
);

NAND2x1p5_ASAP7_75t_L g14752 ( 
.A(n_14265),
.B(n_2124),
.Y(n_14752)
);

INVx2_ASAP7_75t_L g14753 ( 
.A(n_14340),
.Y(n_14753)
);

AOI222xp33_ASAP7_75t_L g14754 ( 
.A1(n_14457),
.A2(n_2126),
.B1(n_2128),
.B2(n_2124),
.C1(n_2125),
.C2(n_2127),
.Y(n_14754)
);

OAI21xp33_ASAP7_75t_SL g14755 ( 
.A1(n_14164),
.A2(n_2125),
.B(n_2126),
.Y(n_14755)
);

INVx1_ASAP7_75t_L g14756 ( 
.A(n_14118),
.Y(n_14756)
);

NAND2xp5_ASAP7_75t_L g14757 ( 
.A(n_14304),
.B(n_2127),
.Y(n_14757)
);

NOR2x1_ASAP7_75t_SL g14758 ( 
.A(n_14142),
.B(n_2128),
.Y(n_14758)
);

AOI21xp5_ASAP7_75t_L g14759 ( 
.A1(n_14210),
.A2(n_2129),
.B(n_2130),
.Y(n_14759)
);

A2O1A1Ixp33_ASAP7_75t_L g14760 ( 
.A1(n_14128),
.A2(n_2131),
.B(n_2129),
.C(n_2130),
.Y(n_14760)
);

INVx3_ASAP7_75t_L g14761 ( 
.A(n_14391),
.Y(n_14761)
);

AND2x2_ASAP7_75t_L g14762 ( 
.A(n_14406),
.B(n_2131),
.Y(n_14762)
);

AND2x2_ASAP7_75t_L g14763 ( 
.A(n_14432),
.B(n_2132),
.Y(n_14763)
);

NAND2xp5_ASAP7_75t_L g14764 ( 
.A(n_14438),
.B(n_2132),
.Y(n_14764)
);

INVx3_ASAP7_75t_L g14765 ( 
.A(n_14249),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14360),
.Y(n_14766)
);

OAI21x1_ASAP7_75t_L g14767 ( 
.A1(n_14062),
.A2(n_2133),
.B(n_2134),
.Y(n_14767)
);

BUFx2_ASAP7_75t_L g14768 ( 
.A(n_14193),
.Y(n_14768)
);

INVx1_ASAP7_75t_L g14769 ( 
.A(n_14424),
.Y(n_14769)
);

BUFx2_ASAP7_75t_L g14770 ( 
.A(n_14287),
.Y(n_14770)
);

AND2x2_ASAP7_75t_L g14771 ( 
.A(n_14446),
.B(n_2134),
.Y(n_14771)
);

NAND2xp5_ASAP7_75t_L g14772 ( 
.A(n_14477),
.B(n_2135),
.Y(n_14772)
);

OAI22xp5_ASAP7_75t_L g14773 ( 
.A1(n_14133),
.A2(n_2137),
.B1(n_2135),
.B2(n_2136),
.Y(n_14773)
);

INVx1_ASAP7_75t_SL g14774 ( 
.A(n_14467),
.Y(n_14774)
);

AND2x4_ASAP7_75t_L g14775 ( 
.A(n_14188),
.B(n_2136),
.Y(n_14775)
);

INVx6_ASAP7_75t_L g14776 ( 
.A(n_14448),
.Y(n_14776)
);

INVx1_ASAP7_75t_L g14777 ( 
.A(n_14230),
.Y(n_14777)
);

NAND2xp5_ASAP7_75t_L g14778 ( 
.A(n_14484),
.B(n_2138),
.Y(n_14778)
);

NOR2xp33_ASAP7_75t_L g14779 ( 
.A(n_14115),
.B(n_2138),
.Y(n_14779)
);

HB1xp67_ASAP7_75t_L g14780 ( 
.A(n_14309),
.Y(n_14780)
);

AO22x1_ASAP7_75t_L g14781 ( 
.A1(n_14163),
.A2(n_2141),
.B1(n_2139),
.B2(n_2140),
.Y(n_14781)
);

NAND2xp5_ASAP7_75t_L g14782 ( 
.A(n_14488),
.B(n_2139),
.Y(n_14782)
);

INVx1_ASAP7_75t_L g14783 ( 
.A(n_14307),
.Y(n_14783)
);

OA21x2_ASAP7_75t_L g14784 ( 
.A1(n_14254),
.A2(n_2141),
.B(n_2142),
.Y(n_14784)
);

NAND2xp5_ASAP7_75t_L g14785 ( 
.A(n_14280),
.B(n_2142),
.Y(n_14785)
);

NAND2xp5_ASAP7_75t_L g14786 ( 
.A(n_14205),
.B(n_2143),
.Y(n_14786)
);

OR2x2_ASAP7_75t_L g14787 ( 
.A(n_14276),
.B(n_2144),
.Y(n_14787)
);

BUFx3_ASAP7_75t_L g14788 ( 
.A(n_14386),
.Y(n_14788)
);

NAND2xp5_ASAP7_75t_SL g14789 ( 
.A(n_14288),
.B(n_2144),
.Y(n_14789)
);

NAND2xp5_ASAP7_75t_L g14790 ( 
.A(n_14324),
.B(n_2145),
.Y(n_14790)
);

OA21x2_ASAP7_75t_L g14791 ( 
.A1(n_14191),
.A2(n_14192),
.B(n_14245),
.Y(n_14791)
);

OAI21x1_ASAP7_75t_L g14792 ( 
.A1(n_14178),
.A2(n_2145),
.B(n_2146),
.Y(n_14792)
);

AOI21x1_ASAP7_75t_L g14793 ( 
.A1(n_14371),
.A2(n_2146),
.B(n_2147),
.Y(n_14793)
);

AOI22xp5_ASAP7_75t_L g14794 ( 
.A1(n_14250),
.A2(n_2149),
.B1(n_2147),
.B2(n_2148),
.Y(n_14794)
);

OAI22xp5_ASAP7_75t_SL g14795 ( 
.A1(n_14269),
.A2(n_2150),
.B1(n_2148),
.B2(n_2149),
.Y(n_14795)
);

AND2x4_ASAP7_75t_L g14796 ( 
.A(n_14357),
.B(n_14372),
.Y(n_14796)
);

BUFx6f_ASAP7_75t_L g14797 ( 
.A(n_14448),
.Y(n_14797)
);

INVx1_ASAP7_75t_L g14798 ( 
.A(n_14261),
.Y(n_14798)
);

CKINVDCx11_ASAP7_75t_R g14799 ( 
.A(n_14396),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_14311),
.Y(n_14800)
);

NOR2x1_ASAP7_75t_SL g14801 ( 
.A(n_14370),
.B(n_2151),
.Y(n_14801)
);

AO31x2_ASAP7_75t_L g14802 ( 
.A1(n_14285),
.A2(n_2153),
.A3(n_2151),
.B(n_2152),
.Y(n_14802)
);

OAI21x1_ASAP7_75t_L g14803 ( 
.A1(n_14212),
.A2(n_2152),
.B(n_2153),
.Y(n_14803)
);

AOI21xp5_ASAP7_75t_L g14804 ( 
.A1(n_14102),
.A2(n_2154),
.B(n_2155),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_14311),
.Y(n_14805)
);

OAI22xp5_ASAP7_75t_L g14806 ( 
.A1(n_14382),
.A2(n_2156),
.B1(n_2154),
.B2(n_2155),
.Y(n_14806)
);

INVx1_ASAP7_75t_L g14807 ( 
.A(n_14251),
.Y(n_14807)
);

AOI21x1_ASAP7_75t_L g14808 ( 
.A1(n_14498),
.A2(n_2156),
.B(n_2157),
.Y(n_14808)
);

OR2x2_ASAP7_75t_L g14809 ( 
.A(n_14211),
.B(n_2157),
.Y(n_14809)
);

CKINVDCx20_ASAP7_75t_R g14810 ( 
.A(n_14271),
.Y(n_14810)
);

AOI21xp5_ASAP7_75t_L g14811 ( 
.A1(n_14314),
.A2(n_2158),
.B(n_2159),
.Y(n_14811)
);

AO21x2_ASAP7_75t_L g14812 ( 
.A1(n_14321),
.A2(n_2158),
.B(n_2159),
.Y(n_14812)
);

NOR2xp33_ASAP7_75t_L g14813 ( 
.A(n_14492),
.B(n_2160),
.Y(n_14813)
);

AND2x2_ASAP7_75t_L g14814 ( 
.A(n_14388),
.B(n_2161),
.Y(n_14814)
);

NAND2xp5_ASAP7_75t_L g14815 ( 
.A(n_14060),
.B(n_2162),
.Y(n_14815)
);

BUFx2_ASAP7_75t_SL g14816 ( 
.A(n_14428),
.Y(n_14816)
);

BUFx2_ASAP7_75t_L g14817 ( 
.A(n_14163),
.Y(n_14817)
);

NAND2xp5_ASAP7_75t_L g14818 ( 
.A(n_14312),
.B(n_2162),
.Y(n_14818)
);

NAND2xp5_ASAP7_75t_L g14819 ( 
.A(n_14299),
.B(n_2163),
.Y(n_14819)
);

AND2x2_ASAP7_75t_L g14820 ( 
.A(n_14327),
.B(n_14417),
.Y(n_14820)
);

AOI22xp5_ASAP7_75t_L g14821 ( 
.A1(n_14163),
.A2(n_2165),
.B1(n_2163),
.B2(n_2164),
.Y(n_14821)
);

AND2x4_ASAP7_75t_SL g14822 ( 
.A(n_14262),
.B(n_2164),
.Y(n_14822)
);

INVx1_ASAP7_75t_L g14823 ( 
.A(n_14407),
.Y(n_14823)
);

BUFx6f_ASAP7_75t_L g14824 ( 
.A(n_14489),
.Y(n_14824)
);

AND2x4_ASAP7_75t_L g14825 ( 
.A(n_14117),
.B(n_2165),
.Y(n_14825)
);

CKINVDCx5p33_ASAP7_75t_R g14826 ( 
.A(n_14293),
.Y(n_14826)
);

INVx2_ASAP7_75t_SL g14827 ( 
.A(n_14305),
.Y(n_14827)
);

OAI21x1_ASAP7_75t_L g14828 ( 
.A1(n_14160),
.A2(n_2166),
.B(n_2167),
.Y(n_14828)
);

OA21x2_ASAP7_75t_L g14829 ( 
.A1(n_14183),
.A2(n_2166),
.B(n_2168),
.Y(n_14829)
);

BUFx3_ASAP7_75t_L g14830 ( 
.A(n_14273),
.Y(n_14830)
);

AND2x2_ASAP7_75t_L g14831 ( 
.A(n_14434),
.B(n_2168),
.Y(n_14831)
);

A2O1A1Ixp33_ASAP7_75t_L g14832 ( 
.A1(n_14322),
.A2(n_2172),
.B(n_2169),
.C(n_2171),
.Y(n_14832)
);

INVx1_ASAP7_75t_L g14833 ( 
.A(n_14426),
.Y(n_14833)
);

INVx1_ASAP7_75t_L g14834 ( 
.A(n_14435),
.Y(n_14834)
);

NOR2xp33_ASAP7_75t_L g14835 ( 
.A(n_14493),
.B(n_2171),
.Y(n_14835)
);

NAND2xp5_ASAP7_75t_L g14836 ( 
.A(n_14490),
.B(n_2172),
.Y(n_14836)
);

AO31x2_ASAP7_75t_L g14837 ( 
.A1(n_14431),
.A2(n_2175),
.A3(n_2173),
.B(n_2174),
.Y(n_14837)
);

NAND2x1p5_ASAP7_75t_L g14838 ( 
.A(n_14381),
.B(n_2173),
.Y(n_14838)
);

AO21x2_ASAP7_75t_L g14839 ( 
.A1(n_14409),
.A2(n_2174),
.B(n_2175),
.Y(n_14839)
);

INVx1_ASAP7_75t_L g14840 ( 
.A(n_14272),
.Y(n_14840)
);

INVx1_ASAP7_75t_L g14841 ( 
.A(n_14274),
.Y(n_14841)
);

INVxp67_ASAP7_75t_L g14842 ( 
.A(n_14320),
.Y(n_14842)
);

INVx3_ASAP7_75t_L g14843 ( 
.A(n_14482),
.Y(n_14843)
);

INVx1_ASAP7_75t_L g14844 ( 
.A(n_14275),
.Y(n_14844)
);

NAND2x1p5_ASAP7_75t_L g14845 ( 
.A(n_14290),
.B(n_2176),
.Y(n_14845)
);

NAND2xp5_ASAP7_75t_L g14846 ( 
.A(n_14175),
.B(n_14445),
.Y(n_14846)
);

INVx1_ASAP7_75t_SL g14847 ( 
.A(n_14422),
.Y(n_14847)
);

INVx1_ASAP7_75t_L g14848 ( 
.A(n_14278),
.Y(n_14848)
);

BUFx3_ASAP7_75t_L g14849 ( 
.A(n_14460),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_14283),
.Y(n_14850)
);

INVx1_ASAP7_75t_L g14851 ( 
.A(n_14263),
.Y(n_14851)
);

NAND2xp5_ASAP7_75t_L g14852 ( 
.A(n_14198),
.B(n_2176),
.Y(n_14852)
);

AND2x2_ASAP7_75t_L g14853 ( 
.A(n_14190),
.B(n_2177),
.Y(n_14853)
);

INVx3_ASAP7_75t_L g14854 ( 
.A(n_14317),
.Y(n_14854)
);

INVx2_ASAP7_75t_L g14855 ( 
.A(n_14326),
.Y(n_14855)
);

OA21x2_ASAP7_75t_L g14856 ( 
.A1(n_14174),
.A2(n_14177),
.B(n_14122),
.Y(n_14856)
);

AOI21xp5_ASAP7_75t_L g14857 ( 
.A1(n_14325),
.A2(n_2177),
.B(n_2178),
.Y(n_14857)
);

AND2x2_ASAP7_75t_L g14858 ( 
.A(n_14136),
.B(n_2179),
.Y(n_14858)
);

AND2x4_ASAP7_75t_L g14859 ( 
.A(n_14131),
.B(n_2180),
.Y(n_14859)
);

AND2x4_ASAP7_75t_L g14860 ( 
.A(n_14161),
.B(n_2181),
.Y(n_14860)
);

INVx1_ASAP7_75t_L g14861 ( 
.A(n_14411),
.Y(n_14861)
);

AOI21xp5_ASAP7_75t_L g14862 ( 
.A1(n_14394),
.A2(n_2181),
.B(n_2182),
.Y(n_14862)
);

OAI21xp5_ASAP7_75t_L g14863 ( 
.A1(n_14359),
.A2(n_2182),
.B(n_2183),
.Y(n_14863)
);

INVx5_ASAP7_75t_L g14864 ( 
.A(n_14486),
.Y(n_14864)
);

AOI22xp33_ASAP7_75t_L g14865 ( 
.A1(n_14167),
.A2(n_2185),
.B1(n_2183),
.B2(n_2184),
.Y(n_14865)
);

NOR2xp33_ASAP7_75t_L g14866 ( 
.A(n_14496),
.B(n_2184),
.Y(n_14866)
);

AO21x2_ASAP7_75t_L g14867 ( 
.A1(n_14298),
.A2(n_2185),
.B(n_2186),
.Y(n_14867)
);

NAND2xp5_ASAP7_75t_L g14868 ( 
.A(n_14420),
.B(n_2186),
.Y(n_14868)
);

INVx1_ASAP7_75t_L g14869 ( 
.A(n_14442),
.Y(n_14869)
);

AOI22xp5_ASAP7_75t_L g14870 ( 
.A1(n_14346),
.A2(n_2189),
.B1(n_2187),
.B2(n_2188),
.Y(n_14870)
);

INVx1_ASAP7_75t_L g14871 ( 
.A(n_14363),
.Y(n_14871)
);

OAI21x1_ASAP7_75t_L g14872 ( 
.A1(n_14082),
.A2(n_2187),
.B(n_2188),
.Y(n_14872)
);

OAI21x1_ASAP7_75t_L g14873 ( 
.A1(n_14292),
.A2(n_2189),
.B(n_2190),
.Y(n_14873)
);

INVx1_ASAP7_75t_L g14874 ( 
.A(n_14473),
.Y(n_14874)
);

AO31x2_ASAP7_75t_L g14875 ( 
.A1(n_14475),
.A2(n_2193),
.A3(n_2191),
.B(n_2192),
.Y(n_14875)
);

AND2x4_ASAP7_75t_L g14876 ( 
.A(n_14397),
.B(n_2191),
.Y(n_14876)
);

AOI21xp33_ASAP7_75t_SL g14877 ( 
.A1(n_14373),
.A2(n_14441),
.B(n_14476),
.Y(n_14877)
);

INVx2_ASAP7_75t_SL g14878 ( 
.A(n_14331),
.Y(n_14878)
);

CKINVDCx20_ASAP7_75t_R g14879 ( 
.A(n_14481),
.Y(n_14879)
);

INVx1_ASAP7_75t_L g14880 ( 
.A(n_14425),
.Y(n_14880)
);

OAI21x1_ASAP7_75t_L g14881 ( 
.A1(n_14367),
.A2(n_2192),
.B(n_2193),
.Y(n_14881)
);

HB1xp67_ASAP7_75t_L g14882 ( 
.A(n_14379),
.Y(n_14882)
);

INVx1_ASAP7_75t_L g14883 ( 
.A(n_14380),
.Y(n_14883)
);

NAND2x1p5_ASAP7_75t_L g14884 ( 
.A(n_14410),
.B(n_2194),
.Y(n_14884)
);

INVx2_ASAP7_75t_SL g14885 ( 
.A(n_14413),
.Y(n_14885)
);

INVx2_ASAP7_75t_L g14886 ( 
.A(n_14166),
.Y(n_14886)
);

BUFx6f_ASAP7_75t_L g14887 ( 
.A(n_14387),
.Y(n_14887)
);

NAND2xp5_ASAP7_75t_SL g14888 ( 
.A(n_14453),
.B(n_14374),
.Y(n_14888)
);

INVx2_ASAP7_75t_L g14889 ( 
.A(n_14345),
.Y(n_14889)
);

NAND2xp5_ASAP7_75t_L g14890 ( 
.A(n_14080),
.B(n_2194),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_14347),
.Y(n_14891)
);

OAI21xp5_ASAP7_75t_L g14892 ( 
.A1(n_14362),
.A2(n_2195),
.B(n_2196),
.Y(n_14892)
);

OR2x2_ASAP7_75t_L g14893 ( 
.A(n_14539),
.B(n_14080),
.Y(n_14893)
);

NAND2xp5_ASAP7_75t_L g14894 ( 
.A(n_14864),
.B(n_14351),
.Y(n_14894)
);

OAI21x1_ASAP7_75t_L g14895 ( 
.A1(n_14703),
.A2(n_14416),
.B(n_14423),
.Y(n_14895)
);

AND2x2_ASAP7_75t_L g14896 ( 
.A(n_14609),
.B(n_14156),
.Y(n_14896)
);

INVx2_ASAP7_75t_L g14897 ( 
.A(n_14596),
.Y(n_14897)
);

INVx1_ASAP7_75t_L g14898 ( 
.A(n_14499),
.Y(n_14898)
);

OA21x2_ASAP7_75t_L g14899 ( 
.A1(n_14720),
.A2(n_14433),
.B(n_14427),
.Y(n_14899)
);

BUFx4f_ASAP7_75t_SL g14900 ( 
.A(n_14679),
.Y(n_14900)
);

NAND2xp5_ASAP7_75t_L g14901 ( 
.A(n_14864),
.B(n_14440),
.Y(n_14901)
);

INVx1_ASAP7_75t_L g14902 ( 
.A(n_14514),
.Y(n_14902)
);

INVx1_ASAP7_75t_L g14903 ( 
.A(n_14520),
.Y(n_14903)
);

CKINVDCx5p33_ASAP7_75t_R g14904 ( 
.A(n_14550),
.Y(n_14904)
);

INVx1_ASAP7_75t_L g14905 ( 
.A(n_14524),
.Y(n_14905)
);

INVx2_ASAP7_75t_L g14906 ( 
.A(n_14737),
.Y(n_14906)
);

CKINVDCx12_ASAP7_75t_R g14907 ( 
.A(n_14690),
.Y(n_14907)
);

INVx2_ASAP7_75t_L g14908 ( 
.A(n_14768),
.Y(n_14908)
);

NOR2xp33_ASAP7_75t_L g14909 ( 
.A(n_14554),
.B(n_14452),
.Y(n_14909)
);

HB1xp67_ASAP7_75t_L g14910 ( 
.A(n_14505),
.Y(n_14910)
);

INVx2_ASAP7_75t_SL g14911 ( 
.A(n_14611),
.Y(n_14911)
);

INVx2_ASAP7_75t_L g14912 ( 
.A(n_14570),
.Y(n_14912)
);

CKINVDCx5p33_ASAP7_75t_R g14913 ( 
.A(n_14638),
.Y(n_14913)
);

INVx2_ASAP7_75t_L g14914 ( 
.A(n_14536),
.Y(n_14914)
);

BUFx2_ASAP7_75t_L g14915 ( 
.A(n_14588),
.Y(n_14915)
);

AO21x1_ASAP7_75t_L g14916 ( 
.A1(n_14540),
.A2(n_14303),
.B(n_14485),
.Y(n_14916)
);

INVx2_ASAP7_75t_L g14917 ( 
.A(n_14504),
.Y(n_14917)
);

INVx3_ASAP7_75t_L g14918 ( 
.A(n_14704),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_14525),
.Y(n_14919)
);

INVx1_ASAP7_75t_L g14920 ( 
.A(n_14533),
.Y(n_14920)
);

INVx1_ASAP7_75t_L g14921 ( 
.A(n_14534),
.Y(n_14921)
);

INVxp67_ASAP7_75t_L g14922 ( 
.A(n_14817),
.Y(n_14922)
);

AND2x2_ASAP7_75t_L g14923 ( 
.A(n_14553),
.B(n_14156),
.Y(n_14923)
);

INVx1_ASAP7_75t_L g14924 ( 
.A(n_14538),
.Y(n_14924)
);

BUFx2_ASAP7_75t_SL g14925 ( 
.A(n_14611),
.Y(n_14925)
);

OR2x2_ASAP7_75t_L g14926 ( 
.A(n_14530),
.B(n_14512),
.Y(n_14926)
);

INVx2_ASAP7_75t_L g14927 ( 
.A(n_14600),
.Y(n_14927)
);

INVx1_ASAP7_75t_L g14928 ( 
.A(n_14544),
.Y(n_14928)
);

INVx1_ASAP7_75t_L g14929 ( 
.A(n_14552),
.Y(n_14929)
);

NAND2xp5_ASAP7_75t_L g14930 ( 
.A(n_14667),
.B(n_14447),
.Y(n_14930)
);

OR2x6_ASAP7_75t_L g14931 ( 
.A(n_14690),
.B(n_14449),
.Y(n_14931)
);

NAND2xp5_ASAP7_75t_L g14932 ( 
.A(n_14513),
.B(n_14454),
.Y(n_14932)
);

OAI21xp5_ASAP7_75t_L g14933 ( 
.A1(n_14560),
.A2(n_14310),
.B(n_14495),
.Y(n_14933)
);

INVx2_ASAP7_75t_L g14934 ( 
.A(n_14681),
.Y(n_14934)
);

INVx2_ASAP7_75t_L g14935 ( 
.A(n_14695),
.Y(n_14935)
);

AND2x2_ASAP7_75t_L g14936 ( 
.A(n_14588),
.B(n_14459),
.Y(n_14936)
);

INVx2_ASAP7_75t_L g14937 ( 
.A(n_14591),
.Y(n_14937)
);

INVx2_ASAP7_75t_SL g14938 ( 
.A(n_14506),
.Y(n_14938)
);

INVx3_ASAP7_75t_L g14939 ( 
.A(n_14728),
.Y(n_14939)
);

AND2x2_ASAP7_75t_L g14940 ( 
.A(n_14556),
.B(n_14461),
.Y(n_14940)
);

INVx2_ASAP7_75t_SL g14941 ( 
.A(n_14640),
.Y(n_14941)
);

BUFx3_ASAP7_75t_L g14942 ( 
.A(n_14523),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_14568),
.Y(n_14943)
);

INVx1_ASAP7_75t_L g14944 ( 
.A(n_14569),
.Y(n_14944)
);

INVx1_ASAP7_75t_L g14945 ( 
.A(n_14573),
.Y(n_14945)
);

INVx1_ASAP7_75t_L g14946 ( 
.A(n_14577),
.Y(n_14946)
);

INVx1_ASAP7_75t_L g14947 ( 
.A(n_14578),
.Y(n_14947)
);

INVx1_ASAP7_75t_L g14948 ( 
.A(n_14597),
.Y(n_14948)
);

INVx1_ASAP7_75t_L g14949 ( 
.A(n_14605),
.Y(n_14949)
);

INVx2_ASAP7_75t_L g14950 ( 
.A(n_14603),
.Y(n_14950)
);

INVx2_ASAP7_75t_L g14951 ( 
.A(n_14561),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14619),
.Y(n_14952)
);

AOI21xp5_ASAP7_75t_L g14953 ( 
.A1(n_14537),
.A2(n_14260),
.B(n_14258),
.Y(n_14953)
);

INVx2_ASAP7_75t_SL g14954 ( 
.A(n_14714),
.Y(n_14954)
);

OAI21x1_ASAP7_75t_L g14955 ( 
.A1(n_14599),
.A2(n_14480),
.B(n_14478),
.Y(n_14955)
);

INVx2_ASAP7_75t_L g14956 ( 
.A(n_14564),
.Y(n_14956)
);

AND2x4_ASAP7_75t_L g14957 ( 
.A(n_14624),
.B(n_14491),
.Y(n_14957)
);

AND2x4_ASAP7_75t_L g14958 ( 
.A(n_14796),
.B(n_14430),
.Y(n_14958)
);

INVx1_ASAP7_75t_L g14959 ( 
.A(n_14630),
.Y(n_14959)
);

AND2x4_ASAP7_75t_L g14960 ( 
.A(n_14532),
.B(n_14462),
.Y(n_14960)
);

INVx2_ASAP7_75t_L g14961 ( 
.A(n_14616),
.Y(n_14961)
);

INVx3_ASAP7_75t_L g14962 ( 
.A(n_14719),
.Y(n_14962)
);

OA21x2_ASAP7_75t_L g14963 ( 
.A1(n_14635),
.A2(n_14316),
.B(n_14268),
.Y(n_14963)
);

AO21x2_ASAP7_75t_L g14964 ( 
.A1(n_14846),
.A2(n_14494),
.B(n_2195),
.Y(n_14964)
);

HB1xp67_ASAP7_75t_L g14965 ( 
.A(n_14543),
.Y(n_14965)
);

INVx1_ASAP7_75t_L g14966 ( 
.A(n_14675),
.Y(n_14966)
);

BUFx2_ASAP7_75t_L g14967 ( 
.A(n_14581),
.Y(n_14967)
);

INVx1_ASAP7_75t_L g14968 ( 
.A(n_14740),
.Y(n_14968)
);

INVx2_ASAP7_75t_L g14969 ( 
.A(n_14660),
.Y(n_14969)
);

INVx2_ASAP7_75t_L g14970 ( 
.A(n_14518),
.Y(n_14970)
);

CKINVDCx6p67_ASAP7_75t_R g14971 ( 
.A(n_14582),
.Y(n_14971)
);

INVx1_ASAP7_75t_L g14972 ( 
.A(n_14653),
.Y(n_14972)
);

HB1xp67_ASAP7_75t_L g14973 ( 
.A(n_14749),
.Y(n_14973)
);

OAI21x1_ASAP7_75t_L g14974 ( 
.A1(n_14589),
.A2(n_2196),
.B(n_2197),
.Y(n_14974)
);

INVx1_ASAP7_75t_L g14975 ( 
.A(n_14671),
.Y(n_14975)
);

INVx2_ASAP7_75t_L g14976 ( 
.A(n_14765),
.Y(n_14976)
);

NOR2x1_ASAP7_75t_SL g14977 ( 
.A(n_14581),
.B(n_2198),
.Y(n_14977)
);

OAI21x1_ASAP7_75t_L g14978 ( 
.A1(n_14693),
.A2(n_2200),
.B(n_2201),
.Y(n_14978)
);

INVx2_ASAP7_75t_L g14979 ( 
.A(n_14735),
.Y(n_14979)
);

INVx1_ASAP7_75t_L g14980 ( 
.A(n_14751),
.Y(n_14980)
);

INVx1_ASAP7_75t_SL g14981 ( 
.A(n_14508),
.Y(n_14981)
);

AND2x2_ASAP7_75t_L g14982 ( 
.A(n_14517),
.B(n_2201),
.Y(n_14982)
);

BUFx6f_ASAP7_75t_L g14983 ( 
.A(n_14647),
.Y(n_14983)
);

INVx2_ASAP7_75t_L g14984 ( 
.A(n_14761),
.Y(n_14984)
);

OR2x2_ASAP7_75t_L g14985 ( 
.A(n_14705),
.B(n_2202),
.Y(n_14985)
);

INVx2_ASAP7_75t_L g14986 ( 
.A(n_14607),
.Y(n_14986)
);

OAI21x1_ASAP7_75t_L g14987 ( 
.A1(n_14618),
.A2(n_2202),
.B(n_2203),
.Y(n_14987)
);

INVx1_ASAP7_75t_L g14988 ( 
.A(n_14766),
.Y(n_14988)
);

NOR2xp33_ASAP7_75t_L g14989 ( 
.A(n_14709),
.B(n_2203),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14747),
.Y(n_14990)
);

INVx1_ASAP7_75t_L g14991 ( 
.A(n_14708),
.Y(n_14991)
);

INVx1_ASAP7_75t_L g14992 ( 
.A(n_14712),
.Y(n_14992)
);

INVxp33_ASAP7_75t_L g14993 ( 
.A(n_14571),
.Y(n_14993)
);

INVx2_ASAP7_75t_L g14994 ( 
.A(n_14579),
.Y(n_14994)
);

NAND2xp5_ASAP7_75t_L g14995 ( 
.A(n_14509),
.B(n_14575),
.Y(n_14995)
);

AOI21xp33_ASAP7_75t_L g14996 ( 
.A1(n_14566),
.A2(n_14510),
.B(n_14580),
.Y(n_14996)
);

INVx1_ASAP7_75t_L g14997 ( 
.A(n_14715),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14634),
.Y(n_14998)
);

INVx1_ASAP7_75t_L g14999 ( 
.A(n_14637),
.Y(n_14999)
);

INVx1_ASAP7_75t_L g15000 ( 
.A(n_14649),
.Y(n_15000)
);

INVx2_ASAP7_75t_L g15001 ( 
.A(n_14673),
.Y(n_15001)
);

INVx1_ASAP7_75t_L g15002 ( 
.A(n_14672),
.Y(n_15002)
);

INVx2_ASAP7_75t_L g15003 ( 
.A(n_14535),
.Y(n_15003)
);

HB1xp67_ASAP7_75t_L g15004 ( 
.A(n_14829),
.Y(n_15004)
);

AO21x2_ASAP7_75t_L g15005 ( 
.A1(n_14815),
.A2(n_2204),
.B(n_2205),
.Y(n_15005)
);

INVx1_ASAP7_75t_L g15006 ( 
.A(n_14823),
.Y(n_15006)
);

HB1xp67_ASAP7_75t_L g15007 ( 
.A(n_14562),
.Y(n_15007)
);

INVx2_ASAP7_75t_L g15008 ( 
.A(n_14797),
.Y(n_15008)
);

OAI21x1_ASAP7_75t_L g15009 ( 
.A1(n_14606),
.A2(n_2204),
.B(n_2205),
.Y(n_15009)
);

INVx3_ASAP7_75t_L g15010 ( 
.A(n_14714),
.Y(n_15010)
);

INVx1_ASAP7_75t_L g15011 ( 
.A(n_14833),
.Y(n_15011)
);

INVx2_ASAP7_75t_L g15012 ( 
.A(n_14797),
.Y(n_15012)
);

NAND2x1p5_ASAP7_75t_L g15013 ( 
.A(n_14559),
.B(n_2206),
.Y(n_15013)
);

OAI21x1_ASAP7_75t_L g15014 ( 
.A1(n_14734),
.A2(n_2206),
.B(n_2207),
.Y(n_15014)
);

INVx1_ASAP7_75t_SL g15015 ( 
.A(n_14799),
.Y(n_15015)
);

INVx3_ASAP7_75t_L g15016 ( 
.A(n_14676),
.Y(n_15016)
);

AND2x4_ASAP7_75t_L g15017 ( 
.A(n_14617),
.B(n_2208),
.Y(n_15017)
);

INVx4_ASAP7_75t_L g15018 ( 
.A(n_14826),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14834),
.Y(n_15019)
);

INVx1_ASAP7_75t_L g15020 ( 
.A(n_14685),
.Y(n_15020)
);

INVx2_ASAP7_75t_L g15021 ( 
.A(n_14724),
.Y(n_15021)
);

AND2x4_ASAP7_75t_L g15022 ( 
.A(n_14736),
.B(n_2208),
.Y(n_15022)
);

OR2x6_ASAP7_75t_L g15023 ( 
.A(n_14759),
.B(n_14558),
.Y(n_15023)
);

CKINVDCx5p33_ASAP7_75t_R g15024 ( 
.A(n_14730),
.Y(n_15024)
);

AO31x2_ASAP7_75t_L g15025 ( 
.A1(n_14777),
.A2(n_2211),
.A3(n_2209),
.B(n_2210),
.Y(n_15025)
);

INVx2_ASAP7_75t_L g15026 ( 
.A(n_14501),
.Y(n_15026)
);

INVx2_ASAP7_75t_L g15027 ( 
.A(n_14825),
.Y(n_15027)
);

BUFx6f_ASAP7_75t_L g15028 ( 
.A(n_14602),
.Y(n_15028)
);

INVx1_ASAP7_75t_L g15029 ( 
.A(n_14692),
.Y(n_15029)
);

OAI21x1_ASAP7_75t_L g15030 ( 
.A1(n_14655),
.A2(n_2210),
.B(n_2211),
.Y(n_15030)
);

AO21x1_ASAP7_75t_SL g15031 ( 
.A1(n_14890),
.A2(n_2212),
.B(n_2213),
.Y(n_15031)
);

INVx1_ASAP7_75t_L g15032 ( 
.A(n_14698),
.Y(n_15032)
);

INVx2_ASAP7_75t_SL g15033 ( 
.A(n_14776),
.Y(n_15033)
);

AOI222xp33_ASAP7_75t_L g15034 ( 
.A1(n_14773),
.A2(n_2215),
.B1(n_2217),
.B2(n_2212),
.C1(n_2214),
.C2(n_2216),
.Y(n_15034)
);

HB1xp67_ASAP7_75t_L g15035 ( 
.A(n_14683),
.Y(n_15035)
);

OAI211xp5_ASAP7_75t_L g15036 ( 
.A1(n_14746),
.A2(n_2217),
.B(n_2214),
.C(n_2215),
.Y(n_15036)
);

INVx1_ASAP7_75t_L g15037 ( 
.A(n_14800),
.Y(n_15037)
);

AND2x4_ASAP7_75t_L g15038 ( 
.A(n_14741),
.B(n_2218),
.Y(n_15038)
);

INVx2_ASAP7_75t_L g15039 ( 
.A(n_14583),
.Y(n_15039)
);

INVx1_ASAP7_75t_L g15040 ( 
.A(n_14805),
.Y(n_15040)
);

INVx2_ASAP7_75t_L g15041 ( 
.A(n_14583),
.Y(n_15041)
);

INVx2_ASAP7_75t_L g15042 ( 
.A(n_14531),
.Y(n_15042)
);

INVx1_ASAP7_75t_L g15043 ( 
.A(n_14636),
.Y(n_15043)
);

INVx1_ASAP7_75t_L g15044 ( 
.A(n_14652),
.Y(n_15044)
);

INVx1_ASAP7_75t_L g15045 ( 
.A(n_14657),
.Y(n_15045)
);

NAND2x1p5_ASAP7_75t_L g15046 ( 
.A(n_14860),
.B(n_2218),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_14670),
.Y(n_15047)
);

INVx1_ASAP7_75t_L g15048 ( 
.A(n_14732),
.Y(n_15048)
);

NAND2x1p5_ASAP7_75t_L g15049 ( 
.A(n_14770),
.B(n_14859),
.Y(n_15049)
);

NAND2xp5_ASAP7_75t_L g15050 ( 
.A(n_14594),
.B(n_14576),
.Y(n_15050)
);

INVx1_ASAP7_75t_L g15051 ( 
.A(n_14662),
.Y(n_15051)
);

AO21x2_ASAP7_75t_L g15052 ( 
.A1(n_14702),
.A2(n_2219),
.B(n_2220),
.Y(n_15052)
);

O2A1O1Ixp33_ASAP7_75t_L g15053 ( 
.A1(n_14707),
.A2(n_2221),
.B(n_2219),
.C(n_2220),
.Y(n_15053)
);

INVx2_ASAP7_75t_L g15054 ( 
.A(n_14500),
.Y(n_15054)
);

INVx2_ASAP7_75t_SL g15055 ( 
.A(n_14586),
.Y(n_15055)
);

INVxp67_ASAP7_75t_L g15056 ( 
.A(n_14801),
.Y(n_15056)
);

INVx1_ASAP7_75t_L g15057 ( 
.A(n_14706),
.Y(n_15057)
);

INVx1_ASAP7_75t_L g15058 ( 
.A(n_14742),
.Y(n_15058)
);

INVx2_ASAP7_75t_L g15059 ( 
.A(n_14849),
.Y(n_15059)
);

AND2x4_ASAP7_75t_L g15060 ( 
.A(n_14507),
.B(n_2221),
.Y(n_15060)
);

INVx2_ASAP7_75t_SL g15061 ( 
.A(n_14830),
.Y(n_15061)
);

INVx2_ASAP7_75t_L g15062 ( 
.A(n_14529),
.Y(n_15062)
);

INVx2_ASAP7_75t_L g15063 ( 
.A(n_14659),
.Y(n_15063)
);

NAND2xp5_ASAP7_75t_L g15064 ( 
.A(n_14840),
.B(n_14841),
.Y(n_15064)
);

NOR2xp33_ASAP7_75t_SL g15065 ( 
.A(n_14590),
.B(n_2223),
.Y(n_15065)
);

INVx1_ASAP7_75t_L g15066 ( 
.A(n_14625),
.Y(n_15066)
);

INVx1_ASAP7_75t_L g15067 ( 
.A(n_14674),
.Y(n_15067)
);

NAND2xp5_ASAP7_75t_L g15068 ( 
.A(n_14844),
.B(n_2223),
.Y(n_15068)
);

OAI21x1_ASAP7_75t_L g15069 ( 
.A1(n_14620),
.A2(n_2225),
.B(n_2226),
.Y(n_15069)
);

INVx1_ASAP7_75t_L g15070 ( 
.A(n_14869),
.Y(n_15070)
);

INVx1_ASAP7_75t_L g15071 ( 
.A(n_14633),
.Y(n_15071)
);

INVx1_ASAP7_75t_L g15072 ( 
.A(n_14633),
.Y(n_15072)
);

INVx1_ASAP7_75t_L g15073 ( 
.A(n_14684),
.Y(n_15073)
);

NOR2x1_ASAP7_75t_R g15074 ( 
.A(n_14816),
.B(n_2225),
.Y(n_15074)
);

INVx1_ASAP7_75t_L g15075 ( 
.A(n_14545),
.Y(n_15075)
);

AND2x2_ASAP7_75t_L g15076 ( 
.A(n_14574),
.B(n_2226),
.Y(n_15076)
);

AO21x2_ASAP7_75t_L g15077 ( 
.A1(n_14852),
.A2(n_2227),
.B(n_2228),
.Y(n_15077)
);

INVx1_ASAP7_75t_L g15078 ( 
.A(n_14646),
.Y(n_15078)
);

HB1xp67_ASAP7_75t_L g15079 ( 
.A(n_14546),
.Y(n_15079)
);

INVx1_ASAP7_75t_L g15080 ( 
.A(n_14793),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_14868),
.Y(n_15081)
);

BUFx3_ASAP7_75t_L g15082 ( 
.A(n_14810),
.Y(n_15082)
);

INVx1_ASAP7_75t_L g15083 ( 
.A(n_14874),
.Y(n_15083)
);

INVx1_ASAP7_75t_L g15084 ( 
.A(n_14880),
.Y(n_15084)
);

INVx3_ASAP7_75t_L g15085 ( 
.A(n_14511),
.Y(n_15085)
);

INVx2_ASAP7_75t_L g15086 ( 
.A(n_14887),
.Y(n_15086)
);

AND2x2_ASAP7_75t_L g15087 ( 
.A(n_14598),
.B(n_14756),
.Y(n_15087)
);

AND2x2_ASAP7_75t_L g15088 ( 
.A(n_14739),
.B(n_14855),
.Y(n_15088)
);

NOR2x1_ASAP7_75t_L g15089 ( 
.A(n_14809),
.B(n_2227),
.Y(n_15089)
);

INVx2_ASAP7_75t_L g15090 ( 
.A(n_14887),
.Y(n_15090)
);

OR2x6_ASAP7_75t_L g15091 ( 
.A(n_14804),
.B(n_2228),
.Y(n_15091)
);

INVx2_ASAP7_75t_SL g15092 ( 
.A(n_14824),
.Y(n_15092)
);

INVx1_ASAP7_75t_L g15093 ( 
.A(n_14861),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_14883),
.Y(n_15094)
);

AND2x2_ASAP7_75t_L g15095 ( 
.A(n_14610),
.B(n_2229),
.Y(n_15095)
);

NAND2xp5_ASAP7_75t_L g15096 ( 
.A(n_14848),
.B(n_14850),
.Y(n_15096)
);

OR2x2_ASAP7_75t_L g15097 ( 
.A(n_14572),
.B(n_2229),
.Y(n_15097)
);

AND2x2_ASAP7_75t_L g15098 ( 
.A(n_14614),
.B(n_14878),
.Y(n_15098)
);

HB1xp67_ASAP7_75t_L g15099 ( 
.A(n_14548),
.Y(n_15099)
);

INVx1_ASAP7_75t_L g15100 ( 
.A(n_14891),
.Y(n_15100)
);

INVx2_ASAP7_75t_L g15101 ( 
.A(n_14519),
.Y(n_15101)
);

A2O1A1Ixp33_ASAP7_75t_SL g15102 ( 
.A1(n_14666),
.A2(n_2232),
.B(n_2230),
.C(n_2231),
.Y(n_15102)
);

INVx1_ASAP7_75t_L g15103 ( 
.A(n_14723),
.Y(n_15103)
);

NAND2xp5_ASAP7_75t_L g15104 ( 
.A(n_14851),
.B(n_2230),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_14882),
.Y(n_15105)
);

INVx1_ASAP7_75t_L g15106 ( 
.A(n_14689),
.Y(n_15106)
);

AOI22xp33_ASAP7_75t_L g15107 ( 
.A1(n_14648),
.A2(n_2234),
.B1(n_2231),
.B2(n_2233),
.Y(n_15107)
);

INVx2_ASAP7_75t_L g15108 ( 
.A(n_14843),
.Y(n_15108)
);

INVx2_ASAP7_75t_L g15109 ( 
.A(n_14567),
.Y(n_15109)
);

INVx2_ASAP7_75t_L g15110 ( 
.A(n_14601),
.Y(n_15110)
);

INVx1_ASAP7_75t_L g15111 ( 
.A(n_14786),
.Y(n_15111)
);

OR2x2_ASAP7_75t_L g15112 ( 
.A(n_14563),
.B(n_2233),
.Y(n_15112)
);

INVx1_ASAP7_75t_L g15113 ( 
.A(n_14803),
.Y(n_15113)
);

INVx1_ASAP7_75t_L g15114 ( 
.A(n_14807),
.Y(n_15114)
);

INVx1_ASAP7_75t_L g15115 ( 
.A(n_14627),
.Y(n_15115)
);

AND2x2_ASAP7_75t_L g15116 ( 
.A(n_14886),
.B(n_2234),
.Y(n_15116)
);

OAI22xp33_ASAP7_75t_L g15117 ( 
.A1(n_14731),
.A2(n_2237),
.B1(n_2235),
.B2(n_2236),
.Y(n_15117)
);

INVx3_ASAP7_75t_L g15118 ( 
.A(n_14824),
.Y(n_15118)
);

INVx1_ASAP7_75t_L g15119 ( 
.A(n_14682),
.Y(n_15119)
);

INVx1_ASAP7_75t_L g15120 ( 
.A(n_14757),
.Y(n_15120)
);

CKINVDCx6p67_ASAP7_75t_R g15121 ( 
.A(n_14565),
.Y(n_15121)
);

NOR2xp33_ASAP7_75t_L g15122 ( 
.A(n_14547),
.B(n_2236),
.Y(n_15122)
);

OA21x2_ASAP7_75t_L g15123 ( 
.A1(n_14613),
.A2(n_2237),
.B(n_2238),
.Y(n_15123)
);

BUFx3_ASAP7_75t_L g15124 ( 
.A(n_14661),
.Y(n_15124)
);

INVx2_ASAP7_75t_L g15125 ( 
.A(n_14604),
.Y(n_15125)
);

CKINVDCx20_ASAP7_75t_R g15126 ( 
.A(n_14788),
.Y(n_15126)
);

INVx3_ASAP7_75t_L g15127 ( 
.A(n_14542),
.Y(n_15127)
);

BUFx3_ASAP7_75t_L g15128 ( 
.A(n_14718),
.Y(n_15128)
);

AND2x2_ASAP7_75t_L g15129 ( 
.A(n_14551),
.B(n_2239),
.Y(n_15129)
);

INVx1_ASAP7_75t_L g15130 ( 
.A(n_14784),
.Y(n_15130)
);

NAND4xp25_ASAP7_75t_SL g15131 ( 
.A(n_14592),
.B(n_2241),
.C(n_2239),
.D(n_2240),
.Y(n_15131)
);

CKINVDCx5p33_ASAP7_75t_R g15132 ( 
.A(n_14827),
.Y(n_15132)
);

INVx1_ASAP7_75t_L g15133 ( 
.A(n_14828),
.Y(n_15133)
);

INVx2_ASAP7_75t_L g15134 ( 
.A(n_14716),
.Y(n_15134)
);

HB1xp67_ASAP7_75t_L g15135 ( 
.A(n_14516),
.Y(n_15135)
);

OR2x2_ASAP7_75t_L g15136 ( 
.A(n_14515),
.B(n_2240),
.Y(n_15136)
);

BUFx2_ASAP7_75t_L g15137 ( 
.A(n_14565),
.Y(n_15137)
);

CKINVDCx20_ASAP7_75t_R g15138 ( 
.A(n_14542),
.Y(n_15138)
);

BUFx3_ASAP7_75t_L g15139 ( 
.A(n_14722),
.Y(n_15139)
);

INVx1_ASAP7_75t_L g15140 ( 
.A(n_14767),
.Y(n_15140)
);

INVx2_ASAP7_75t_SL g15141 ( 
.A(n_14669),
.Y(n_15141)
);

BUFx3_ASAP7_75t_L g15142 ( 
.A(n_14775),
.Y(n_15142)
);

INVx1_ASAP7_75t_L g15143 ( 
.A(n_14889),
.Y(n_15143)
);

HB1xp67_ASAP7_75t_L g15144 ( 
.A(n_14780),
.Y(n_15144)
);

INVx2_ASAP7_75t_L g15145 ( 
.A(n_14856),
.Y(n_15145)
);

INVx1_ASAP7_75t_L g15146 ( 
.A(n_14798),
.Y(n_15146)
);

INVx2_ASAP7_75t_L g15147 ( 
.A(n_14791),
.Y(n_15147)
);

BUFx2_ASAP7_75t_L g15148 ( 
.A(n_14565),
.Y(n_15148)
);

OA21x2_ASAP7_75t_L g15149 ( 
.A1(n_14842),
.A2(n_2241),
.B(n_2242),
.Y(n_15149)
);

INVx1_ASAP7_75t_L g15150 ( 
.A(n_14783),
.Y(n_15150)
);

INVx1_ASAP7_75t_L g15151 ( 
.A(n_14764),
.Y(n_15151)
);

BUFx2_ASAP7_75t_L g15152 ( 
.A(n_14854),
.Y(n_15152)
);

INVx1_ASAP7_75t_L g15153 ( 
.A(n_14772),
.Y(n_15153)
);

BUFx8_ASAP7_75t_SL g15154 ( 
.A(n_14814),
.Y(n_15154)
);

INVx1_ASAP7_75t_L g15155 ( 
.A(n_14778),
.Y(n_15155)
);

INVx1_ASAP7_75t_L g15156 ( 
.A(n_14782),
.Y(n_15156)
);

INVx2_ASAP7_75t_L g15157 ( 
.A(n_14792),
.Y(n_15157)
);

INVx1_ASAP7_75t_L g15158 ( 
.A(n_14641),
.Y(n_15158)
);

HB1xp67_ASAP7_75t_L g15159 ( 
.A(n_14885),
.Y(n_15159)
);

INVx1_ASAP7_75t_L g15160 ( 
.A(n_14871),
.Y(n_15160)
);

INVx2_ASAP7_75t_L g15161 ( 
.A(n_14526),
.Y(n_15161)
);

OAI21x1_ASAP7_75t_L g15162 ( 
.A1(n_14615),
.A2(n_2242),
.B(n_2243),
.Y(n_15162)
);

INVx1_ASAP7_75t_L g15163 ( 
.A(n_14612),
.Y(n_15163)
);

INVx1_ASAP7_75t_L g15164 ( 
.A(n_14651),
.Y(n_15164)
);

INVx4_ASAP7_75t_SL g15165 ( 
.A(n_14750),
.Y(n_15165)
);

INVx1_ASAP7_75t_L g15166 ( 
.A(n_14858),
.Y(n_15166)
);

OAI21x1_ASAP7_75t_L g15167 ( 
.A1(n_14541),
.A2(n_2243),
.B(n_2244),
.Y(n_15167)
);

AND2x2_ASAP7_75t_L g15168 ( 
.A(n_14522),
.B(n_2245),
.Y(n_15168)
);

AND2x4_ASAP7_75t_L g15169 ( 
.A(n_14628),
.B(n_14758),
.Y(n_15169)
);

INVx1_ASAP7_75t_L g15170 ( 
.A(n_14853),
.Y(n_15170)
);

AND2x2_ASAP7_75t_L g15171 ( 
.A(n_14608),
.B(n_2246),
.Y(n_15171)
);

INVx1_ASAP7_75t_L g15172 ( 
.A(n_14753),
.Y(n_15172)
);

AND2x4_ASAP7_75t_L g15173 ( 
.A(n_14820),
.B(n_2246),
.Y(n_15173)
);

BUFx3_ASAP7_75t_L g15174 ( 
.A(n_14700),
.Y(n_15174)
);

INVx2_ASAP7_75t_L g15175 ( 
.A(n_14555),
.Y(n_15175)
);

INVx2_ASAP7_75t_L g15176 ( 
.A(n_14549),
.Y(n_15176)
);

INVx1_ASAP7_75t_L g15177 ( 
.A(n_14872),
.Y(n_15177)
);

INVx2_ASAP7_75t_L g15178 ( 
.A(n_14769),
.Y(n_15178)
);

INVx1_ASAP7_75t_L g15179 ( 
.A(n_14818),
.Y(n_15179)
);

INVx2_ASAP7_75t_L g15180 ( 
.A(n_14626),
.Y(n_15180)
);

OAI21xp5_ASAP7_75t_L g15181 ( 
.A1(n_14557),
.A2(n_2247),
.B(n_2248),
.Y(n_15181)
);

INVx1_ASAP7_75t_L g15182 ( 
.A(n_14836),
.Y(n_15182)
);

HB1xp67_ASAP7_75t_L g15183 ( 
.A(n_14738),
.Y(n_15183)
);

OAI21x1_ASAP7_75t_L g15184 ( 
.A1(n_14584),
.A2(n_2247),
.B(n_2248),
.Y(n_15184)
);

INVx2_ASAP7_75t_L g15185 ( 
.A(n_14521),
.Y(n_15185)
);

INVx1_ASAP7_75t_L g15186 ( 
.A(n_14642),
.Y(n_15186)
);

BUFx3_ASAP7_75t_L g15187 ( 
.A(n_14822),
.Y(n_15187)
);

INVx2_ASAP7_75t_L g15188 ( 
.A(n_14527),
.Y(n_15188)
);

INVx1_ASAP7_75t_L g15189 ( 
.A(n_14680),
.Y(n_15189)
);

INVx2_ASAP7_75t_SL g15190 ( 
.A(n_14639),
.Y(n_15190)
);

HB1xp67_ASAP7_75t_L g15191 ( 
.A(n_14528),
.Y(n_15191)
);

BUFx2_ASAP7_75t_L g15192 ( 
.A(n_14503),
.Y(n_15192)
);

AO21x1_ASAP7_75t_L g15193 ( 
.A1(n_14888),
.A2(n_2249),
.B(n_2250),
.Y(n_15193)
);

INVx2_ASAP7_75t_L g15194 ( 
.A(n_14748),
.Y(n_15194)
);

AND2x4_ASAP7_75t_L g15195 ( 
.A(n_14677),
.B(n_2249),
.Y(n_15195)
);

BUFx10_ASAP7_75t_L g15196 ( 
.A(n_14686),
.Y(n_15196)
);

INVx2_ASAP7_75t_L g15197 ( 
.A(n_14701),
.Y(n_15197)
);

HB1xp67_ASAP7_75t_L g15198 ( 
.A(n_14876),
.Y(n_15198)
);

NAND2xp5_ASAP7_75t_L g15199 ( 
.A(n_14631),
.B(n_14650),
.Y(n_15199)
);

NAND2xp5_ASAP7_75t_L g15200 ( 
.A(n_14656),
.B(n_14632),
.Y(n_15200)
);

OR2x2_ASAP7_75t_L g15201 ( 
.A(n_14585),
.B(n_2251),
.Y(n_15201)
);

INVx1_ASAP7_75t_L g15202 ( 
.A(n_14710),
.Y(n_15202)
);

BUFx2_ASAP7_75t_SL g15203 ( 
.A(n_14774),
.Y(n_15203)
);

INVx2_ASAP7_75t_L g15204 ( 
.A(n_14726),
.Y(n_15204)
);

INVx1_ASAP7_75t_L g15205 ( 
.A(n_14644),
.Y(n_15205)
);

HB1xp67_ASAP7_75t_L g15206 ( 
.A(n_14729),
.Y(n_15206)
);

AND2x2_ASAP7_75t_L g15207 ( 
.A(n_14745),
.B(n_2251),
.Y(n_15207)
);

AND2x4_ASAP7_75t_L g15208 ( 
.A(n_14762),
.B(n_2252),
.Y(n_15208)
);

INVx1_ASAP7_75t_L g15209 ( 
.A(n_14787),
.Y(n_15209)
);

INVx1_ASAP7_75t_L g15210 ( 
.A(n_14725),
.Y(n_15210)
);

INVx2_ASAP7_75t_L g15211 ( 
.A(n_14694),
.Y(n_15211)
);

AND2x4_ASAP7_75t_L g15212 ( 
.A(n_14763),
.B(n_14771),
.Y(n_15212)
);

BUFx2_ASAP7_75t_L g15213 ( 
.A(n_14678),
.Y(n_15213)
);

INVx1_ASAP7_75t_L g15214 ( 
.A(n_14727),
.Y(n_15214)
);

INVx1_ASAP7_75t_L g15215 ( 
.A(n_14881),
.Y(n_15215)
);

INVx1_ASAP7_75t_L g15216 ( 
.A(n_14658),
.Y(n_15216)
);

NAND2xp5_ASAP7_75t_L g15217 ( 
.A(n_14663),
.B(n_2252),
.Y(n_15217)
);

NAND2xp5_ASAP7_75t_L g15218 ( 
.A(n_14691),
.B(n_2253),
.Y(n_15218)
);

AND2x2_ASAP7_75t_L g15219 ( 
.A(n_14713),
.B(n_2253),
.Y(n_15219)
);

BUFx4f_ASAP7_75t_SL g15220 ( 
.A(n_14645),
.Y(n_15220)
);

INVx1_ASAP7_75t_L g15221 ( 
.A(n_14593),
.Y(n_15221)
);

INVx2_ASAP7_75t_L g15222 ( 
.A(n_14884),
.Y(n_15222)
);

HB1xp67_ASAP7_75t_L g15223 ( 
.A(n_14711),
.Y(n_15223)
);

INVx1_ASAP7_75t_L g15224 ( 
.A(n_14743),
.Y(n_15224)
);

AOI22xp5_ASAP7_75t_L g15225 ( 
.A1(n_14755),
.A2(n_2256),
.B1(n_2254),
.B2(n_2255),
.Y(n_15225)
);

INVx3_ASAP7_75t_L g15226 ( 
.A(n_14847),
.Y(n_15226)
);

INVx1_ASAP7_75t_L g15227 ( 
.A(n_14743),
.Y(n_15227)
);

INVx3_ASAP7_75t_L g15228 ( 
.A(n_14838),
.Y(n_15228)
);

INVx2_ASAP7_75t_L g15229 ( 
.A(n_14808),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_14733),
.Y(n_15230)
);

NOR2xp67_ASAP7_75t_L g15231 ( 
.A(n_14877),
.B(n_2254),
.Y(n_15231)
);

INVx1_ASAP7_75t_L g15232 ( 
.A(n_14654),
.Y(n_15232)
);

BUFx2_ASAP7_75t_L g15233 ( 
.A(n_14845),
.Y(n_15233)
);

INVx2_ASAP7_75t_L g15234 ( 
.A(n_14622),
.Y(n_15234)
);

INVx2_ASAP7_75t_L g15235 ( 
.A(n_14873),
.Y(n_15235)
);

INVx2_ASAP7_75t_L g15236 ( 
.A(n_14867),
.Y(n_15236)
);

INVx2_ASAP7_75t_L g15237 ( 
.A(n_14839),
.Y(n_15237)
);

NAND2xp5_ASAP7_75t_L g15238 ( 
.A(n_14595),
.B(n_2255),
.Y(n_15238)
);

INVxp33_ASAP7_75t_SL g15239 ( 
.A(n_14643),
.Y(n_15239)
);

BUFx3_ASAP7_75t_L g15240 ( 
.A(n_14831),
.Y(n_15240)
);

OA21x2_ASAP7_75t_L g15241 ( 
.A1(n_14697),
.A2(n_14502),
.B(n_14587),
.Y(n_15241)
);

AND2x2_ASAP7_75t_L g15242 ( 
.A(n_14813),
.B(n_2256),
.Y(n_15242)
);

BUFx6f_ASAP7_75t_L g15243 ( 
.A(n_14752),
.Y(n_15243)
);

INVx2_ASAP7_75t_SL g15244 ( 
.A(n_14781),
.Y(n_15244)
);

INVx1_ASAP7_75t_L g15245 ( 
.A(n_14654),
.Y(n_15245)
);

AO21x2_ASAP7_75t_L g15246 ( 
.A1(n_14821),
.A2(n_2257),
.B(n_2258),
.Y(n_15246)
);

BUFx3_ASAP7_75t_L g15247 ( 
.A(n_14790),
.Y(n_15247)
);

OR2x2_ASAP7_75t_L g15248 ( 
.A(n_14819),
.B(n_2259),
.Y(n_15248)
);

AND2x2_ASAP7_75t_L g15249 ( 
.A(n_14835),
.B(n_2259),
.Y(n_15249)
);

INVx2_ASAP7_75t_L g15250 ( 
.A(n_14879),
.Y(n_15250)
);

AND2x2_ASAP7_75t_L g15251 ( 
.A(n_14717),
.B(n_2260),
.Y(n_15251)
);

INVx2_ASAP7_75t_L g15252 ( 
.A(n_14629),
.Y(n_15252)
);

INVx2_ASAP7_75t_SL g15253 ( 
.A(n_14785),
.Y(n_15253)
);

NAND2xp5_ASAP7_75t_L g15254 ( 
.A(n_14750),
.B(n_2261),
.Y(n_15254)
);

INVx1_ASAP7_75t_L g15255 ( 
.A(n_14875),
.Y(n_15255)
);

NAND2xp5_ASAP7_75t_L g15256 ( 
.A(n_15244),
.B(n_14687),
.Y(n_15256)
);

AOI22xp33_ASAP7_75t_SL g15257 ( 
.A1(n_14923),
.A2(n_14664),
.B1(n_14863),
.B2(n_14621),
.Y(n_15257)
);

INVx2_ASAP7_75t_L g15258 ( 
.A(n_14983),
.Y(n_15258)
);

AOI22xp33_ASAP7_75t_L g15259 ( 
.A1(n_14996),
.A2(n_14857),
.B1(n_14811),
.B2(n_14754),
.Y(n_15259)
);

BUFx3_ASAP7_75t_L g15260 ( 
.A(n_14900),
.Y(n_15260)
);

OAI221xp5_ASAP7_75t_L g15261 ( 
.A1(n_15181),
.A2(n_14794),
.B1(n_14665),
.B2(n_14760),
.C(n_14699),
.Y(n_15261)
);

INVx1_ASAP7_75t_L g15262 ( 
.A(n_14965),
.Y(n_15262)
);

OAI221xp5_ASAP7_75t_L g15263 ( 
.A1(n_14995),
.A2(n_14865),
.B1(n_14688),
.B2(n_14721),
.C(n_14668),
.Y(n_15263)
);

AOI22xp33_ASAP7_75t_L g15264 ( 
.A1(n_14916),
.A2(n_14795),
.B1(n_14892),
.B2(n_14812),
.Y(n_15264)
);

INVx2_ASAP7_75t_SL g15265 ( 
.A(n_14918),
.Y(n_15265)
);

CKINVDCx6p67_ASAP7_75t_R g15266 ( 
.A(n_14925),
.Y(n_15266)
);

AOI22xp33_ASAP7_75t_SL g15267 ( 
.A1(n_15241),
.A2(n_15192),
.B1(n_15050),
.B2(n_15213),
.Y(n_15267)
);

AOI221xp5_ASAP7_75t_L g15268 ( 
.A1(n_14953),
.A2(n_15183),
.B1(n_15206),
.B2(n_15117),
.C(n_15223),
.Y(n_15268)
);

NAND2xp5_ASAP7_75t_L g15269 ( 
.A(n_15203),
.B(n_14862),
.Y(n_15269)
);

AND2x2_ASAP7_75t_L g15270 ( 
.A(n_15127),
.B(n_14866),
.Y(n_15270)
);

OAI221xp5_ASAP7_75t_L g15271 ( 
.A1(n_14933),
.A2(n_14623),
.B1(n_14832),
.B2(n_14870),
.C(n_14779),
.Y(n_15271)
);

OAI22xp5_ASAP7_75t_L g15272 ( 
.A1(n_15199),
.A2(n_14789),
.B1(n_14744),
.B2(n_14696),
.Y(n_15272)
);

AOI21xp33_ASAP7_75t_L g15273 ( 
.A1(n_14993),
.A2(n_14806),
.B(n_14875),
.Y(n_15273)
);

INVx1_ASAP7_75t_L g15274 ( 
.A(n_14910),
.Y(n_15274)
);

AOI221xp5_ASAP7_75t_L g15275 ( 
.A1(n_15131),
.A2(n_14802),
.B1(n_14837),
.B2(n_2264),
.C(n_2262),
.Y(n_15275)
);

HB1xp67_ASAP7_75t_L g15276 ( 
.A(n_15198),
.Y(n_15276)
);

AOI222xp33_ASAP7_75t_L g15277 ( 
.A1(n_15200),
.A2(n_14802),
.B1(n_14837),
.B2(n_2264),
.C1(n_2266),
.C2(n_2262),
.Y(n_15277)
);

INVx2_ASAP7_75t_L g15278 ( 
.A(n_14983),
.Y(n_15278)
);

INVx1_ASAP7_75t_SL g15279 ( 
.A(n_15220),
.Y(n_15279)
);

INVx2_ASAP7_75t_L g15280 ( 
.A(n_14911),
.Y(n_15280)
);

AND2x4_ASAP7_75t_L g15281 ( 
.A(n_14938),
.B(n_2263),
.Y(n_15281)
);

A2O1A1Ixp33_ASAP7_75t_L g15282 ( 
.A1(n_15231),
.A2(n_2266),
.B(n_2263),
.C(n_2265),
.Y(n_15282)
);

AOI22xp33_ASAP7_75t_L g15283 ( 
.A1(n_14963),
.A2(n_2268),
.B1(n_2265),
.B2(n_2267),
.Y(n_15283)
);

OR2x6_ASAP7_75t_L g15284 ( 
.A(n_15137),
.B(n_2267),
.Y(n_15284)
);

INVx1_ASAP7_75t_L g15285 ( 
.A(n_15037),
.Y(n_15285)
);

NAND3xp33_ASAP7_75t_L g15286 ( 
.A(n_14973),
.B(n_15004),
.C(n_14932),
.Y(n_15286)
);

BUFx4f_ASAP7_75t_SL g15287 ( 
.A(n_15138),
.Y(n_15287)
);

AND2x2_ASAP7_75t_L g15288 ( 
.A(n_14967),
.B(n_14897),
.Y(n_15288)
);

AND2x2_ASAP7_75t_L g15289 ( 
.A(n_14908),
.B(n_2268),
.Y(n_15289)
);

NAND2xp5_ASAP7_75t_L g15290 ( 
.A(n_14896),
.B(n_2269),
.Y(n_15290)
);

OAI211xp5_ASAP7_75t_SL g15291 ( 
.A1(n_14922),
.A2(n_15111),
.B(n_15036),
.C(n_15120),
.Y(n_15291)
);

INVx1_ASAP7_75t_L g15292 ( 
.A(n_15040),
.Y(n_15292)
);

AOI21xp5_ASAP7_75t_L g15293 ( 
.A1(n_14894),
.A2(n_2269),
.B(n_2270),
.Y(n_15293)
);

OR2x2_ASAP7_75t_L g15294 ( 
.A(n_14926),
.B(n_2272),
.Y(n_15294)
);

AOI22xp33_ASAP7_75t_SL g15295 ( 
.A1(n_15236),
.A2(n_2274),
.B1(n_2272),
.B2(n_2273),
.Y(n_15295)
);

CKINVDCx20_ASAP7_75t_R g15296 ( 
.A(n_15024),
.Y(n_15296)
);

OAI22xp5_ASAP7_75t_L g15297 ( 
.A1(n_15237),
.A2(n_2275),
.B1(n_2273),
.B2(n_2274),
.Y(n_15297)
);

AOI22xp5_ASAP7_75t_L g15298 ( 
.A1(n_15193),
.A2(n_2278),
.B1(n_2276),
.B2(n_2277),
.Y(n_15298)
);

INVx1_ASAP7_75t_L g15299 ( 
.A(n_15007),
.Y(n_15299)
);

OAI22xp5_ASAP7_75t_L g15300 ( 
.A1(n_14901),
.A2(n_2278),
.B1(n_2276),
.B2(n_2277),
.Y(n_15300)
);

OAI211xp5_ASAP7_75t_L g15301 ( 
.A1(n_15053),
.A2(n_2281),
.B(n_2279),
.C(n_2280),
.Y(n_15301)
);

AND2x2_ASAP7_75t_L g15302 ( 
.A(n_15148),
.B(n_2279),
.Y(n_15302)
);

OAI221xp5_ASAP7_75t_L g15303 ( 
.A1(n_15023),
.A2(n_2283),
.B1(n_2280),
.B2(n_2282),
.C(n_2284),
.Y(n_15303)
);

AND2x2_ASAP7_75t_L g15304 ( 
.A(n_14915),
.B(n_2283),
.Y(n_15304)
);

AOI22xp33_ASAP7_75t_L g15305 ( 
.A1(n_14971),
.A2(n_2287),
.B1(n_2285),
.B2(n_2286),
.Y(n_15305)
);

OAI22xp5_ASAP7_75t_L g15306 ( 
.A1(n_15057),
.A2(n_2288),
.B1(n_2285),
.B2(n_2286),
.Y(n_15306)
);

AOI22xp33_ASAP7_75t_L g15307 ( 
.A1(n_14899),
.A2(n_2290),
.B1(n_2288),
.B2(n_2289),
.Y(n_15307)
);

AND2x2_ASAP7_75t_L g15308 ( 
.A(n_15021),
.B(n_14942),
.Y(n_15308)
);

AND2x2_ASAP7_75t_L g15309 ( 
.A(n_14981),
.B(n_2289),
.Y(n_15309)
);

OR2x2_ASAP7_75t_L g15310 ( 
.A(n_15209),
.B(n_2290),
.Y(n_15310)
);

AOI22xp33_ASAP7_75t_SL g15311 ( 
.A1(n_15239),
.A2(n_2293),
.B1(n_2291),
.B2(n_2292),
.Y(n_15311)
);

OAI21x1_ASAP7_75t_L g15312 ( 
.A1(n_14895),
.A2(n_2291),
.B(n_2292),
.Y(n_15312)
);

AND2x2_ASAP7_75t_L g15313 ( 
.A(n_15226),
.B(n_15152),
.Y(n_15313)
);

INVx1_ASAP7_75t_L g15314 ( 
.A(n_15058),
.Y(n_15314)
);

NAND2xp33_ASAP7_75t_R g15315 ( 
.A(n_15123),
.B(n_2293),
.Y(n_15315)
);

NOR3xp33_ASAP7_75t_L g15316 ( 
.A(n_14927),
.B(n_2294),
.C(n_2295),
.Y(n_15316)
);

AOI221xp5_ASAP7_75t_L g15317 ( 
.A1(n_15066),
.A2(n_2296),
.B1(n_2294),
.B2(n_2295),
.C(n_2297),
.Y(n_15317)
);

BUFx6f_ASAP7_75t_L g15318 ( 
.A(n_15028),
.Y(n_15318)
);

AND2x2_ASAP7_75t_L g15319 ( 
.A(n_14962),
.B(n_2296),
.Y(n_15319)
);

OAI221xp5_ASAP7_75t_L g15320 ( 
.A1(n_15023),
.A2(n_2299),
.B1(n_2297),
.B2(n_2298),
.C(n_2300),
.Y(n_15320)
);

AOI22xp5_ASAP7_75t_L g15321 ( 
.A1(n_15052),
.A2(n_2300),
.B1(n_2298),
.B2(n_2299),
.Y(n_15321)
);

AOI22xp33_ASAP7_75t_L g15322 ( 
.A1(n_15121),
.A2(n_2303),
.B1(n_2301),
.B2(n_2302),
.Y(n_15322)
);

INVx2_ASAP7_75t_L g15323 ( 
.A(n_15028),
.Y(n_15323)
);

AND2x6_ASAP7_75t_L g15324 ( 
.A(n_14939),
.B(n_15015),
.Y(n_15324)
);

AOI22xp5_ASAP7_75t_L g15325 ( 
.A1(n_14950),
.A2(n_2304),
.B1(n_2301),
.B2(n_2302),
.Y(n_15325)
);

OAI22xp5_ASAP7_75t_L g15326 ( 
.A1(n_15067),
.A2(n_2306),
.B1(n_2304),
.B2(n_2305),
.Y(n_15326)
);

NAND2xp5_ASAP7_75t_L g15327 ( 
.A(n_15056),
.B(n_2305),
.Y(n_15327)
);

INVx1_ASAP7_75t_L g15328 ( 
.A(n_15070),
.Y(n_15328)
);

AND2x2_ASAP7_75t_L g15329 ( 
.A(n_14934),
.B(n_2306),
.Y(n_15329)
);

INVx1_ASAP7_75t_L g15330 ( 
.A(n_14898),
.Y(n_15330)
);

BUFx6f_ASAP7_75t_L g15331 ( 
.A(n_15082),
.Y(n_15331)
);

OAI21xp5_ASAP7_75t_L g15332 ( 
.A1(n_15188),
.A2(n_2307),
.B(n_2308),
.Y(n_15332)
);

OAI221xp5_ASAP7_75t_L g15333 ( 
.A1(n_14989),
.A2(n_2309),
.B1(n_2307),
.B2(n_2308),
.C(n_2310),
.Y(n_15333)
);

AOI22xp33_ASAP7_75t_SL g15334 ( 
.A1(n_15233),
.A2(n_2312),
.B1(n_2309),
.B2(n_2311),
.Y(n_15334)
);

AOI22xp33_ASAP7_75t_L g15335 ( 
.A1(n_15054),
.A2(n_2313),
.B1(n_2311),
.B2(n_2312),
.Y(n_15335)
);

AND2x2_ASAP7_75t_L g15336 ( 
.A(n_14935),
.B(n_2313),
.Y(n_15336)
);

AND2x4_ASAP7_75t_L g15337 ( 
.A(n_14941),
.B(n_2314),
.Y(n_15337)
);

AND2x2_ASAP7_75t_L g15338 ( 
.A(n_14906),
.B(n_2315),
.Y(n_15338)
);

OAI22xp5_ASAP7_75t_L g15339 ( 
.A1(n_15225),
.A2(n_2319),
.B1(n_2316),
.B2(n_2317),
.Y(n_15339)
);

BUFx2_ASAP7_75t_L g15340 ( 
.A(n_15154),
.Y(n_15340)
);

INVx2_ASAP7_75t_L g15341 ( 
.A(n_15016),
.Y(n_15341)
);

OAI21x1_ASAP7_75t_L g15342 ( 
.A1(n_14978),
.A2(n_2317),
.B(n_2320),
.Y(n_15342)
);

AND2x2_ASAP7_75t_L g15343 ( 
.A(n_15055),
.B(n_2320),
.Y(n_15343)
);

CKINVDCx5p33_ASAP7_75t_R g15344 ( 
.A(n_14904),
.Y(n_15344)
);

NOR2xp33_ASAP7_75t_L g15345 ( 
.A(n_15250),
.B(n_2321),
.Y(n_15345)
);

AOI21xp5_ASAP7_75t_L g15346 ( 
.A1(n_14930),
.A2(n_14909),
.B(n_15102),
.Y(n_15346)
);

NAND2x1_ASAP7_75t_L g15347 ( 
.A(n_15085),
.B(n_2321),
.Y(n_15347)
);

AOI22xp33_ASAP7_75t_L g15348 ( 
.A1(n_14914),
.A2(n_2324),
.B1(n_2322),
.B2(n_2323),
.Y(n_15348)
);

OAI221xp5_ASAP7_75t_L g15349 ( 
.A1(n_15130),
.A2(n_2325),
.B1(n_2322),
.B2(n_2324),
.C(n_2326),
.Y(n_15349)
);

OAI22xp33_ASAP7_75t_L g15350 ( 
.A1(n_14893),
.A2(n_2327),
.B1(n_2325),
.B2(n_2326),
.Y(n_15350)
);

OAI211xp5_ASAP7_75t_L g15351 ( 
.A1(n_15135),
.A2(n_2329),
.B(n_2327),
.C(n_2328),
.Y(n_15351)
);

INVx1_ASAP7_75t_L g15352 ( 
.A(n_14902),
.Y(n_15352)
);

AOI22xp33_ASAP7_75t_L g15353 ( 
.A1(n_14912),
.A2(n_2330),
.B1(n_2328),
.B2(n_2329),
.Y(n_15353)
);

AOI22xp33_ASAP7_75t_L g15354 ( 
.A1(n_15108),
.A2(n_2332),
.B1(n_2330),
.B2(n_2331),
.Y(n_15354)
);

OAI22xp33_ASAP7_75t_L g15355 ( 
.A1(n_14931),
.A2(n_2334),
.B1(n_2332),
.B2(n_2333),
.Y(n_15355)
);

AOI22xp33_ASAP7_75t_L g15356 ( 
.A1(n_14937),
.A2(n_2336),
.B1(n_2333),
.B2(n_2335),
.Y(n_15356)
);

NAND2xp5_ASAP7_75t_L g15357 ( 
.A(n_15190),
.B(n_2336),
.Y(n_15357)
);

INVx1_ASAP7_75t_L g15358 ( 
.A(n_14903),
.Y(n_15358)
);

AOI222xp33_ASAP7_75t_L g15359 ( 
.A1(n_15165),
.A2(n_2339),
.B1(n_2341),
.B2(n_2337),
.C1(n_2338),
.C2(n_2340),
.Y(n_15359)
);

INVx1_ASAP7_75t_L g15360 ( 
.A(n_14905),
.Y(n_15360)
);

AND2x2_ASAP7_75t_L g15361 ( 
.A(n_15061),
.B(n_2337),
.Y(n_15361)
);

OR2x6_ASAP7_75t_L g15362 ( 
.A(n_15141),
.B(n_2338),
.Y(n_15362)
);

OAI21x1_ASAP7_75t_L g15363 ( 
.A1(n_15234),
.A2(n_2339),
.B(n_2340),
.Y(n_15363)
);

AOI22xp33_ASAP7_75t_L g15364 ( 
.A1(n_15003),
.A2(n_2343),
.B1(n_2341),
.B2(n_2342),
.Y(n_15364)
);

HB1xp67_ASAP7_75t_L g15365 ( 
.A(n_15035),
.Y(n_15365)
);

CKINVDCx5p33_ASAP7_75t_R g15366 ( 
.A(n_14913),
.Y(n_15366)
);

AOI22xp33_ASAP7_75t_L g15367 ( 
.A1(n_14936),
.A2(n_2345),
.B1(n_2342),
.B2(n_2344),
.Y(n_15367)
);

AOI22xp33_ASAP7_75t_L g15368 ( 
.A1(n_15059),
.A2(n_2346),
.B1(n_2344),
.B2(n_2345),
.Y(n_15368)
);

AOI22xp33_ASAP7_75t_L g15369 ( 
.A1(n_14957),
.A2(n_2348),
.B1(n_2346),
.B2(n_2347),
.Y(n_15369)
);

BUFx3_ASAP7_75t_L g15370 ( 
.A(n_15187),
.Y(n_15370)
);

AND2x2_ASAP7_75t_L g15371 ( 
.A(n_15118),
.B(n_2348),
.Y(n_15371)
);

OAI22xp5_ASAP7_75t_L g15372 ( 
.A1(n_15013),
.A2(n_2351),
.B1(n_2349),
.B2(n_2350),
.Y(n_15372)
);

AOI221xp5_ASAP7_75t_L g15373 ( 
.A1(n_15255),
.A2(n_2351),
.B1(n_2349),
.B2(n_2350),
.C(n_2352),
.Y(n_15373)
);

AOI22xp33_ASAP7_75t_L g15374 ( 
.A1(n_14917),
.A2(n_2354),
.B1(n_2352),
.B2(n_2353),
.Y(n_15374)
);

OR2x2_ASAP7_75t_L g15375 ( 
.A(n_15253),
.B(n_2353),
.Y(n_15375)
);

NAND2xp5_ASAP7_75t_L g15376 ( 
.A(n_15077),
.B(n_2354),
.Y(n_15376)
);

INVx1_ASAP7_75t_L g15377 ( 
.A(n_14919),
.Y(n_15377)
);

OAI22xp33_ASAP7_75t_L g15378 ( 
.A1(n_14931),
.A2(n_2357),
.B1(n_2355),
.B2(n_2356),
.Y(n_15378)
);

INVx1_ASAP7_75t_L g15379 ( 
.A(n_14920),
.Y(n_15379)
);

AND2x2_ASAP7_75t_L g15380 ( 
.A(n_14976),
.B(n_14984),
.Y(n_15380)
);

AOI222xp33_ASAP7_75t_L g15381 ( 
.A1(n_15165),
.A2(n_2357),
.B1(n_2359),
.B2(n_2355),
.C1(n_2356),
.C2(n_2358),
.Y(n_15381)
);

AOI221xp5_ASAP7_75t_L g15382 ( 
.A1(n_15185),
.A2(n_2361),
.B1(n_2358),
.B2(n_2359),
.C(n_2362),
.Y(n_15382)
);

AOI22xp33_ASAP7_75t_L g15383 ( 
.A1(n_15163),
.A2(n_2364),
.B1(n_2362),
.B2(n_2363),
.Y(n_15383)
);

AND2x2_ASAP7_75t_L g15384 ( 
.A(n_15092),
.B(n_2363),
.Y(n_15384)
);

AND2x2_ASAP7_75t_L g15385 ( 
.A(n_14979),
.B(n_2364),
.Y(n_15385)
);

INVx1_ASAP7_75t_L g15386 ( 
.A(n_14921),
.Y(n_15386)
);

AOI22xp33_ASAP7_75t_L g15387 ( 
.A1(n_15186),
.A2(n_2367),
.B1(n_2365),
.B2(n_2366),
.Y(n_15387)
);

OAI22xp5_ASAP7_75t_L g15388 ( 
.A1(n_15049),
.A2(n_2367),
.B1(n_2365),
.B2(n_2366),
.Y(n_15388)
);

A2O1A1Ixp33_ASAP7_75t_L g15389 ( 
.A1(n_15229),
.A2(n_2370),
.B(n_2368),
.C(n_2369),
.Y(n_15389)
);

NOR2xp33_ASAP7_75t_L g15390 ( 
.A(n_15018),
.B(n_2369),
.Y(n_15390)
);

AOI221xp5_ASAP7_75t_L g15391 ( 
.A1(n_15079),
.A2(n_2372),
.B1(n_2370),
.B2(n_2371),
.C(n_2373),
.Y(n_15391)
);

INVx1_ASAP7_75t_L g15392 ( 
.A(n_14924),
.Y(n_15392)
);

NOR2xp33_ASAP7_75t_L g15393 ( 
.A(n_15132),
.B(n_2372),
.Y(n_15393)
);

AOI22xp33_ASAP7_75t_SL g15394 ( 
.A1(n_15243),
.A2(n_2376),
.B1(n_2374),
.B2(n_2375),
.Y(n_15394)
);

INVx2_ASAP7_75t_L g15395 ( 
.A(n_15124),
.Y(n_15395)
);

AOI22xp33_ASAP7_75t_L g15396 ( 
.A1(n_15189),
.A2(n_2377),
.B1(n_2374),
.B2(n_2376),
.Y(n_15396)
);

INVx1_ASAP7_75t_L g15397 ( 
.A(n_14928),
.Y(n_15397)
);

INVx1_ASAP7_75t_L g15398 ( 
.A(n_14929),
.Y(n_15398)
);

AOI21xp33_ASAP7_75t_L g15399 ( 
.A1(n_15099),
.A2(n_2378),
.B(n_2379),
.Y(n_15399)
);

NOR2xp33_ASAP7_75t_L g15400 ( 
.A(n_15196),
.B(n_2378),
.Y(n_15400)
);

OAI21xp33_ASAP7_75t_L g15401 ( 
.A1(n_15087),
.A2(n_2379),
.B(n_2380),
.Y(n_15401)
);

AOI22xp33_ASAP7_75t_L g15402 ( 
.A1(n_15202),
.A2(n_2382),
.B1(n_2380),
.B2(n_2381),
.Y(n_15402)
);

BUFx2_ASAP7_75t_L g15403 ( 
.A(n_15169),
.Y(n_15403)
);

AND2x4_ASAP7_75t_L g15404 ( 
.A(n_15033),
.B(n_2381),
.Y(n_15404)
);

AOI22xp33_ASAP7_75t_L g15405 ( 
.A1(n_14970),
.A2(n_2384),
.B1(n_2382),
.B2(n_2383),
.Y(n_15405)
);

NAND2xp5_ASAP7_75t_L g15406 ( 
.A(n_15197),
.B(n_2383),
.Y(n_15406)
);

OAI22xp5_ASAP7_75t_SL g15407 ( 
.A1(n_14907),
.A2(n_2387),
.B1(n_2385),
.B2(n_2386),
.Y(n_15407)
);

NAND2xp5_ASAP7_75t_SL g15408 ( 
.A(n_15243),
.B(n_2385),
.Y(n_15408)
);

OAI21x1_ASAP7_75t_L g15409 ( 
.A1(n_15145),
.A2(n_2386),
.B(n_2387),
.Y(n_15409)
);

OAI22xp5_ASAP7_75t_L g15410 ( 
.A1(n_14951),
.A2(n_2390),
.B1(n_2388),
.B2(n_2389),
.Y(n_15410)
);

AOI21xp33_ASAP7_75t_L g15411 ( 
.A1(n_15064),
.A2(n_2388),
.B(n_2390),
.Y(n_15411)
);

AOI21x1_ASAP7_75t_L g15412 ( 
.A1(n_15191),
.A2(n_2391),
.B(n_2392),
.Y(n_15412)
);

AOI22xp33_ASAP7_75t_L g15413 ( 
.A1(n_15247),
.A2(n_2393),
.B1(n_2391),
.B2(n_2392),
.Y(n_15413)
);

AOI21xp33_ASAP7_75t_L g15414 ( 
.A1(n_15096),
.A2(n_2394),
.B(n_2395),
.Y(n_15414)
);

AOI221xp5_ASAP7_75t_L g15415 ( 
.A1(n_15224),
.A2(n_2398),
.B1(n_2396),
.B2(n_2397),
.C(n_2399),
.Y(n_15415)
);

NAND2xp5_ASAP7_75t_L g15416 ( 
.A(n_15194),
.B(n_2396),
.Y(n_15416)
);

AOI22xp33_ASAP7_75t_L g15417 ( 
.A1(n_14940),
.A2(n_2399),
.B1(n_2397),
.B2(n_2398),
.Y(n_15417)
);

HB1xp67_ASAP7_75t_L g15418 ( 
.A(n_15144),
.Y(n_15418)
);

INVx1_ASAP7_75t_L g15419 ( 
.A(n_14943),
.Y(n_15419)
);

OAI22xp33_ASAP7_75t_L g15420 ( 
.A1(n_15091),
.A2(n_2402),
.B1(n_2400),
.B2(n_2401),
.Y(n_15420)
);

INVx4_ASAP7_75t_SL g15421 ( 
.A(n_15025),
.Y(n_15421)
);

AOI21xp5_ASAP7_75t_L g15422 ( 
.A1(n_15238),
.A2(n_15074),
.B(n_15217),
.Y(n_15422)
);

INVxp67_ASAP7_75t_L g15423 ( 
.A(n_14977),
.Y(n_15423)
);

CKINVDCx20_ASAP7_75t_R g15424 ( 
.A(n_15126),
.Y(n_15424)
);

AOI221xp5_ASAP7_75t_L g15425 ( 
.A1(n_15227),
.A2(n_2403),
.B1(n_2401),
.B2(n_2402),
.C(n_2404),
.Y(n_15425)
);

AOI22xp33_ASAP7_75t_L g15426 ( 
.A1(n_15230),
.A2(n_15166),
.B1(n_15151),
.B2(n_15155),
.Y(n_15426)
);

OR2x2_ASAP7_75t_L g15427 ( 
.A(n_15097),
.B(n_2403),
.Y(n_15427)
);

OAI22xp5_ASAP7_75t_L g15428 ( 
.A1(n_14956),
.A2(n_2406),
.B1(n_2404),
.B2(n_2405),
.Y(n_15428)
);

NAND2xp5_ASAP7_75t_L g15429 ( 
.A(n_15170),
.B(n_2405),
.Y(n_15429)
);

AOI221xp5_ASAP7_75t_L g15430 ( 
.A1(n_15232),
.A2(n_2408),
.B1(n_2406),
.B2(n_2407),
.C(n_2409),
.Y(n_15430)
);

OR2x2_ASAP7_75t_L g15431 ( 
.A(n_15153),
.B(n_2407),
.Y(n_15431)
);

AOI22xp33_ASAP7_75t_SL g15432 ( 
.A1(n_14964),
.A2(n_2413),
.B1(n_2411),
.B2(n_2412),
.Y(n_15432)
);

BUFx3_ASAP7_75t_L g15433 ( 
.A(n_15142),
.Y(n_15433)
);

NAND2xp5_ASAP7_75t_L g15434 ( 
.A(n_15204),
.B(n_2411),
.Y(n_15434)
);

NAND2xp5_ASAP7_75t_L g15435 ( 
.A(n_15134),
.B(n_15005),
.Y(n_15435)
);

AOI22xp33_ASAP7_75t_L g15436 ( 
.A1(n_15156),
.A2(n_15081),
.B1(n_15103),
.B2(n_15179),
.Y(n_15436)
);

INVx2_ASAP7_75t_L g15437 ( 
.A(n_15010),
.Y(n_15437)
);

AOI21xp5_ASAP7_75t_L g15438 ( 
.A1(n_15218),
.A2(n_2412),
.B(n_2414),
.Y(n_15438)
);

INVx2_ASAP7_75t_L g15439 ( 
.A(n_15128),
.Y(n_15439)
);

AOI21xp5_ASAP7_75t_L g15440 ( 
.A1(n_15254),
.A2(n_2414),
.B(n_2415),
.Y(n_15440)
);

BUFx3_ASAP7_75t_L g15441 ( 
.A(n_15139),
.Y(n_15441)
);

OAI22xp33_ASAP7_75t_L g15442 ( 
.A1(n_15091),
.A2(n_2417),
.B1(n_2415),
.B2(n_2416),
.Y(n_15442)
);

NOR2xp33_ASAP7_75t_L g15443 ( 
.A(n_15228),
.B(n_2416),
.Y(n_15443)
);

INVx2_ASAP7_75t_L g15444 ( 
.A(n_15174),
.Y(n_15444)
);

OR2x2_ASAP7_75t_L g15445 ( 
.A(n_15026),
.B(n_2417),
.Y(n_15445)
);

AOI22xp33_ASAP7_75t_L g15446 ( 
.A1(n_15182),
.A2(n_2420),
.B1(n_2418),
.B2(n_2419),
.Y(n_15446)
);

AOI22xp33_ASAP7_75t_L g15447 ( 
.A1(n_15080),
.A2(n_2420),
.B1(n_2418),
.B2(n_2419),
.Y(n_15447)
);

AOI21xp5_ASAP7_75t_L g15448 ( 
.A1(n_15068),
.A2(n_15104),
.B(n_15252),
.Y(n_15448)
);

AOI22xp33_ASAP7_75t_L g15449 ( 
.A1(n_15216),
.A2(n_2423),
.B1(n_2421),
.B2(n_2422),
.Y(n_15449)
);

NAND2xp5_ASAP7_75t_L g15450 ( 
.A(n_15180),
.B(n_2421),
.Y(n_15450)
);

AOI22xp33_ASAP7_75t_L g15451 ( 
.A1(n_15205),
.A2(n_2424),
.B1(n_2422),
.B2(n_2423),
.Y(n_15451)
);

INVxp67_ASAP7_75t_SL g15452 ( 
.A(n_15089),
.Y(n_15452)
);

OAI33xp33_ASAP7_75t_L g15453 ( 
.A1(n_15071),
.A2(n_2426),
.A3(n_2428),
.B1(n_2424),
.B2(n_2425),
.B3(n_2427),
.Y(n_15453)
);

INVx1_ASAP7_75t_L g15454 ( 
.A(n_14944),
.Y(n_15454)
);

NAND2xp5_ASAP7_75t_L g15455 ( 
.A(n_15210),
.B(n_15214),
.Y(n_15455)
);

INVx2_ASAP7_75t_L g15456 ( 
.A(n_15240),
.Y(n_15456)
);

AOI221x1_ASAP7_75t_SL g15457 ( 
.A1(n_15072),
.A2(n_2428),
.B1(n_2425),
.B2(n_2427),
.C(n_2429),
.Y(n_15457)
);

AOI21xp5_ASAP7_75t_L g15458 ( 
.A1(n_15065),
.A2(n_2429),
.B(n_2430),
.Y(n_15458)
);

OAI211xp5_ASAP7_75t_L g15459 ( 
.A1(n_15034),
.A2(n_15107),
.B(n_15245),
.C(n_15083),
.Y(n_15459)
);

AOI22xp33_ASAP7_75t_L g15460 ( 
.A1(n_14960),
.A2(n_2432),
.B1(n_2430),
.B2(n_2431),
.Y(n_15460)
);

AOI22xp33_ASAP7_75t_L g15461 ( 
.A1(n_14961),
.A2(n_2434),
.B1(n_2431),
.B2(n_2433),
.Y(n_15461)
);

OAI22xp5_ASAP7_75t_L g15462 ( 
.A1(n_14969),
.A2(n_15001),
.B1(n_15027),
.B2(n_15222),
.Y(n_15462)
);

NOR2xp33_ASAP7_75t_L g15463 ( 
.A(n_14954),
.B(n_15212),
.Y(n_15463)
);

OA21x2_ASAP7_75t_L g15464 ( 
.A1(n_15039),
.A2(n_2433),
.B(n_2434),
.Y(n_15464)
);

INVx3_ASAP7_75t_L g15465 ( 
.A(n_15017),
.Y(n_15465)
);

BUFx4f_ASAP7_75t_SL g15466 ( 
.A(n_15022),
.Y(n_15466)
);

AOI22xp33_ASAP7_75t_SL g15467 ( 
.A1(n_15246),
.A2(n_2437),
.B1(n_2435),
.B2(n_2436),
.Y(n_15467)
);

AOI21xp5_ASAP7_75t_L g15468 ( 
.A1(n_15215),
.A2(n_2436),
.B(n_2437),
.Y(n_15468)
);

AOI22xp33_ASAP7_75t_L g15469 ( 
.A1(n_15086),
.A2(n_2441),
.B1(n_2438),
.B2(n_2439),
.Y(n_15469)
);

OAI221xp5_ASAP7_75t_L g15470 ( 
.A1(n_15090),
.A2(n_2441),
.B1(n_2438),
.B2(n_2439),
.C(n_2442),
.Y(n_15470)
);

OAI22xp33_ASAP7_75t_L g15471 ( 
.A1(n_15211),
.A2(n_2444),
.B1(n_2442),
.B2(n_2443),
.Y(n_15471)
);

AND2x2_ASAP7_75t_L g15472 ( 
.A(n_15008),
.B(n_2443),
.Y(n_15472)
);

OAI221xp5_ASAP7_75t_L g15473 ( 
.A1(n_15006),
.A2(n_2447),
.B1(n_2445),
.B2(n_2446),
.C(n_2448),
.Y(n_15473)
);

BUFx2_ASAP7_75t_L g15474 ( 
.A(n_14958),
.Y(n_15474)
);

OAI221xp5_ASAP7_75t_L g15475 ( 
.A1(n_15011),
.A2(n_2448),
.B1(n_2445),
.B2(n_2447),
.C(n_2449),
.Y(n_15475)
);

OAI22xp5_ASAP7_75t_L g15476 ( 
.A1(n_15012),
.A2(n_15136),
.B1(n_15063),
.B2(n_15073),
.Y(n_15476)
);

INVx1_ASAP7_75t_L g15477 ( 
.A(n_14945),
.Y(n_15477)
);

AND2x4_ASAP7_75t_L g15478 ( 
.A(n_15060),
.B(n_2449),
.Y(n_15478)
);

OAI22xp5_ASAP7_75t_L g15479 ( 
.A1(n_15140),
.A2(n_2452),
.B1(n_2450),
.B2(n_2451),
.Y(n_15479)
);

OR2x2_ASAP7_75t_L g15480 ( 
.A(n_15112),
.B(n_2450),
.Y(n_15480)
);

HB1xp67_ASAP7_75t_L g15481 ( 
.A(n_15149),
.Y(n_15481)
);

AOI22xp33_ASAP7_75t_L g15482 ( 
.A1(n_15051),
.A2(n_2453),
.B1(n_2451),
.B2(n_2452),
.Y(n_15482)
);

INVxp67_ASAP7_75t_L g15483 ( 
.A(n_15031),
.Y(n_15483)
);

AOI22xp33_ASAP7_75t_L g15484 ( 
.A1(n_15157),
.A2(n_2455),
.B1(n_2453),
.B2(n_2454),
.Y(n_15484)
);

AOI22xp33_ASAP7_75t_L g15485 ( 
.A1(n_14968),
.A2(n_2457),
.B1(n_2455),
.B2(n_2456),
.Y(n_15485)
);

AND2x2_ASAP7_75t_L g15486 ( 
.A(n_15098),
.B(n_15168),
.Y(n_15486)
);

INVx1_ASAP7_75t_L g15487 ( 
.A(n_14946),
.Y(n_15487)
);

AOI22xp33_ASAP7_75t_L g15488 ( 
.A1(n_15019),
.A2(n_2458),
.B1(n_2456),
.B2(n_2457),
.Y(n_15488)
);

AO21x2_ASAP7_75t_L g15489 ( 
.A1(n_15041),
.A2(n_2458),
.B(n_2459),
.Y(n_15489)
);

OR2x2_ASAP7_75t_L g15490 ( 
.A(n_15201),
.B(n_2459),
.Y(n_15490)
);

AND2x2_ASAP7_75t_SL g15491 ( 
.A(n_14985),
.B(n_2461),
.Y(n_15491)
);

AOI22xp33_ASAP7_75t_L g15492 ( 
.A1(n_15235),
.A2(n_2463),
.B1(n_2461),
.B2(n_2462),
.Y(n_15492)
);

AND2x2_ASAP7_75t_L g15493 ( 
.A(n_15088),
.B(n_15076),
.Y(n_15493)
);

INVxp67_ASAP7_75t_SL g15494 ( 
.A(n_15046),
.Y(n_15494)
);

AND2x4_ASAP7_75t_L g15495 ( 
.A(n_14982),
.B(n_2462),
.Y(n_15495)
);

OAI22x1_ASAP7_75t_L g15496 ( 
.A1(n_15158),
.A2(n_15164),
.B1(n_14988),
.B2(n_15119),
.Y(n_15496)
);

AOI22xp33_ASAP7_75t_L g15497 ( 
.A1(n_15176),
.A2(n_15221),
.B1(n_15133),
.B2(n_15042),
.Y(n_15497)
);

OR2x6_ASAP7_75t_L g15498 ( 
.A(n_15195),
.B(n_2463),
.Y(n_15498)
);

AOI222xp33_ASAP7_75t_L g15499 ( 
.A1(n_15093),
.A2(n_2466),
.B1(n_2468),
.B2(n_2464),
.C1(n_2465),
.C2(n_2467),
.Y(n_15499)
);

NAND2x1_ASAP7_75t_L g15500 ( 
.A(n_15147),
.B(n_2464),
.Y(n_15500)
);

AND2x2_ASAP7_75t_L g15501 ( 
.A(n_15171),
.B(n_2465),
.Y(n_15501)
);

OAI22xp33_ASAP7_75t_L g15502 ( 
.A1(n_15115),
.A2(n_2469),
.B1(n_2466),
.B2(n_2468),
.Y(n_15502)
);

INVx1_ASAP7_75t_L g15503 ( 
.A(n_14947),
.Y(n_15503)
);

NOR4xp25_ASAP7_75t_L g15504 ( 
.A(n_15105),
.B(n_2471),
.C(n_2469),
.D(n_2470),
.Y(n_15504)
);

AND2x2_ASAP7_75t_L g15505 ( 
.A(n_15009),
.B(n_2470),
.Y(n_15505)
);

AOI21xp5_ASAP7_75t_L g15506 ( 
.A1(n_15106),
.A2(n_15177),
.B(n_15113),
.Y(n_15506)
);

AOI22xp5_ASAP7_75t_L g15507 ( 
.A1(n_15078),
.A2(n_2473),
.B1(n_2471),
.B2(n_2472),
.Y(n_15507)
);

AOI22xp33_ASAP7_75t_L g15508 ( 
.A1(n_15101),
.A2(n_2476),
.B1(n_2472),
.B2(n_2474),
.Y(n_15508)
);

OAI211xp5_ASAP7_75t_L g15509 ( 
.A1(n_15160),
.A2(n_2477),
.B(n_2474),
.C(n_2476),
.Y(n_15509)
);

O2A1O1Ixp33_ASAP7_75t_L g15510 ( 
.A1(n_15122),
.A2(n_2480),
.B(n_2478),
.C(n_2479),
.Y(n_15510)
);

NAND2xp5_ASAP7_75t_L g15511 ( 
.A(n_15116),
.B(n_2478),
.Y(n_15511)
);

OAI21xp5_ASAP7_75t_L g15512 ( 
.A1(n_14974),
.A2(n_2479),
.B(n_2480),
.Y(n_15512)
);

AOI22xp33_ASAP7_75t_L g15513 ( 
.A1(n_15175),
.A2(n_2483),
.B1(n_2481),
.B2(n_2482),
.Y(n_15513)
);

AOI22xp33_ASAP7_75t_L g15514 ( 
.A1(n_15161),
.A2(n_2483),
.B1(n_2481),
.B2(n_2482),
.Y(n_15514)
);

OAI22xp5_ASAP7_75t_L g15515 ( 
.A1(n_15159),
.A2(n_2486),
.B1(n_2484),
.B2(n_2485),
.Y(n_15515)
);

AOI221xp5_ASAP7_75t_SL g15516 ( 
.A1(n_15084),
.A2(n_2486),
.B1(n_2484),
.B2(n_2485),
.C(n_2487),
.Y(n_15516)
);

AOI22xp33_ASAP7_75t_SL g15517 ( 
.A1(n_15162),
.A2(n_2489),
.B1(n_2487),
.B2(n_2488),
.Y(n_15517)
);

AOI221xp5_ASAP7_75t_SL g15518 ( 
.A1(n_15094),
.A2(n_15114),
.B1(n_15150),
.B2(n_15146),
.C(n_15100),
.Y(n_15518)
);

NAND2xp5_ASAP7_75t_L g15519 ( 
.A(n_15095),
.B(n_2488),
.Y(n_15519)
);

HB1xp67_ASAP7_75t_L g15520 ( 
.A(n_15184),
.Y(n_15520)
);

AND2x2_ASAP7_75t_L g15521 ( 
.A(n_15219),
.B(n_2490),
.Y(n_15521)
);

HB1xp67_ASAP7_75t_L g15522 ( 
.A(n_15365),
.Y(n_15522)
);

INVx2_ASAP7_75t_L g15523 ( 
.A(n_15318),
.Y(n_15523)
);

INVx2_ASAP7_75t_L g15524 ( 
.A(n_15318),
.Y(n_15524)
);

AND2x2_ASAP7_75t_L g15525 ( 
.A(n_15340),
.B(n_15129),
.Y(n_15525)
);

INVx1_ASAP7_75t_L g15526 ( 
.A(n_15276),
.Y(n_15526)
);

BUFx3_ASAP7_75t_L g15527 ( 
.A(n_15260),
.Y(n_15527)
);

AND2x2_ASAP7_75t_L g15528 ( 
.A(n_15266),
.B(n_15075),
.Y(n_15528)
);

INVx1_ASAP7_75t_L g15529 ( 
.A(n_15418),
.Y(n_15529)
);

NAND2xp5_ASAP7_75t_L g15530 ( 
.A(n_15452),
.B(n_15242),
.Y(n_15530)
);

AND2x2_ASAP7_75t_L g15531 ( 
.A(n_15313),
.B(n_15062),
.Y(n_15531)
);

NAND2xp5_ASAP7_75t_L g15532 ( 
.A(n_15264),
.B(n_15249),
.Y(n_15532)
);

AND2x2_ASAP7_75t_L g15533 ( 
.A(n_15403),
.B(n_15109),
.Y(n_15533)
);

HB1xp67_ASAP7_75t_L g15534 ( 
.A(n_15284),
.Y(n_15534)
);

INVx1_ASAP7_75t_L g15535 ( 
.A(n_15299),
.Y(n_15535)
);

INVx4_ASAP7_75t_L g15536 ( 
.A(n_15287),
.Y(n_15536)
);

NAND2xp5_ASAP7_75t_L g15537 ( 
.A(n_15474),
.B(n_14992),
.Y(n_15537)
);

NAND2xp5_ASAP7_75t_L g15538 ( 
.A(n_15283),
.B(n_14997),
.Y(n_15538)
);

AND2x2_ASAP7_75t_L g15539 ( 
.A(n_15265),
.B(n_15110),
.Y(n_15539)
);

CKINVDCx6p67_ASAP7_75t_R g15540 ( 
.A(n_15324),
.Y(n_15540)
);

INVx1_ASAP7_75t_L g15541 ( 
.A(n_15274),
.Y(n_15541)
);

NAND2xp5_ASAP7_75t_L g15542 ( 
.A(n_15267),
.B(n_15002),
.Y(n_15542)
);

NAND2xp5_ASAP7_75t_L g15543 ( 
.A(n_15483),
.B(n_15167),
.Y(n_15543)
);

OR2x2_ASAP7_75t_L g15544 ( 
.A(n_15256),
.B(n_15043),
.Y(n_15544)
);

AND2x2_ASAP7_75t_L g15545 ( 
.A(n_15370),
.B(n_15125),
.Y(n_15545)
);

AOI22xp33_ASAP7_75t_L g15546 ( 
.A1(n_15268),
.A2(n_14994),
.B1(n_15172),
.B2(n_15143),
.Y(n_15546)
);

OR2x2_ASAP7_75t_L g15547 ( 
.A(n_15294),
.B(n_15044),
.Y(n_15547)
);

AND2x2_ASAP7_75t_L g15548 ( 
.A(n_15288),
.B(n_15045),
.Y(n_15548)
);

INVx2_ASAP7_75t_L g15549 ( 
.A(n_15331),
.Y(n_15549)
);

INVx1_ASAP7_75t_L g15550 ( 
.A(n_15262),
.Y(n_15550)
);

INVx2_ASAP7_75t_L g15551 ( 
.A(n_15331),
.Y(n_15551)
);

BUFx2_ASAP7_75t_L g15552 ( 
.A(n_15324),
.Y(n_15552)
);

INVx2_ASAP7_75t_L g15553 ( 
.A(n_15466),
.Y(n_15553)
);

AND2x2_ASAP7_75t_L g15554 ( 
.A(n_15308),
.B(n_15047),
.Y(n_15554)
);

INVx2_ASAP7_75t_L g15555 ( 
.A(n_15296),
.Y(n_15555)
);

AND2x2_ASAP7_75t_L g15556 ( 
.A(n_15280),
.B(n_15048),
.Y(n_15556)
);

INVxp67_ASAP7_75t_L g15557 ( 
.A(n_15324),
.Y(n_15557)
);

INVx1_ASAP7_75t_L g15558 ( 
.A(n_15314),
.Y(n_15558)
);

NOR2x1_ASAP7_75t_L g15559 ( 
.A(n_15500),
.B(n_15038),
.Y(n_15559)
);

OR2x2_ASAP7_75t_L g15560 ( 
.A(n_15290),
.B(n_14991),
.Y(n_15560)
);

INVx2_ASAP7_75t_L g15561 ( 
.A(n_15424),
.Y(n_15561)
);

AND2x2_ASAP7_75t_L g15562 ( 
.A(n_15323),
.B(n_15207),
.Y(n_15562)
);

HB1xp67_ASAP7_75t_L g15563 ( 
.A(n_15284),
.Y(n_15563)
);

INVx1_ASAP7_75t_L g15564 ( 
.A(n_15375),
.Y(n_15564)
);

BUFx2_ASAP7_75t_L g15565 ( 
.A(n_15423),
.Y(n_15565)
);

INVx2_ASAP7_75t_L g15566 ( 
.A(n_15433),
.Y(n_15566)
);

NAND2xp5_ASAP7_75t_L g15567 ( 
.A(n_15302),
.B(n_14948),
.Y(n_15567)
);

AND2x2_ASAP7_75t_L g15568 ( 
.A(n_15258),
.B(n_15173),
.Y(n_15568)
);

INVx1_ASAP7_75t_L g15569 ( 
.A(n_15285),
.Y(n_15569)
);

OAI22xp5_ASAP7_75t_L g15570 ( 
.A1(n_15257),
.A2(n_14990),
.B1(n_14980),
.B2(n_14998),
.Y(n_15570)
);

INVx2_ASAP7_75t_L g15571 ( 
.A(n_15441),
.Y(n_15571)
);

BUFx6f_ASAP7_75t_L g15572 ( 
.A(n_15404),
.Y(n_15572)
);

BUFx2_ASAP7_75t_L g15573 ( 
.A(n_15362),
.Y(n_15573)
);

INVx2_ASAP7_75t_L g15574 ( 
.A(n_15278),
.Y(n_15574)
);

HB1xp67_ASAP7_75t_L g15575 ( 
.A(n_15421),
.Y(n_15575)
);

AND2x2_ASAP7_75t_L g15576 ( 
.A(n_15270),
.B(n_15208),
.Y(n_15576)
);

NAND2xp5_ASAP7_75t_L g15577 ( 
.A(n_15432),
.B(n_14949),
.Y(n_15577)
);

INVx1_ASAP7_75t_L g15578 ( 
.A(n_15292),
.Y(n_15578)
);

INVx5_ASAP7_75t_SL g15579 ( 
.A(n_15362),
.Y(n_15579)
);

INVxp67_ASAP7_75t_SL g15580 ( 
.A(n_15347),
.Y(n_15580)
);

INVx2_ASAP7_75t_L g15581 ( 
.A(n_15395),
.Y(n_15581)
);

AND2x2_ASAP7_75t_L g15582 ( 
.A(n_15279),
.B(n_15251),
.Y(n_15582)
);

INVxp67_ASAP7_75t_L g15583 ( 
.A(n_15481),
.Y(n_15583)
);

HB1xp67_ASAP7_75t_L g15584 ( 
.A(n_15421),
.Y(n_15584)
);

NAND2xp5_ASAP7_75t_L g15585 ( 
.A(n_15504),
.B(n_14952),
.Y(n_15585)
);

INVx2_ASAP7_75t_L g15586 ( 
.A(n_15465),
.Y(n_15586)
);

BUFx3_ASAP7_75t_L g15587 ( 
.A(n_15344),
.Y(n_15587)
);

INVx2_ASAP7_75t_L g15588 ( 
.A(n_15341),
.Y(n_15588)
);

AND2x4_ASAP7_75t_SL g15589 ( 
.A(n_15281),
.B(n_15337),
.Y(n_15589)
);

INVx2_ASAP7_75t_L g15590 ( 
.A(n_15439),
.Y(n_15590)
);

NAND2xp5_ASAP7_75t_L g15591 ( 
.A(n_15346),
.B(n_14959),
.Y(n_15591)
);

HB1xp67_ASAP7_75t_L g15592 ( 
.A(n_15464),
.Y(n_15592)
);

INVx1_ASAP7_75t_L g15593 ( 
.A(n_15328),
.Y(n_15593)
);

AND2x2_ASAP7_75t_L g15594 ( 
.A(n_15493),
.B(n_14999),
.Y(n_15594)
);

INVx1_ASAP7_75t_L g15595 ( 
.A(n_15445),
.Y(n_15595)
);

BUFx3_ASAP7_75t_L g15596 ( 
.A(n_15478),
.Y(n_15596)
);

INVx3_ASAP7_75t_L g15597 ( 
.A(n_15444),
.Y(n_15597)
);

INVx2_ASAP7_75t_L g15598 ( 
.A(n_15437),
.Y(n_15598)
);

HB1xp67_ASAP7_75t_L g15599 ( 
.A(n_15464),
.Y(n_15599)
);

OR2x2_ASAP7_75t_L g15600 ( 
.A(n_15269),
.B(n_15000),
.Y(n_15600)
);

INVx2_ASAP7_75t_L g15601 ( 
.A(n_15456),
.Y(n_15601)
);

HB1xp67_ASAP7_75t_L g15602 ( 
.A(n_15520),
.Y(n_15602)
);

AND2x2_ASAP7_75t_L g15603 ( 
.A(n_15486),
.B(n_15020),
.Y(n_15603)
);

INVx2_ASAP7_75t_L g15604 ( 
.A(n_15380),
.Y(n_15604)
);

BUFx3_ASAP7_75t_L g15605 ( 
.A(n_15498),
.Y(n_15605)
);

AND2x2_ASAP7_75t_L g15606 ( 
.A(n_15494),
.B(n_15029),
.Y(n_15606)
);

AND2x2_ASAP7_75t_L g15607 ( 
.A(n_15463),
.B(n_15032),
.Y(n_15607)
);

OR2x2_ASAP7_75t_L g15608 ( 
.A(n_15435),
.B(n_14966),
.Y(n_15608)
);

NAND2xp5_ASAP7_75t_L g15609 ( 
.A(n_15277),
.B(n_14972),
.Y(n_15609)
);

INVx3_ASAP7_75t_L g15610 ( 
.A(n_15366),
.Y(n_15610)
);

INVx1_ASAP7_75t_L g15611 ( 
.A(n_15310),
.Y(n_15611)
);

INVx2_ASAP7_75t_L g15612 ( 
.A(n_15343),
.Y(n_15612)
);

INVx3_ASAP7_75t_SL g15613 ( 
.A(n_15498),
.Y(n_15613)
);

INVx2_ASAP7_75t_L g15614 ( 
.A(n_15289),
.Y(n_15614)
);

AND2x2_ASAP7_75t_L g15615 ( 
.A(n_15304),
.B(n_15069),
.Y(n_15615)
);

INVx2_ASAP7_75t_L g15616 ( 
.A(n_15338),
.Y(n_15616)
);

INVx2_ASAP7_75t_L g15617 ( 
.A(n_15329),
.Y(n_15617)
);

AND2x2_ASAP7_75t_L g15618 ( 
.A(n_15491),
.B(n_14975),
.Y(n_15618)
);

INVx1_ASAP7_75t_L g15619 ( 
.A(n_15330),
.Y(n_15619)
);

INVxp67_ASAP7_75t_L g15620 ( 
.A(n_15315),
.Y(n_15620)
);

HB1xp67_ASAP7_75t_L g15621 ( 
.A(n_15489),
.Y(n_15621)
);

AND2x2_ASAP7_75t_L g15622 ( 
.A(n_15309),
.B(n_15030),
.Y(n_15622)
);

INVx2_ASAP7_75t_L g15623 ( 
.A(n_15336),
.Y(n_15623)
);

INVx1_ASAP7_75t_L g15624 ( 
.A(n_15352),
.Y(n_15624)
);

NOR2x1_ASAP7_75t_L g15625 ( 
.A(n_15291),
.B(n_15248),
.Y(n_15625)
);

INVx1_ASAP7_75t_L g15626 ( 
.A(n_15358),
.Y(n_15626)
);

OR2x2_ASAP7_75t_L g15627 ( 
.A(n_15455),
.B(n_15178),
.Y(n_15627)
);

INVx1_ASAP7_75t_L g15628 ( 
.A(n_15360),
.Y(n_15628)
);

AND2x2_ASAP7_75t_L g15629 ( 
.A(n_15501),
.B(n_14955),
.Y(n_15629)
);

INVx1_ASAP7_75t_L g15630 ( 
.A(n_15377),
.Y(n_15630)
);

INVxp67_ASAP7_75t_SL g15631 ( 
.A(n_15408),
.Y(n_15631)
);

AND2x4_ASAP7_75t_L g15632 ( 
.A(n_15361),
.B(n_14987),
.Y(n_15632)
);

INVx2_ASAP7_75t_L g15633 ( 
.A(n_15385),
.Y(n_15633)
);

NAND2x1p5_ASAP7_75t_L g15634 ( 
.A(n_15312),
.B(n_15014),
.Y(n_15634)
);

INVx3_ASAP7_75t_L g15635 ( 
.A(n_15495),
.Y(n_15635)
);

BUFx6f_ASAP7_75t_L g15636 ( 
.A(n_15384),
.Y(n_15636)
);

INVx1_ASAP7_75t_L g15637 ( 
.A(n_15379),
.Y(n_15637)
);

AND2x2_ASAP7_75t_L g15638 ( 
.A(n_15462),
.B(n_14986),
.Y(n_15638)
);

NAND2xp5_ASAP7_75t_L g15639 ( 
.A(n_15422),
.B(n_15025),
.Y(n_15639)
);

AND2x2_ASAP7_75t_L g15640 ( 
.A(n_15521),
.B(n_2490),
.Y(n_15640)
);

NAND2xp5_ASAP7_75t_L g15641 ( 
.A(n_15259),
.B(n_2491),
.Y(n_15641)
);

INVx2_ASAP7_75t_L g15642 ( 
.A(n_15371),
.Y(n_15642)
);

INVx2_ASAP7_75t_L g15643 ( 
.A(n_15319),
.Y(n_15643)
);

AND2x2_ASAP7_75t_L g15644 ( 
.A(n_15426),
.B(n_2491),
.Y(n_15644)
);

INVx1_ASAP7_75t_L g15645 ( 
.A(n_15386),
.Y(n_15645)
);

INVx1_ASAP7_75t_L g15646 ( 
.A(n_15392),
.Y(n_15646)
);

NAND4xp25_ASAP7_75t_L g15647 ( 
.A(n_15436),
.B(n_2494),
.C(n_2492),
.D(n_2493),
.Y(n_15647)
);

NAND2xp5_ASAP7_75t_L g15648 ( 
.A(n_15293),
.B(n_2492),
.Y(n_15648)
);

HB1xp67_ASAP7_75t_L g15649 ( 
.A(n_15496),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_15397),
.Y(n_15650)
);

INVx2_ASAP7_75t_R g15651 ( 
.A(n_15398),
.Y(n_15651)
);

NOR2xp33_ASAP7_75t_L g15652 ( 
.A(n_15271),
.B(n_2493),
.Y(n_15652)
);

OR2x2_ASAP7_75t_L g15653 ( 
.A(n_15476),
.B(n_2494),
.Y(n_15653)
);

AND2x2_ASAP7_75t_L g15654 ( 
.A(n_15472),
.B(n_2495),
.Y(n_15654)
);

AND2x4_ASAP7_75t_L g15655 ( 
.A(n_15327),
.B(n_2495),
.Y(n_15655)
);

INVx2_ASAP7_75t_L g15656 ( 
.A(n_15409),
.Y(n_15656)
);

INVx2_ASAP7_75t_L g15657 ( 
.A(n_15480),
.Y(n_15657)
);

INVx1_ASAP7_75t_L g15658 ( 
.A(n_15419),
.Y(n_15658)
);

INVx1_ASAP7_75t_L g15659 ( 
.A(n_15454),
.Y(n_15659)
);

INVx2_ASAP7_75t_L g15660 ( 
.A(n_15427),
.Y(n_15660)
);

NAND2xp5_ASAP7_75t_L g15661 ( 
.A(n_15438),
.B(n_2496),
.Y(n_15661)
);

BUFx6f_ASAP7_75t_L g15662 ( 
.A(n_15357),
.Y(n_15662)
);

INVx1_ASAP7_75t_L g15663 ( 
.A(n_15477),
.Y(n_15663)
);

AOI22xp33_ASAP7_75t_L g15664 ( 
.A1(n_15263),
.A2(n_2499),
.B1(n_2497),
.B2(n_2498),
.Y(n_15664)
);

INVx1_ASAP7_75t_L g15665 ( 
.A(n_15487),
.Y(n_15665)
);

INVx2_ASAP7_75t_SL g15666 ( 
.A(n_15505),
.Y(n_15666)
);

INVx1_ASAP7_75t_L g15667 ( 
.A(n_15503),
.Y(n_15667)
);

NAND2xp5_ASAP7_75t_L g15668 ( 
.A(n_15440),
.B(n_15468),
.Y(n_15668)
);

INVx3_ASAP7_75t_L g15669 ( 
.A(n_15490),
.Y(n_15669)
);

INVxp67_ASAP7_75t_R g15670 ( 
.A(n_15407),
.Y(n_15670)
);

INVx2_ASAP7_75t_L g15671 ( 
.A(n_15363),
.Y(n_15671)
);

OR2x2_ASAP7_75t_L g15672 ( 
.A(n_15286),
.B(n_2498),
.Y(n_15672)
);

AND2x2_ASAP7_75t_L g15673 ( 
.A(n_15345),
.B(n_2500),
.Y(n_15673)
);

INVxp67_ASAP7_75t_SL g15674 ( 
.A(n_15400),
.Y(n_15674)
);

INVx3_ASAP7_75t_L g15675 ( 
.A(n_15431),
.Y(n_15675)
);

AND2x2_ASAP7_75t_L g15676 ( 
.A(n_15390),
.B(n_2500),
.Y(n_15676)
);

INVx2_ASAP7_75t_L g15677 ( 
.A(n_15342),
.Y(n_15677)
);

INVx1_ASAP7_75t_L g15678 ( 
.A(n_15416),
.Y(n_15678)
);

NAND2xp5_ASAP7_75t_L g15679 ( 
.A(n_15401),
.B(n_2501),
.Y(n_15679)
);

INVx2_ASAP7_75t_L g15680 ( 
.A(n_15412),
.Y(n_15680)
);

INVx1_ASAP7_75t_L g15681 ( 
.A(n_15406),
.Y(n_15681)
);

INVx1_ASAP7_75t_L g15682 ( 
.A(n_15434),
.Y(n_15682)
);

AND2x2_ASAP7_75t_L g15683 ( 
.A(n_15393),
.B(n_2502),
.Y(n_15683)
);

AND2x2_ASAP7_75t_L g15684 ( 
.A(n_15429),
.B(n_2502),
.Y(n_15684)
);

INVx1_ASAP7_75t_SL g15685 ( 
.A(n_15511),
.Y(n_15685)
);

AND2x2_ASAP7_75t_L g15686 ( 
.A(n_15443),
.B(n_2503),
.Y(n_15686)
);

NAND2xp5_ASAP7_75t_L g15687 ( 
.A(n_15355),
.B(n_2503),
.Y(n_15687)
);

NAND2xp5_ASAP7_75t_L g15688 ( 
.A(n_15378),
.B(n_2504),
.Y(n_15688)
);

INVx4_ASAP7_75t_L g15689 ( 
.A(n_15519),
.Y(n_15689)
);

AOI22xp33_ASAP7_75t_L g15690 ( 
.A1(n_15261),
.A2(n_2507),
.B1(n_2505),
.B2(n_2506),
.Y(n_15690)
);

INVx2_ASAP7_75t_L g15691 ( 
.A(n_15450),
.Y(n_15691)
);

AND2x2_ASAP7_75t_L g15692 ( 
.A(n_15497),
.B(n_2505),
.Y(n_15692)
);

INVx2_ASAP7_75t_L g15693 ( 
.A(n_15376),
.Y(n_15693)
);

AND2x2_ASAP7_75t_L g15694 ( 
.A(n_15307),
.B(n_2506),
.Y(n_15694)
);

INVx1_ASAP7_75t_L g15695 ( 
.A(n_15515),
.Y(n_15695)
);

INVx1_ASAP7_75t_L g15696 ( 
.A(n_15297),
.Y(n_15696)
);

INVx1_ASAP7_75t_L g15697 ( 
.A(n_15506),
.Y(n_15697)
);

INVx1_ASAP7_75t_L g15698 ( 
.A(n_15306),
.Y(n_15698)
);

NOR2xp33_ASAP7_75t_L g15699 ( 
.A(n_15303),
.B(n_2507),
.Y(n_15699)
);

INVx5_ASAP7_75t_L g15700 ( 
.A(n_15359),
.Y(n_15700)
);

INVx2_ASAP7_75t_L g15701 ( 
.A(n_15388),
.Y(n_15701)
);

AND2x2_ASAP7_75t_L g15702 ( 
.A(n_15272),
.B(n_2508),
.Y(n_15702)
);

INVx1_ASAP7_75t_L g15703 ( 
.A(n_15326),
.Y(n_15703)
);

INVx1_ASAP7_75t_L g15704 ( 
.A(n_15350),
.Y(n_15704)
);

INVx2_ASAP7_75t_L g15705 ( 
.A(n_15298),
.Y(n_15705)
);

AND2x4_ASAP7_75t_L g15706 ( 
.A(n_15332),
.B(n_2508),
.Y(n_15706)
);

AND2x2_ASAP7_75t_L g15707 ( 
.A(n_15273),
.B(n_2509),
.Y(n_15707)
);

INVx2_ASAP7_75t_L g15708 ( 
.A(n_15321),
.Y(n_15708)
);

INVxp67_ASAP7_75t_R g15709 ( 
.A(n_15372),
.Y(n_15709)
);

INVx1_ASAP7_75t_L g15710 ( 
.A(n_15300),
.Y(n_15710)
);

INVx1_ASAP7_75t_L g15711 ( 
.A(n_15459),
.Y(n_15711)
);

INVx3_ASAP7_75t_SL g15712 ( 
.A(n_15394),
.Y(n_15712)
);

BUFx2_ASAP7_75t_SL g15713 ( 
.A(n_15458),
.Y(n_15713)
);

BUFx2_ASAP7_75t_L g15714 ( 
.A(n_15512),
.Y(n_15714)
);

AND2x2_ASAP7_75t_L g15715 ( 
.A(n_15448),
.B(n_2510),
.Y(n_15715)
);

AND2x2_ASAP7_75t_L g15716 ( 
.A(n_15518),
.B(n_2510),
.Y(n_15716)
);

NAND2xp5_ASAP7_75t_L g15717 ( 
.A(n_15275),
.B(n_2511),
.Y(n_15717)
);

OR2x2_ASAP7_75t_L g15718 ( 
.A(n_15320),
.B(n_2511),
.Y(n_15718)
);

AND2x2_ASAP7_75t_L g15719 ( 
.A(n_15311),
.B(n_2512),
.Y(n_15719)
);

INVx2_ASAP7_75t_L g15720 ( 
.A(n_15507),
.Y(n_15720)
);

NAND2xp5_ASAP7_75t_L g15721 ( 
.A(n_15381),
.B(n_2512),
.Y(n_15721)
);

AND2x2_ASAP7_75t_L g15722 ( 
.A(n_15334),
.B(n_2513),
.Y(n_15722)
);

AND2x2_ASAP7_75t_L g15723 ( 
.A(n_15467),
.B(n_2513),
.Y(n_15723)
);

INVx3_ASAP7_75t_L g15724 ( 
.A(n_15420),
.Y(n_15724)
);

INVx2_ASAP7_75t_L g15725 ( 
.A(n_15325),
.Y(n_15725)
);

AND2x2_ASAP7_75t_L g15726 ( 
.A(n_15417),
.B(n_15367),
.Y(n_15726)
);

INVx2_ASAP7_75t_L g15727 ( 
.A(n_15527),
.Y(n_15727)
);

AND2x2_ASAP7_75t_L g15728 ( 
.A(n_15536),
.B(n_15369),
.Y(n_15728)
);

INVx1_ASAP7_75t_L g15729 ( 
.A(n_15522),
.Y(n_15729)
);

INVx1_ASAP7_75t_L g15730 ( 
.A(n_15592),
.Y(n_15730)
);

INVx2_ASAP7_75t_SL g15731 ( 
.A(n_15589),
.Y(n_15731)
);

AND2x2_ASAP7_75t_L g15732 ( 
.A(n_15525),
.B(n_15316),
.Y(n_15732)
);

INVx1_ASAP7_75t_L g15733 ( 
.A(n_15599),
.Y(n_15733)
);

INVx2_ASAP7_75t_L g15734 ( 
.A(n_15572),
.Y(n_15734)
);

BUFx12f_ASAP7_75t_L g15735 ( 
.A(n_15587),
.Y(n_15735)
);

HB1xp67_ASAP7_75t_L g15736 ( 
.A(n_15573),
.Y(n_15736)
);

INVx1_ASAP7_75t_L g15737 ( 
.A(n_15526),
.Y(n_15737)
);

AND2x2_ASAP7_75t_L g15738 ( 
.A(n_15540),
.B(n_15282),
.Y(n_15738)
);

OR2x2_ASAP7_75t_L g15739 ( 
.A(n_15620),
.B(n_15339),
.Y(n_15739)
);

INVx2_ASAP7_75t_L g15740 ( 
.A(n_15572),
.Y(n_15740)
);

AND2x2_ASAP7_75t_L g15741 ( 
.A(n_15579),
.B(n_15305),
.Y(n_15741)
);

INVx1_ASAP7_75t_L g15742 ( 
.A(n_15575),
.Y(n_15742)
);

INVx2_ASAP7_75t_L g15743 ( 
.A(n_15561),
.Y(n_15743)
);

INVx2_ASAP7_75t_L g15744 ( 
.A(n_15582),
.Y(n_15744)
);

AND2x2_ASAP7_75t_L g15745 ( 
.A(n_15579),
.B(n_15295),
.Y(n_15745)
);

INVx1_ASAP7_75t_L g15746 ( 
.A(n_15584),
.Y(n_15746)
);

OR2x2_ASAP7_75t_L g15747 ( 
.A(n_15530),
.B(n_15389),
.Y(n_15747)
);

INVx2_ASAP7_75t_L g15748 ( 
.A(n_15605),
.Y(n_15748)
);

INVx1_ASAP7_75t_L g15749 ( 
.A(n_15529),
.Y(n_15749)
);

INVx2_ASAP7_75t_SL g15750 ( 
.A(n_15559),
.Y(n_15750)
);

AND2x2_ASAP7_75t_L g15751 ( 
.A(n_15613),
.B(n_15322),
.Y(n_15751)
);

INVx1_ASAP7_75t_L g15752 ( 
.A(n_15602),
.Y(n_15752)
);

INVx2_ASAP7_75t_L g15753 ( 
.A(n_15555),
.Y(n_15753)
);

INVx1_ASAP7_75t_L g15754 ( 
.A(n_15669),
.Y(n_15754)
);

AND2x2_ASAP7_75t_L g15755 ( 
.A(n_15552),
.B(n_15411),
.Y(n_15755)
);

INVx1_ASAP7_75t_L g15756 ( 
.A(n_15534),
.Y(n_15756)
);

NAND2xp5_ASAP7_75t_L g15757 ( 
.A(n_15700),
.B(n_15516),
.Y(n_15757)
);

NAND2xp33_ASAP7_75t_SL g15758 ( 
.A(n_15712),
.B(n_15460),
.Y(n_15758)
);

HB1xp67_ASAP7_75t_L g15759 ( 
.A(n_15651),
.Y(n_15759)
);

INVx2_ASAP7_75t_L g15760 ( 
.A(n_15553),
.Y(n_15760)
);

INVx2_ASAP7_75t_L g15761 ( 
.A(n_15596),
.Y(n_15761)
);

INVx1_ASAP7_75t_L g15762 ( 
.A(n_15563),
.Y(n_15762)
);

OR2x2_ASAP7_75t_L g15763 ( 
.A(n_15724),
.B(n_15479),
.Y(n_15763)
);

AOI22xp5_ASAP7_75t_L g15764 ( 
.A1(n_15711),
.A2(n_15301),
.B1(n_15351),
.B2(n_15391),
.Y(n_15764)
);

BUFx3_ASAP7_75t_L g15765 ( 
.A(n_15636),
.Y(n_15765)
);

NOR2x1_ASAP7_75t_L g15766 ( 
.A(n_15672),
.B(n_15509),
.Y(n_15766)
);

INVx1_ASAP7_75t_L g15767 ( 
.A(n_15657),
.Y(n_15767)
);

INVxp67_ASAP7_75t_SL g15768 ( 
.A(n_15580),
.Y(n_15768)
);

INVx1_ASAP7_75t_L g15769 ( 
.A(n_15660),
.Y(n_15769)
);

INVx1_ASAP7_75t_L g15770 ( 
.A(n_15564),
.Y(n_15770)
);

BUFx3_ASAP7_75t_L g15771 ( 
.A(n_15636),
.Y(n_15771)
);

INVx1_ASAP7_75t_L g15772 ( 
.A(n_15621),
.Y(n_15772)
);

NAND2xp5_ASAP7_75t_L g15773 ( 
.A(n_15700),
.B(n_15457),
.Y(n_15773)
);

INVx2_ASAP7_75t_SL g15774 ( 
.A(n_15528),
.Y(n_15774)
);

OR2x2_ASAP7_75t_L g15775 ( 
.A(n_15565),
.B(n_15410),
.Y(n_15775)
);

INVx1_ASAP7_75t_L g15776 ( 
.A(n_15611),
.Y(n_15776)
);

AOI22xp33_ASAP7_75t_L g15777 ( 
.A1(n_15570),
.A2(n_15317),
.B1(n_15382),
.B2(n_15373),
.Y(n_15777)
);

INVx1_ASAP7_75t_L g15778 ( 
.A(n_15547),
.Y(n_15778)
);

AOI22xp33_ASAP7_75t_L g15779 ( 
.A1(n_15625),
.A2(n_15415),
.B1(n_15430),
.B2(n_15425),
.Y(n_15779)
);

NAND2xp5_ASAP7_75t_L g15780 ( 
.A(n_15635),
.B(n_15442),
.Y(n_15780)
);

INVx1_ASAP7_75t_L g15781 ( 
.A(n_15595),
.Y(n_15781)
);

AND2x2_ASAP7_75t_L g15782 ( 
.A(n_15557),
.B(n_15414),
.Y(n_15782)
);

AND2x2_ASAP7_75t_L g15783 ( 
.A(n_15670),
.B(n_15576),
.Y(n_15783)
);

NAND2xp5_ASAP7_75t_L g15784 ( 
.A(n_15723),
.B(n_15502),
.Y(n_15784)
);

INVx1_ASAP7_75t_L g15785 ( 
.A(n_15537),
.Y(n_15785)
);

INVx2_ASAP7_75t_L g15786 ( 
.A(n_15597),
.Y(n_15786)
);

INVx1_ASAP7_75t_L g15787 ( 
.A(n_15535),
.Y(n_15787)
);

INVx2_ASAP7_75t_L g15788 ( 
.A(n_15566),
.Y(n_15788)
);

AND2x2_ASAP7_75t_L g15789 ( 
.A(n_15571),
.B(n_15517),
.Y(n_15789)
);

AND2x2_ASAP7_75t_L g15790 ( 
.A(n_15533),
.B(n_15356),
.Y(n_15790)
);

INVx1_ASAP7_75t_L g15791 ( 
.A(n_15541),
.Y(n_15791)
);

OR2x2_ASAP7_75t_L g15792 ( 
.A(n_15704),
.B(n_15428),
.Y(n_15792)
);

HB1xp67_ASAP7_75t_L g15793 ( 
.A(n_15618),
.Y(n_15793)
);

INVx1_ASAP7_75t_L g15794 ( 
.A(n_15550),
.Y(n_15794)
);

OR2x2_ASAP7_75t_L g15795 ( 
.A(n_15577),
.B(n_15471),
.Y(n_15795)
);

AND2x2_ASAP7_75t_L g15796 ( 
.A(n_15622),
.B(n_15374),
.Y(n_15796)
);

AND2x2_ASAP7_75t_L g15797 ( 
.A(n_15545),
.B(n_15405),
.Y(n_15797)
);

AOI22xp33_ASAP7_75t_L g15798 ( 
.A1(n_15714),
.A2(n_15453),
.B1(n_15499),
.B2(n_15399),
.Y(n_15798)
);

OR2x2_ASAP7_75t_L g15799 ( 
.A(n_15639),
.B(n_15333),
.Y(n_15799)
);

HB1xp67_ASAP7_75t_L g15800 ( 
.A(n_15634),
.Y(n_15800)
);

INVx1_ASAP7_75t_L g15801 ( 
.A(n_15594),
.Y(n_15801)
);

INVx3_ASAP7_75t_L g15802 ( 
.A(n_15549),
.Y(n_15802)
);

OR2x2_ASAP7_75t_L g15803 ( 
.A(n_15591),
.B(n_15484),
.Y(n_15803)
);

INVx2_ASAP7_75t_L g15804 ( 
.A(n_15551),
.Y(n_15804)
);

INVx3_ASAP7_75t_L g15805 ( 
.A(n_15523),
.Y(n_15805)
);

INVx2_ASAP7_75t_L g15806 ( 
.A(n_15524),
.Y(n_15806)
);

INVx2_ASAP7_75t_L g15807 ( 
.A(n_15568),
.Y(n_15807)
);

AND2x2_ASAP7_75t_L g15808 ( 
.A(n_15531),
.B(n_15364),
.Y(n_15808)
);

AOI22xp33_ASAP7_75t_L g15809 ( 
.A1(n_15708),
.A2(n_15349),
.B1(n_15470),
.B2(n_15508),
.Y(n_15809)
);

INVx1_ASAP7_75t_L g15810 ( 
.A(n_15675),
.Y(n_15810)
);

AND2x2_ASAP7_75t_L g15811 ( 
.A(n_15562),
.B(n_15492),
.Y(n_15811)
);

AND2x2_ASAP7_75t_L g15812 ( 
.A(n_15539),
.B(n_15469),
.Y(n_15812)
);

NAND2xp5_ASAP7_75t_L g15813 ( 
.A(n_15631),
.B(n_15510),
.Y(n_15813)
);

AND2x2_ASAP7_75t_L g15814 ( 
.A(n_15586),
.B(n_15335),
.Y(n_15814)
);

NOR2xp33_ASAP7_75t_L g15815 ( 
.A(n_15610),
.B(n_15473),
.Y(n_15815)
);

NAND2xp5_ASAP7_75t_L g15816 ( 
.A(n_15692),
.B(n_15413),
.Y(n_15816)
);

OR2x6_ASAP7_75t_SL g15817 ( 
.A(n_15532),
.B(n_15475),
.Y(n_15817)
);

HB1xp67_ASAP7_75t_L g15818 ( 
.A(n_15583),
.Y(n_15818)
);

AND2x2_ASAP7_75t_L g15819 ( 
.A(n_15615),
.B(n_15461),
.Y(n_15819)
);

AND2x2_ASAP7_75t_L g15820 ( 
.A(n_15548),
.B(n_15354),
.Y(n_15820)
);

INVx1_ASAP7_75t_L g15821 ( 
.A(n_15603),
.Y(n_15821)
);

AND2x2_ASAP7_75t_L g15822 ( 
.A(n_15709),
.B(n_15383),
.Y(n_15822)
);

INVx1_ASAP7_75t_L g15823 ( 
.A(n_15640),
.Y(n_15823)
);

AND2x2_ASAP7_75t_L g15824 ( 
.A(n_15554),
.B(n_15348),
.Y(n_15824)
);

INVx1_ASAP7_75t_L g15825 ( 
.A(n_15614),
.Y(n_15825)
);

INVx1_ASAP7_75t_L g15826 ( 
.A(n_15616),
.Y(n_15826)
);

INVxp67_ASAP7_75t_SL g15827 ( 
.A(n_15649),
.Y(n_15827)
);

INVx1_ASAP7_75t_L g15828 ( 
.A(n_15560),
.Y(n_15828)
);

INVx1_ASAP7_75t_L g15829 ( 
.A(n_15567),
.Y(n_15829)
);

BUFx3_ASAP7_75t_L g15830 ( 
.A(n_15612),
.Y(n_15830)
);

NAND2xp5_ASAP7_75t_L g15831 ( 
.A(n_15716),
.B(n_15674),
.Y(n_15831)
);

OR2x2_ASAP7_75t_L g15832 ( 
.A(n_15695),
.B(n_15513),
.Y(n_15832)
);

AND2x2_ASAP7_75t_L g15833 ( 
.A(n_15629),
.B(n_15514),
.Y(n_15833)
);

OR2x2_ASAP7_75t_L g15834 ( 
.A(n_15585),
.B(n_15387),
.Y(n_15834)
);

NAND2xp5_ASAP7_75t_L g15835 ( 
.A(n_15666),
.B(n_15396),
.Y(n_15835)
);

AND2x2_ASAP7_75t_L g15836 ( 
.A(n_15607),
.B(n_15368),
.Y(n_15836)
);

AOI22xp5_ASAP7_75t_SL g15837 ( 
.A1(n_15713),
.A2(n_15447),
.B1(n_15402),
.B2(n_15446),
.Y(n_15837)
);

INVx2_ASAP7_75t_L g15838 ( 
.A(n_15590),
.Y(n_15838)
);

NOR2xp67_ASAP7_75t_L g15839 ( 
.A(n_15656),
.B(n_15671),
.Y(n_15839)
);

AOI22xp33_ASAP7_75t_L g15840 ( 
.A1(n_15705),
.A2(n_15488),
.B1(n_15485),
.B2(n_15482),
.Y(n_15840)
);

HB1xp67_ASAP7_75t_L g15841 ( 
.A(n_15632),
.Y(n_15841)
);

INVxp67_ASAP7_75t_L g15842 ( 
.A(n_15543),
.Y(n_15842)
);

INVx1_ASAP7_75t_L g15843 ( 
.A(n_15606),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_15643),
.B(n_15642),
.Y(n_15844)
);

INVx2_ASAP7_75t_L g15845 ( 
.A(n_15604),
.Y(n_15845)
);

NAND2xp5_ASAP7_75t_L g15846 ( 
.A(n_15644),
.B(n_15449),
.Y(n_15846)
);

AOI22xp5_ASAP7_75t_L g15847 ( 
.A1(n_15652),
.A2(n_15726),
.B1(n_15546),
.B2(n_15609),
.Y(n_15847)
);

INVxp67_ASAP7_75t_SL g15848 ( 
.A(n_15680),
.Y(n_15848)
);

INVx2_ASAP7_75t_L g15849 ( 
.A(n_15581),
.Y(n_15849)
);

INVx1_ASAP7_75t_L g15850 ( 
.A(n_15633),
.Y(n_15850)
);

NOR2xp67_ASAP7_75t_L g15851 ( 
.A(n_15677),
.B(n_15353),
.Y(n_15851)
);

OR2x2_ASAP7_75t_L g15852 ( 
.A(n_15653),
.B(n_15451),
.Y(n_15852)
);

AND2x4_ASAP7_75t_L g15853 ( 
.A(n_15617),
.B(n_2514),
.Y(n_15853)
);

INVx2_ASAP7_75t_L g15854 ( 
.A(n_15623),
.Y(n_15854)
);

BUFx2_ASAP7_75t_L g15855 ( 
.A(n_15689),
.Y(n_15855)
);

INVx2_ASAP7_75t_L g15856 ( 
.A(n_15574),
.Y(n_15856)
);

OR2x2_ASAP7_75t_L g15857 ( 
.A(n_15698),
.B(n_2515),
.Y(n_15857)
);

BUFx6f_ASAP7_75t_L g15858 ( 
.A(n_15654),
.Y(n_15858)
);

INVx2_ASAP7_75t_L g15859 ( 
.A(n_15588),
.Y(n_15859)
);

INVx1_ASAP7_75t_L g15860 ( 
.A(n_15684),
.Y(n_15860)
);

NAND2xp5_ASAP7_75t_L g15861 ( 
.A(n_15715),
.B(n_2515),
.Y(n_15861)
);

INVx2_ASAP7_75t_L g15862 ( 
.A(n_15601),
.Y(n_15862)
);

AND2x4_ASAP7_75t_L g15863 ( 
.A(n_15598),
.B(n_2516),
.Y(n_15863)
);

INVx1_ASAP7_75t_L g15864 ( 
.A(n_15558),
.Y(n_15864)
);

INVx1_ASAP7_75t_L g15865 ( 
.A(n_15569),
.Y(n_15865)
);

BUFx6f_ASAP7_75t_L g15866 ( 
.A(n_15655),
.Y(n_15866)
);

AOI221xp5_ASAP7_75t_L g15867 ( 
.A1(n_15542),
.A2(n_2518),
.B1(n_2516),
.B2(n_2517),
.C(n_2519),
.Y(n_15867)
);

NAND2xp5_ASAP7_75t_L g15868 ( 
.A(n_15702),
.B(n_15664),
.Y(n_15868)
);

INVx2_ASAP7_75t_SL g15869 ( 
.A(n_15556),
.Y(n_15869)
);

AND2x2_ASAP7_75t_L g15870 ( 
.A(n_15638),
.B(n_2517),
.Y(n_15870)
);

INVx1_ASAP7_75t_L g15871 ( 
.A(n_15578),
.Y(n_15871)
);

OR2x2_ASAP7_75t_L g15872 ( 
.A(n_15703),
.B(n_2519),
.Y(n_15872)
);

INVx1_ASAP7_75t_L g15873 ( 
.A(n_15593),
.Y(n_15873)
);

NAND2xp5_ASAP7_75t_L g15874 ( 
.A(n_15694),
.B(n_2520),
.Y(n_15874)
);

AOI22xp33_ASAP7_75t_L g15875 ( 
.A1(n_15720),
.A2(n_2522),
.B1(n_2520),
.B2(n_2521),
.Y(n_15875)
);

AND2x2_ASAP7_75t_L g15876 ( 
.A(n_15701),
.B(n_2522),
.Y(n_15876)
);

NAND2xp5_ASAP7_75t_SL g15877 ( 
.A(n_15662),
.B(n_2523),
.Y(n_15877)
);

AND2x2_ASAP7_75t_L g15878 ( 
.A(n_15685),
.B(n_2523),
.Y(n_15878)
);

INVx2_ASAP7_75t_L g15879 ( 
.A(n_15662),
.Y(n_15879)
);

NAND2xp5_ASAP7_75t_L g15880 ( 
.A(n_15707),
.B(n_2524),
.Y(n_15880)
);

NAND2xp5_ASAP7_75t_L g15881 ( 
.A(n_15690),
.B(n_2525),
.Y(n_15881)
);

INVx1_ASAP7_75t_L g15882 ( 
.A(n_15619),
.Y(n_15882)
);

AND2x2_ASAP7_75t_L g15883 ( 
.A(n_15783),
.B(n_15696),
.Y(n_15883)
);

NAND2xp5_ASAP7_75t_L g15884 ( 
.A(n_15768),
.B(n_15710),
.Y(n_15884)
);

AND2x4_ASAP7_75t_L g15885 ( 
.A(n_15774),
.B(n_15691),
.Y(n_15885)
);

INVx2_ASAP7_75t_L g15886 ( 
.A(n_15750),
.Y(n_15886)
);

AND2x2_ASAP7_75t_L g15887 ( 
.A(n_15736),
.B(n_15693),
.Y(n_15887)
);

AND2x2_ASAP7_75t_L g15888 ( 
.A(n_15731),
.B(n_15745),
.Y(n_15888)
);

AND2x2_ASAP7_75t_L g15889 ( 
.A(n_15727),
.B(n_15725),
.Y(n_15889)
);

INVx1_ASAP7_75t_L g15890 ( 
.A(n_15759),
.Y(n_15890)
);

INVx2_ASAP7_75t_L g15891 ( 
.A(n_15765),
.Y(n_15891)
);

INVx1_ASAP7_75t_L g15892 ( 
.A(n_15756),
.Y(n_15892)
);

OR2x2_ASAP7_75t_L g15893 ( 
.A(n_15827),
.B(n_15538),
.Y(n_15893)
);

HB1xp67_ASAP7_75t_L g15894 ( 
.A(n_15793),
.Y(n_15894)
);

INVx1_ASAP7_75t_SL g15895 ( 
.A(n_15855),
.Y(n_15895)
);

AND2x2_ASAP7_75t_L g15896 ( 
.A(n_15741),
.B(n_15678),
.Y(n_15896)
);

INVxp33_ASAP7_75t_SL g15897 ( 
.A(n_15818),
.Y(n_15897)
);

INVx2_ASAP7_75t_L g15898 ( 
.A(n_15771),
.Y(n_15898)
);

INVx1_ASAP7_75t_L g15899 ( 
.A(n_15762),
.Y(n_15899)
);

NAND2xp5_ASAP7_75t_L g15900 ( 
.A(n_15841),
.B(n_15697),
.Y(n_15900)
);

NAND2xp5_ASAP7_75t_L g15901 ( 
.A(n_15744),
.B(n_15706),
.Y(n_15901)
);

NAND2xp5_ASAP7_75t_L g15902 ( 
.A(n_15748),
.B(n_15732),
.Y(n_15902)
);

NAND2xp5_ASAP7_75t_L g15903 ( 
.A(n_15761),
.B(n_15641),
.Y(n_15903)
);

NAND2xp5_ASAP7_75t_L g15904 ( 
.A(n_15843),
.B(n_15681),
.Y(n_15904)
);

INVx2_ASAP7_75t_L g15905 ( 
.A(n_15858),
.Y(n_15905)
);

INVx2_ASAP7_75t_L g15906 ( 
.A(n_15858),
.Y(n_15906)
);

INVx2_ASAP7_75t_L g15907 ( 
.A(n_15866),
.Y(n_15907)
);

INVx2_ASAP7_75t_L g15908 ( 
.A(n_15866),
.Y(n_15908)
);

AND2x2_ASAP7_75t_L g15909 ( 
.A(n_15738),
.B(n_15682),
.Y(n_15909)
);

NAND2xp5_ASAP7_75t_L g15910 ( 
.A(n_15734),
.B(n_15717),
.Y(n_15910)
);

OR2x2_ASAP7_75t_L g15911 ( 
.A(n_15831),
.B(n_15544),
.Y(n_15911)
);

AOI22xp33_ASAP7_75t_L g15912 ( 
.A1(n_15758),
.A2(n_15668),
.B1(n_15600),
.B2(n_15721),
.Y(n_15912)
);

AND2x2_ASAP7_75t_L g15913 ( 
.A(n_15740),
.B(n_15683),
.Y(n_15913)
);

NAND2xp5_ASAP7_75t_L g15914 ( 
.A(n_15839),
.B(n_15742),
.Y(n_15914)
);

NAND2xp5_ASAP7_75t_L g15915 ( 
.A(n_15746),
.B(n_15719),
.Y(n_15915)
);

BUFx2_ASAP7_75t_L g15916 ( 
.A(n_15735),
.Y(n_15916)
);

AND2x4_ASAP7_75t_L g15917 ( 
.A(n_15869),
.B(n_15676),
.Y(n_15917)
);

AOI22xp33_ASAP7_75t_SL g15918 ( 
.A1(n_15757),
.A2(n_15722),
.B1(n_15648),
.B2(n_15699),
.Y(n_15918)
);

INVx1_ASAP7_75t_L g15919 ( 
.A(n_15730),
.Y(n_15919)
);

HB1xp67_ASAP7_75t_L g15920 ( 
.A(n_15733),
.Y(n_15920)
);

NOR2xp33_ASAP7_75t_L g15921 ( 
.A(n_15760),
.B(n_15773),
.Y(n_15921)
);

INVx3_ASAP7_75t_L g15922 ( 
.A(n_15830),
.Y(n_15922)
);

NOR2x1_ASAP7_75t_L g15923 ( 
.A(n_15772),
.B(n_15661),
.Y(n_15923)
);

AND2x2_ASAP7_75t_L g15924 ( 
.A(n_15789),
.B(n_15673),
.Y(n_15924)
);

INVx2_ASAP7_75t_L g15925 ( 
.A(n_15805),
.Y(n_15925)
);

INVx1_ASAP7_75t_L g15926 ( 
.A(n_15729),
.Y(n_15926)
);

INVx1_ASAP7_75t_L g15927 ( 
.A(n_15844),
.Y(n_15927)
);

BUFx2_ASAP7_75t_L g15928 ( 
.A(n_15800),
.Y(n_15928)
);

NOR2xp33_ASAP7_75t_L g15929 ( 
.A(n_15775),
.B(n_15647),
.Y(n_15929)
);

INVxp67_ASAP7_75t_SL g15930 ( 
.A(n_15766),
.Y(n_15930)
);

NAND2xp5_ASAP7_75t_L g15931 ( 
.A(n_15802),
.B(n_15687),
.Y(n_15931)
);

AND2x2_ASAP7_75t_L g15932 ( 
.A(n_15751),
.B(n_15686),
.Y(n_15932)
);

HB1xp67_ASAP7_75t_L g15933 ( 
.A(n_15786),
.Y(n_15933)
);

AND2x2_ASAP7_75t_L g15934 ( 
.A(n_15807),
.B(n_15608),
.Y(n_15934)
);

AND2x2_ASAP7_75t_L g15935 ( 
.A(n_15728),
.B(n_15624),
.Y(n_15935)
);

AND2x2_ASAP7_75t_L g15936 ( 
.A(n_15743),
.B(n_15626),
.Y(n_15936)
);

INVx1_ASAP7_75t_L g15937 ( 
.A(n_15801),
.Y(n_15937)
);

AND2x2_ASAP7_75t_L g15938 ( 
.A(n_15814),
.B(n_15628),
.Y(n_15938)
);

HB1xp67_ASAP7_75t_L g15939 ( 
.A(n_15878),
.Y(n_15939)
);

OR2x2_ASAP7_75t_L g15940 ( 
.A(n_15763),
.B(n_15627),
.Y(n_15940)
);

AND2x2_ASAP7_75t_L g15941 ( 
.A(n_15753),
.B(n_15630),
.Y(n_15941)
);

INVx1_ASAP7_75t_L g15942 ( 
.A(n_15821),
.Y(n_15942)
);

NAND2xp5_ASAP7_75t_L g15943 ( 
.A(n_15796),
.B(n_15688),
.Y(n_15943)
);

NAND2xp5_ASAP7_75t_L g15944 ( 
.A(n_15870),
.B(n_15637),
.Y(n_15944)
);

INVx1_ASAP7_75t_L g15945 ( 
.A(n_15752),
.Y(n_15945)
);

INVx1_ASAP7_75t_L g15946 ( 
.A(n_15754),
.Y(n_15946)
);

AND2x2_ASAP7_75t_L g15947 ( 
.A(n_15876),
.B(n_15645),
.Y(n_15947)
);

INVx2_ASAP7_75t_L g15948 ( 
.A(n_15853),
.Y(n_15948)
);

BUFx2_ASAP7_75t_L g15949 ( 
.A(n_15848),
.Y(n_15949)
);

INVx2_ASAP7_75t_L g15950 ( 
.A(n_15863),
.Y(n_15950)
);

NAND2xp5_ASAP7_75t_L g15951 ( 
.A(n_15790),
.B(n_15646),
.Y(n_15951)
);

INVx2_ASAP7_75t_L g15952 ( 
.A(n_15788),
.Y(n_15952)
);

OR2x2_ASAP7_75t_L g15953 ( 
.A(n_15739),
.B(n_15718),
.Y(n_15953)
);

NAND2xp5_ASAP7_75t_L g15954 ( 
.A(n_15819),
.B(n_15808),
.Y(n_15954)
);

INVxp67_ASAP7_75t_SL g15955 ( 
.A(n_15877),
.Y(n_15955)
);

INVx1_ASAP7_75t_L g15956 ( 
.A(n_15810),
.Y(n_15956)
);

INVx1_ASAP7_75t_L g15957 ( 
.A(n_15823),
.Y(n_15957)
);

HB1xp67_ASAP7_75t_L g15958 ( 
.A(n_15778),
.Y(n_15958)
);

INVx1_ASAP7_75t_L g15959 ( 
.A(n_15860),
.Y(n_15959)
);

AND2x2_ASAP7_75t_L g15960 ( 
.A(n_15755),
.B(n_15650),
.Y(n_15960)
);

INVx1_ASAP7_75t_L g15961 ( 
.A(n_15767),
.Y(n_15961)
);

AND2x2_ASAP7_75t_L g15962 ( 
.A(n_15797),
.B(n_15658),
.Y(n_15962)
);

AND2x2_ASAP7_75t_L g15963 ( 
.A(n_15782),
.B(n_15659),
.Y(n_15963)
);

INVx2_ASAP7_75t_L g15964 ( 
.A(n_15806),
.Y(n_15964)
);

NAND2xp5_ASAP7_75t_L g15965 ( 
.A(n_15811),
.B(n_15663),
.Y(n_15965)
);

INVx1_ASAP7_75t_L g15966 ( 
.A(n_15769),
.Y(n_15966)
);

INVxp67_ASAP7_75t_SL g15967 ( 
.A(n_15780),
.Y(n_15967)
);

INVx1_ASAP7_75t_SL g15968 ( 
.A(n_15857),
.Y(n_15968)
);

INVx1_ASAP7_75t_L g15969 ( 
.A(n_15854),
.Y(n_15969)
);

INVx1_ASAP7_75t_L g15970 ( 
.A(n_15770),
.Y(n_15970)
);

HB1xp67_ASAP7_75t_L g15971 ( 
.A(n_15879),
.Y(n_15971)
);

INVx3_ASAP7_75t_L g15972 ( 
.A(n_15804),
.Y(n_15972)
);

NAND2xp5_ASAP7_75t_L g15973 ( 
.A(n_15812),
.B(n_15665),
.Y(n_15973)
);

INVx2_ASAP7_75t_L g15974 ( 
.A(n_15845),
.Y(n_15974)
);

INVx1_ASAP7_75t_L g15975 ( 
.A(n_15737),
.Y(n_15975)
);

NOR2xp33_ASAP7_75t_L g15976 ( 
.A(n_15784),
.B(n_15679),
.Y(n_15976)
);

BUFx2_ASAP7_75t_L g15977 ( 
.A(n_15828),
.Y(n_15977)
);

AOI22xp33_ASAP7_75t_L g15978 ( 
.A1(n_15834),
.A2(n_15667),
.B1(n_2527),
.B2(n_2525),
.Y(n_15978)
);

OR2x2_ASAP7_75t_L g15979 ( 
.A(n_15792),
.B(n_2526),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15749),
.Y(n_15980)
);

INVx2_ASAP7_75t_L g15981 ( 
.A(n_15856),
.Y(n_15981)
);

AND2x4_ASAP7_75t_L g15982 ( 
.A(n_15825),
.B(n_2526),
.Y(n_15982)
);

INVx1_ASAP7_75t_L g15983 ( 
.A(n_15776),
.Y(n_15983)
);

AND2x2_ASAP7_75t_L g15984 ( 
.A(n_15824),
.B(n_2528),
.Y(n_15984)
);

NAND2xp5_ASAP7_75t_L g15985 ( 
.A(n_15851),
.B(n_2528),
.Y(n_15985)
);

INVx2_ASAP7_75t_L g15986 ( 
.A(n_15838),
.Y(n_15986)
);

INVx3_ASAP7_75t_L g15987 ( 
.A(n_15849),
.Y(n_15987)
);

BUFx2_ASAP7_75t_L g15988 ( 
.A(n_15781),
.Y(n_15988)
);

INVx2_ASAP7_75t_L g15989 ( 
.A(n_15862),
.Y(n_15989)
);

NAND2xp5_ASAP7_75t_L g15990 ( 
.A(n_15820),
.B(n_2529),
.Y(n_15990)
);

OR2x2_ASAP7_75t_L g15991 ( 
.A(n_15795),
.B(n_2529),
.Y(n_15991)
);

AND2x2_ASAP7_75t_L g15992 ( 
.A(n_15822),
.B(n_2531),
.Y(n_15992)
);

INVx2_ASAP7_75t_L g15993 ( 
.A(n_15859),
.Y(n_15993)
);

INVx2_ASAP7_75t_L g15994 ( 
.A(n_15826),
.Y(n_15994)
);

AND2x2_ASAP7_75t_L g15995 ( 
.A(n_15836),
.B(n_2531),
.Y(n_15995)
);

AND2x4_ASAP7_75t_SL g15996 ( 
.A(n_15850),
.B(n_2532),
.Y(n_15996)
);

NAND2xp5_ASAP7_75t_L g15997 ( 
.A(n_15764),
.B(n_2533),
.Y(n_15997)
);

AND2x2_ASAP7_75t_L g15998 ( 
.A(n_15833),
.B(n_2533),
.Y(n_15998)
);

NAND2xp5_ASAP7_75t_L g15999 ( 
.A(n_15798),
.B(n_2534),
.Y(n_15999)
);

AND2x4_ASAP7_75t_L g16000 ( 
.A(n_15785),
.B(n_15872),
.Y(n_16000)
);

INVx2_ASAP7_75t_L g16001 ( 
.A(n_15787),
.Y(n_16001)
);

AND2x2_ASAP7_75t_L g16002 ( 
.A(n_15815),
.B(n_15829),
.Y(n_16002)
);

OR2x2_ASAP7_75t_L g16003 ( 
.A(n_15832),
.B(n_15813),
.Y(n_16003)
);

INVx1_ASAP7_75t_L g16004 ( 
.A(n_15861),
.Y(n_16004)
);

INVx2_ASAP7_75t_L g16005 ( 
.A(n_15791),
.Y(n_16005)
);

INVx1_ASAP7_75t_SL g16006 ( 
.A(n_15747),
.Y(n_16006)
);

INVx1_ASAP7_75t_L g16007 ( 
.A(n_15880),
.Y(n_16007)
);

AND2x2_ASAP7_75t_L g16008 ( 
.A(n_15837),
.B(n_2534),
.Y(n_16008)
);

NAND2xp5_ASAP7_75t_L g16009 ( 
.A(n_15779),
.B(n_2535),
.Y(n_16009)
);

AND2x2_ASAP7_75t_L g16010 ( 
.A(n_15842),
.B(n_2535),
.Y(n_16010)
);

HB1xp67_ASAP7_75t_L g16011 ( 
.A(n_15794),
.Y(n_16011)
);

AND2x4_ASAP7_75t_L g16012 ( 
.A(n_15882),
.B(n_2536),
.Y(n_16012)
);

NAND2xp5_ASAP7_75t_L g16013 ( 
.A(n_15847),
.B(n_2536),
.Y(n_16013)
);

INVx2_ASAP7_75t_L g16014 ( 
.A(n_15864),
.Y(n_16014)
);

AND2x2_ASAP7_75t_L g16015 ( 
.A(n_15809),
.B(n_2537),
.Y(n_16015)
);

NAND3xp33_ASAP7_75t_L g16016 ( 
.A(n_15930),
.B(n_15777),
.C(n_15867),
.Y(n_16016)
);

INVx2_ASAP7_75t_L g16017 ( 
.A(n_15916),
.Y(n_16017)
);

AND2x2_ASAP7_75t_L g16018 ( 
.A(n_15888),
.B(n_15835),
.Y(n_16018)
);

AND2x4_ASAP7_75t_L g16019 ( 
.A(n_15886),
.B(n_15865),
.Y(n_16019)
);

HB1xp67_ASAP7_75t_L g16020 ( 
.A(n_15894),
.Y(n_16020)
);

INVx2_ASAP7_75t_L g16021 ( 
.A(n_15949),
.Y(n_16021)
);

AND2x2_ASAP7_75t_L g16022 ( 
.A(n_15883),
.B(n_15840),
.Y(n_16022)
);

INVx1_ASAP7_75t_L g16023 ( 
.A(n_15890),
.Y(n_16023)
);

INVx2_ASAP7_75t_L g16024 ( 
.A(n_15922),
.Y(n_16024)
);

OR2x2_ASAP7_75t_L g16025 ( 
.A(n_15893),
.B(n_15895),
.Y(n_16025)
);

AND2x4_ASAP7_75t_L g16026 ( 
.A(n_15885),
.B(n_15871),
.Y(n_16026)
);

AND2x4_ASAP7_75t_L g16027 ( 
.A(n_15917),
.B(n_15873),
.Y(n_16027)
);

OR2x2_ASAP7_75t_L g16028 ( 
.A(n_15954),
.B(n_15852),
.Y(n_16028)
);

AOI22xp33_ASAP7_75t_L g16029 ( 
.A1(n_15897),
.A2(n_15803),
.B1(n_15799),
.B2(n_15868),
.Y(n_16029)
);

OAI33xp33_ASAP7_75t_L g16030 ( 
.A1(n_15919),
.A2(n_15846),
.A3(n_15816),
.B1(n_15881),
.B2(n_15817),
.B3(n_15874),
.Y(n_16030)
);

NAND2xp5_ASAP7_75t_L g16031 ( 
.A(n_15924),
.B(n_15875),
.Y(n_16031)
);

BUFx2_ASAP7_75t_L g16032 ( 
.A(n_15928),
.Y(n_16032)
);

AND2x2_ASAP7_75t_L g16033 ( 
.A(n_15932),
.B(n_2537),
.Y(n_16033)
);

OR2x2_ASAP7_75t_L g16034 ( 
.A(n_15915),
.B(n_2538),
.Y(n_16034)
);

AND2x2_ASAP7_75t_L g16035 ( 
.A(n_15913),
.B(n_2538),
.Y(n_16035)
);

NAND4xp25_ASAP7_75t_L g16036 ( 
.A(n_15912),
.B(n_2541),
.C(n_2539),
.D(n_2540),
.Y(n_16036)
);

BUFx2_ASAP7_75t_L g16037 ( 
.A(n_15977),
.Y(n_16037)
);

HB1xp67_ASAP7_75t_L g16038 ( 
.A(n_15958),
.Y(n_16038)
);

AND2x4_ASAP7_75t_L g16039 ( 
.A(n_15907),
.B(n_2539),
.Y(n_16039)
);

INVx2_ASAP7_75t_SL g16040 ( 
.A(n_15996),
.Y(n_16040)
);

OAI31xp33_ASAP7_75t_L g16041 ( 
.A1(n_16008),
.A2(n_2543),
.A3(n_2541),
.B(n_2542),
.Y(n_16041)
);

INVx1_ASAP7_75t_L g16042 ( 
.A(n_15920),
.Y(n_16042)
);

NOR3xp33_ASAP7_75t_SL g16043 ( 
.A(n_15921),
.B(n_2542),
.C(n_2543),
.Y(n_16043)
);

INVx2_ASAP7_75t_L g16044 ( 
.A(n_15887),
.Y(n_16044)
);

AND2x2_ASAP7_75t_L g16045 ( 
.A(n_15998),
.B(n_2544),
.Y(n_16045)
);

INVx1_ASAP7_75t_L g16046 ( 
.A(n_15939),
.Y(n_16046)
);

AND2x2_ASAP7_75t_L g16047 ( 
.A(n_15984),
.B(n_2544),
.Y(n_16047)
);

INVx2_ASAP7_75t_L g16048 ( 
.A(n_15908),
.Y(n_16048)
);

BUFx2_ASAP7_75t_L g16049 ( 
.A(n_15988),
.Y(n_16049)
);

HB1xp67_ASAP7_75t_L g16050 ( 
.A(n_15933),
.Y(n_16050)
);

INVx2_ASAP7_75t_SL g16051 ( 
.A(n_15982),
.Y(n_16051)
);

OR2x2_ASAP7_75t_L g16052 ( 
.A(n_15953),
.B(n_2545),
.Y(n_16052)
);

AND2x2_ASAP7_75t_L g16053 ( 
.A(n_15995),
.B(n_15889),
.Y(n_16053)
);

AND2x2_ASAP7_75t_L g16054 ( 
.A(n_15909),
.B(n_2545),
.Y(n_16054)
);

INVx2_ASAP7_75t_L g16055 ( 
.A(n_15905),
.Y(n_16055)
);

AND2x2_ASAP7_75t_L g16056 ( 
.A(n_15992),
.B(n_2546),
.Y(n_16056)
);

INVxp67_ASAP7_75t_SL g16057 ( 
.A(n_15923),
.Y(n_16057)
);

INVx5_ASAP7_75t_SL g16058 ( 
.A(n_16012),
.Y(n_16058)
);

INVx1_ASAP7_75t_L g16059 ( 
.A(n_15971),
.Y(n_16059)
);

BUFx6f_ASAP7_75t_L g16060 ( 
.A(n_15906),
.Y(n_16060)
);

NOR2x1_ASAP7_75t_SL g16061 ( 
.A(n_15940),
.B(n_15925),
.Y(n_16061)
);

INVx5_ASAP7_75t_L g16062 ( 
.A(n_15972),
.Y(n_16062)
);

INVx2_ASAP7_75t_L g16063 ( 
.A(n_15891),
.Y(n_16063)
);

AND2x2_ASAP7_75t_L g16064 ( 
.A(n_15962),
.B(n_2547),
.Y(n_16064)
);

NAND2xp5_ASAP7_75t_L g16065 ( 
.A(n_15918),
.B(n_2548),
.Y(n_16065)
);

INVx1_ASAP7_75t_L g16066 ( 
.A(n_15927),
.Y(n_16066)
);

AND2x2_ASAP7_75t_L g16067 ( 
.A(n_15898),
.B(n_2548),
.Y(n_16067)
);

INVx2_ASAP7_75t_L g16068 ( 
.A(n_15948),
.Y(n_16068)
);

AND2x2_ASAP7_75t_L g16069 ( 
.A(n_15935),
.B(n_2549),
.Y(n_16069)
);

INVx1_ASAP7_75t_L g16070 ( 
.A(n_15884),
.Y(n_16070)
);

AND2x2_ASAP7_75t_L g16071 ( 
.A(n_15938),
.B(n_2550),
.Y(n_16071)
);

AND2x2_ASAP7_75t_L g16072 ( 
.A(n_15896),
.B(n_2550),
.Y(n_16072)
);

AND2x2_ASAP7_75t_L g16073 ( 
.A(n_15950),
.B(n_2551),
.Y(n_16073)
);

NAND2xp5_ASAP7_75t_L g16074 ( 
.A(n_16006),
.B(n_2551),
.Y(n_16074)
);

OAI221xp5_ASAP7_75t_SL g16075 ( 
.A1(n_16003),
.A2(n_15999),
.B1(n_15943),
.B2(n_16013),
.C(n_15967),
.Y(n_16075)
);

AND2x2_ASAP7_75t_L g16076 ( 
.A(n_15934),
.B(n_2552),
.Y(n_16076)
);

AND2x2_ASAP7_75t_L g16077 ( 
.A(n_15960),
.B(n_2553),
.Y(n_16077)
);

BUFx2_ASAP7_75t_L g16078 ( 
.A(n_15955),
.Y(n_16078)
);

INVx2_ASAP7_75t_L g16079 ( 
.A(n_15987),
.Y(n_16079)
);

NAND3xp33_ASAP7_75t_SL g16080 ( 
.A(n_15968),
.B(n_2553),
.C(n_2554),
.Y(n_16080)
);

NOR2x1_ASAP7_75t_L g16081 ( 
.A(n_15914),
.B(n_2554),
.Y(n_16081)
);

INVx1_ASAP7_75t_L g16082 ( 
.A(n_15947),
.Y(n_16082)
);

INVx2_ASAP7_75t_SL g16083 ( 
.A(n_15936),
.Y(n_16083)
);

INVx2_ASAP7_75t_L g16084 ( 
.A(n_15979),
.Y(n_16084)
);

BUFx6f_ASAP7_75t_L g16085 ( 
.A(n_15964),
.Y(n_16085)
);

INVx1_ASAP7_75t_L g16086 ( 
.A(n_15944),
.Y(n_16086)
);

OAI21xp33_ASAP7_75t_L g16087 ( 
.A1(n_15929),
.A2(n_2555),
.B(n_2556),
.Y(n_16087)
);

INVx1_ASAP7_75t_L g16088 ( 
.A(n_16011),
.Y(n_16088)
);

INVx3_ASAP7_75t_L g16089 ( 
.A(n_15974),
.Y(n_16089)
);

BUFx2_ASAP7_75t_L g16090 ( 
.A(n_16000),
.Y(n_16090)
);

OR2x2_ASAP7_75t_L g16091 ( 
.A(n_15991),
.B(n_2557),
.Y(n_16091)
);

AOI22xp5_ASAP7_75t_L g16092 ( 
.A1(n_16015),
.A2(n_2560),
.B1(n_2558),
.B2(n_2559),
.Y(n_16092)
);

AO21x2_ASAP7_75t_L g16093 ( 
.A1(n_15985),
.A2(n_15997),
.B(n_16009),
.Y(n_16093)
);

INVx2_ASAP7_75t_L g16094 ( 
.A(n_15941),
.Y(n_16094)
);

NAND2xp5_ASAP7_75t_L g16095 ( 
.A(n_15892),
.B(n_2559),
.Y(n_16095)
);

OAI211xp5_ASAP7_75t_SL g16096 ( 
.A1(n_15902),
.A2(n_2562),
.B(n_2560),
.C(n_2561),
.Y(n_16096)
);

AND2x4_ASAP7_75t_L g16097 ( 
.A(n_15899),
.B(n_2561),
.Y(n_16097)
);

INVx1_ASAP7_75t_L g16098 ( 
.A(n_15963),
.Y(n_16098)
);

INVx1_ASAP7_75t_L g16099 ( 
.A(n_15901),
.Y(n_16099)
);

OAI221xp5_ASAP7_75t_L g16100 ( 
.A1(n_15978),
.A2(n_2564),
.B1(n_2562),
.B2(n_2563),
.C(n_2565),
.Y(n_16100)
);

INVx3_ASAP7_75t_L g16101 ( 
.A(n_15952),
.Y(n_16101)
);

AND2x2_ASAP7_75t_L g16102 ( 
.A(n_16002),
.B(n_2563),
.Y(n_16102)
);

AND2x4_ASAP7_75t_L g16103 ( 
.A(n_15946),
.B(n_2564),
.Y(n_16103)
);

OR2x2_ASAP7_75t_L g16104 ( 
.A(n_15900),
.B(n_2565),
.Y(n_16104)
);

INVx1_ASAP7_75t_L g16105 ( 
.A(n_15926),
.Y(n_16105)
);

INVx2_ASAP7_75t_L g16106 ( 
.A(n_15945),
.Y(n_16106)
);

AOI22xp5_ASAP7_75t_L g16107 ( 
.A1(n_15976),
.A2(n_2568),
.B1(n_2566),
.B2(n_2567),
.Y(n_16107)
);

OR2x2_ASAP7_75t_L g16108 ( 
.A(n_15911),
.B(n_2566),
.Y(n_16108)
);

NAND2xp5_ASAP7_75t_L g16109 ( 
.A(n_16010),
.B(n_2567),
.Y(n_16109)
);

INVx2_ASAP7_75t_L g16110 ( 
.A(n_15957),
.Y(n_16110)
);

OR2x2_ASAP7_75t_L g16111 ( 
.A(n_15931),
.B(n_2568),
.Y(n_16111)
);

INVx1_ASAP7_75t_L g16112 ( 
.A(n_15956),
.Y(n_16112)
);

INVx1_ASAP7_75t_L g16113 ( 
.A(n_15910),
.Y(n_16113)
);

NOR2x1_ASAP7_75t_L g16114 ( 
.A(n_15990),
.B(n_2569),
.Y(n_16114)
);

OR2x2_ASAP7_75t_L g16115 ( 
.A(n_15951),
.B(n_2569),
.Y(n_16115)
);

AND2x2_ASAP7_75t_L g16116 ( 
.A(n_15959),
.B(n_2570),
.Y(n_16116)
);

AND2x2_ASAP7_75t_L g16117 ( 
.A(n_16004),
.B(n_2570),
.Y(n_16117)
);

AND2x2_ASAP7_75t_L g16118 ( 
.A(n_16007),
.B(n_2571),
.Y(n_16118)
);

NAND2xp5_ASAP7_75t_L g16119 ( 
.A(n_15937),
.B(n_2571),
.Y(n_16119)
);

OR2x6_ASAP7_75t_L g16120 ( 
.A(n_15981),
.B(n_2572),
.Y(n_16120)
);

INVxp67_ASAP7_75t_SL g16121 ( 
.A(n_15973),
.Y(n_16121)
);

XNOR2xp5_ASAP7_75t_L g16122 ( 
.A(n_15903),
.B(n_2572),
.Y(n_16122)
);

NAND2xp5_ASAP7_75t_L g16123 ( 
.A(n_15942),
.B(n_2573),
.Y(n_16123)
);

NAND2x1p5_ASAP7_75t_SL g16124 ( 
.A(n_15994),
.B(n_2573),
.Y(n_16124)
);

HB1xp67_ASAP7_75t_L g16125 ( 
.A(n_15969),
.Y(n_16125)
);

NAND2xp5_ASAP7_75t_L g16126 ( 
.A(n_15961),
.B(n_15966),
.Y(n_16126)
);

OAI321xp33_ASAP7_75t_L g16127 ( 
.A1(n_15965),
.A2(n_15904),
.A3(n_15983),
.B1(n_15970),
.B2(n_15980),
.C(n_15975),
.Y(n_16127)
);

INVx1_ASAP7_75t_L g16128 ( 
.A(n_15986),
.Y(n_16128)
);

AND2x2_ASAP7_75t_L g16129 ( 
.A(n_15989),
.B(n_2574),
.Y(n_16129)
);

AND2x2_ASAP7_75t_L g16130 ( 
.A(n_15993),
.B(n_2574),
.Y(n_16130)
);

OAI22xp5_ASAP7_75t_L g16131 ( 
.A1(n_16014),
.A2(n_2577),
.B1(n_2575),
.B2(n_2576),
.Y(n_16131)
);

INVx1_ASAP7_75t_L g16132 ( 
.A(n_16037),
.Y(n_16132)
);

OR2x2_ASAP7_75t_L g16133 ( 
.A(n_16124),
.B(n_16001),
.Y(n_16133)
);

OR2x2_ASAP7_75t_L g16134 ( 
.A(n_16032),
.B(n_16005),
.Y(n_16134)
);

INVx3_ASAP7_75t_L g16135 ( 
.A(n_16062),
.Y(n_16135)
);

NAND2xp5_ASAP7_75t_SL g16136 ( 
.A(n_16062),
.B(n_2575),
.Y(n_16136)
);

NAND2xp5_ASAP7_75t_L g16137 ( 
.A(n_16058),
.B(n_2576),
.Y(n_16137)
);

AND2x4_ASAP7_75t_SL g16138 ( 
.A(n_16053),
.B(n_16026),
.Y(n_16138)
);

AND2x4_ASAP7_75t_L g16139 ( 
.A(n_16090),
.B(n_2577),
.Y(n_16139)
);

INVx2_ASAP7_75t_L g16140 ( 
.A(n_16061),
.Y(n_16140)
);

INVx2_ASAP7_75t_SL g16141 ( 
.A(n_16050),
.Y(n_16141)
);

NAND2xp5_ASAP7_75t_L g16142 ( 
.A(n_16040),
.B(n_2578),
.Y(n_16142)
);

INVx1_ASAP7_75t_L g16143 ( 
.A(n_16038),
.Y(n_16143)
);

INVx1_ASAP7_75t_L g16144 ( 
.A(n_16049),
.Y(n_16144)
);

AND2x2_ASAP7_75t_L g16145 ( 
.A(n_16018),
.B(n_2578),
.Y(n_16145)
);

BUFx2_ASAP7_75t_SL g16146 ( 
.A(n_16021),
.Y(n_16146)
);

INVx1_ASAP7_75t_L g16147 ( 
.A(n_16020),
.Y(n_16147)
);

INVx1_ASAP7_75t_L g16148 ( 
.A(n_16081),
.Y(n_16148)
);

NAND2xp5_ASAP7_75t_L g16149 ( 
.A(n_16057),
.B(n_16017),
.Y(n_16149)
);

INVx1_ASAP7_75t_L g16150 ( 
.A(n_16033),
.Y(n_16150)
);

OR2x2_ASAP7_75t_L g16151 ( 
.A(n_16025),
.B(n_2579),
.Y(n_16151)
);

NAND2xp5_ASAP7_75t_L g16152 ( 
.A(n_16051),
.B(n_2579),
.Y(n_16152)
);

NAND2xp5_ASAP7_75t_L g16153 ( 
.A(n_16022),
.B(n_2580),
.Y(n_16153)
);

INVx1_ASAP7_75t_L g16154 ( 
.A(n_16054),
.Y(n_16154)
);

HB1xp67_ASAP7_75t_L g16155 ( 
.A(n_16120),
.Y(n_16155)
);

INVx2_ASAP7_75t_L g16156 ( 
.A(n_16120),
.Y(n_16156)
);

INVx1_ASAP7_75t_L g16157 ( 
.A(n_16035),
.Y(n_16157)
);

NAND2xp5_ASAP7_75t_L g16158 ( 
.A(n_16027),
.B(n_2580),
.Y(n_16158)
);

AND2x4_ASAP7_75t_L g16159 ( 
.A(n_16044),
.B(n_16024),
.Y(n_16159)
);

AND2x2_ASAP7_75t_L g16160 ( 
.A(n_16078),
.B(n_2581),
.Y(n_16160)
);

NAND2xp5_ASAP7_75t_L g16161 ( 
.A(n_16056),
.B(n_2581),
.Y(n_16161)
);

AND2x2_ASAP7_75t_L g16162 ( 
.A(n_16068),
.B(n_2582),
.Y(n_16162)
);

AND2x2_ASAP7_75t_L g16163 ( 
.A(n_16098),
.B(n_2582),
.Y(n_16163)
);

AND2x2_ASAP7_75t_L g16164 ( 
.A(n_16082),
.B(n_2583),
.Y(n_16164)
);

AND2x2_ASAP7_75t_L g16165 ( 
.A(n_16072),
.B(n_2583),
.Y(n_16165)
);

AND2x4_ASAP7_75t_L g16166 ( 
.A(n_16083),
.B(n_2584),
.Y(n_16166)
);

NAND2xp5_ASAP7_75t_SL g16167 ( 
.A(n_16085),
.B(n_2584),
.Y(n_16167)
);

INVx1_ASAP7_75t_L g16168 ( 
.A(n_16064),
.Y(n_16168)
);

NAND2xp5_ASAP7_75t_L g16169 ( 
.A(n_16045),
.B(n_2585),
.Y(n_16169)
);

AND2x2_ASAP7_75t_L g16170 ( 
.A(n_16063),
.B(n_2585),
.Y(n_16170)
);

NAND2xp5_ASAP7_75t_L g16171 ( 
.A(n_16047),
.B(n_2586),
.Y(n_16171)
);

INVx1_ASAP7_75t_L g16172 ( 
.A(n_16069),
.Y(n_16172)
);

NAND2xp5_ASAP7_75t_L g16173 ( 
.A(n_16059),
.B(n_16071),
.Y(n_16173)
);

INVx3_ASAP7_75t_L g16174 ( 
.A(n_16085),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_16102),
.B(n_2586),
.Y(n_16175)
);

INVx2_ASAP7_75t_L g16176 ( 
.A(n_16060),
.Y(n_16176)
);

OR2x2_ASAP7_75t_L g16177 ( 
.A(n_16028),
.B(n_2587),
.Y(n_16177)
);

AND2x2_ASAP7_75t_L g16178 ( 
.A(n_16048),
.B(n_2587),
.Y(n_16178)
);

INVx1_ASAP7_75t_L g16179 ( 
.A(n_16077),
.Y(n_16179)
);

AND2x4_ASAP7_75t_SL g16180 ( 
.A(n_16060),
.B(n_2588),
.Y(n_16180)
);

BUFx2_ASAP7_75t_L g16181 ( 
.A(n_16114),
.Y(n_16181)
);

INVx1_ASAP7_75t_L g16182 ( 
.A(n_16076),
.Y(n_16182)
);

AND2x2_ASAP7_75t_L g16183 ( 
.A(n_16073),
.B(n_2589),
.Y(n_16183)
);

BUFx2_ASAP7_75t_L g16184 ( 
.A(n_16042),
.Y(n_16184)
);

HB1xp67_ASAP7_75t_L g16185 ( 
.A(n_16046),
.Y(n_16185)
);

OR2x2_ASAP7_75t_L g16186 ( 
.A(n_16080),
.B(n_16036),
.Y(n_16186)
);

AND2x2_ASAP7_75t_L g16187 ( 
.A(n_16055),
.B(n_2589),
.Y(n_16187)
);

NAND2xp5_ASAP7_75t_L g16188 ( 
.A(n_16029),
.B(n_16023),
.Y(n_16188)
);

AND2x2_ASAP7_75t_L g16189 ( 
.A(n_16079),
.B(n_2590),
.Y(n_16189)
);

NAND3xp33_ASAP7_75t_L g16190 ( 
.A(n_16016),
.B(n_2591),
.C(n_2592),
.Y(n_16190)
);

NAND2xp5_ASAP7_75t_L g16191 ( 
.A(n_16019),
.B(n_2591),
.Y(n_16191)
);

INVx1_ASAP7_75t_L g16192 ( 
.A(n_16052),
.Y(n_16192)
);

INVx3_ASAP7_75t_L g16193 ( 
.A(n_16039),
.Y(n_16193)
);

AND2x2_ASAP7_75t_L g16194 ( 
.A(n_16094),
.B(n_2592),
.Y(n_16194)
);

INVx2_ASAP7_75t_L g16195 ( 
.A(n_16091),
.Y(n_16195)
);

OR2x2_ASAP7_75t_L g16196 ( 
.A(n_16065),
.B(n_2593),
.Y(n_16196)
);

NAND2xp5_ASAP7_75t_L g16197 ( 
.A(n_16067),
.B(n_2594),
.Y(n_16197)
);

AND2x4_ASAP7_75t_L g16198 ( 
.A(n_16084),
.B(n_2594),
.Y(n_16198)
);

INVx1_ASAP7_75t_L g16199 ( 
.A(n_16125),
.Y(n_16199)
);

AND2x2_ASAP7_75t_L g16200 ( 
.A(n_16043),
.B(n_2595),
.Y(n_16200)
);

INVx1_ASAP7_75t_L g16201 ( 
.A(n_16108),
.Y(n_16201)
);

NAND2xp5_ASAP7_75t_L g16202 ( 
.A(n_16088),
.B(n_2595),
.Y(n_16202)
);

INVx3_ASAP7_75t_L g16203 ( 
.A(n_16089),
.Y(n_16203)
);

INVx1_ASAP7_75t_L g16204 ( 
.A(n_16116),
.Y(n_16204)
);

AND2x2_ASAP7_75t_L g16205 ( 
.A(n_16093),
.B(n_2596),
.Y(n_16205)
);

OR2x2_ASAP7_75t_L g16206 ( 
.A(n_16031),
.B(n_2596),
.Y(n_16206)
);

AND2x4_ASAP7_75t_L g16207 ( 
.A(n_16101),
.B(n_16066),
.Y(n_16207)
);

AND2x2_ASAP7_75t_L g16208 ( 
.A(n_16121),
.B(n_2597),
.Y(n_16208)
);

AND2x4_ASAP7_75t_L g16209 ( 
.A(n_16129),
.B(n_2597),
.Y(n_16209)
);

AND2x2_ASAP7_75t_L g16210 ( 
.A(n_16099),
.B(n_2598),
.Y(n_16210)
);

INVx1_ASAP7_75t_L g16211 ( 
.A(n_16130),
.Y(n_16211)
);

NOR2x1_ASAP7_75t_L g16212 ( 
.A(n_16074),
.B(n_2598),
.Y(n_16212)
);

INVx2_ASAP7_75t_L g16213 ( 
.A(n_16097),
.Y(n_16213)
);

INVx1_ASAP7_75t_L g16214 ( 
.A(n_16109),
.Y(n_16214)
);

INVx2_ASAP7_75t_L g16215 ( 
.A(n_16103),
.Y(n_16215)
);

OR3x2_ASAP7_75t_L g16216 ( 
.A(n_16034),
.B(n_2599),
.C(n_2600),
.Y(n_16216)
);

INVx1_ASAP7_75t_L g16217 ( 
.A(n_16104),
.Y(n_16217)
);

INVx2_ASAP7_75t_L g16218 ( 
.A(n_16111),
.Y(n_16218)
);

OR2x2_ASAP7_75t_SL g16219 ( 
.A(n_16115),
.B(n_2600),
.Y(n_16219)
);

AND2x2_ASAP7_75t_L g16220 ( 
.A(n_16070),
.B(n_2601),
.Y(n_16220)
);

OR2x2_ASAP7_75t_L g16221 ( 
.A(n_16128),
.B(n_2601),
.Y(n_16221)
);

INVx2_ASAP7_75t_L g16222 ( 
.A(n_16117),
.Y(n_16222)
);

OR2x2_ASAP7_75t_L g16223 ( 
.A(n_16075),
.B(n_16106),
.Y(n_16223)
);

INVxp67_ASAP7_75t_L g16224 ( 
.A(n_16118),
.Y(n_16224)
);

AND2x2_ASAP7_75t_L g16225 ( 
.A(n_16086),
.B(n_2602),
.Y(n_16225)
);

INVx1_ASAP7_75t_L g16226 ( 
.A(n_16122),
.Y(n_16226)
);

AND2x2_ASAP7_75t_L g16227 ( 
.A(n_16113),
.B(n_2602),
.Y(n_16227)
);

INVxp67_ASAP7_75t_L g16228 ( 
.A(n_16119),
.Y(n_16228)
);

INVx2_ASAP7_75t_L g16229 ( 
.A(n_16110),
.Y(n_16229)
);

AND2x2_ASAP7_75t_L g16230 ( 
.A(n_16087),
.B(n_2603),
.Y(n_16230)
);

HB1xp67_ASAP7_75t_L g16231 ( 
.A(n_16123),
.Y(n_16231)
);

INVx2_ASAP7_75t_L g16232 ( 
.A(n_16105),
.Y(n_16232)
);

AND2x2_ASAP7_75t_L g16233 ( 
.A(n_16041),
.B(n_2603),
.Y(n_16233)
);

INVx1_ASAP7_75t_L g16234 ( 
.A(n_16095),
.Y(n_16234)
);

AND2x2_ASAP7_75t_L g16235 ( 
.A(n_16112),
.B(n_2604),
.Y(n_16235)
);

AND2x2_ASAP7_75t_L g16236 ( 
.A(n_16092),
.B(n_2604),
.Y(n_16236)
);

INVx1_ASAP7_75t_L g16237 ( 
.A(n_16126),
.Y(n_16237)
);

OR2x2_ASAP7_75t_L g16238 ( 
.A(n_16100),
.B(n_2605),
.Y(n_16238)
);

NAND2x1_ASAP7_75t_L g16239 ( 
.A(n_16127),
.B(n_2605),
.Y(n_16239)
);

AND2x2_ASAP7_75t_L g16240 ( 
.A(n_16107),
.B(n_2606),
.Y(n_16240)
);

OR2x2_ASAP7_75t_L g16241 ( 
.A(n_16131),
.B(n_2607),
.Y(n_16241)
);

AND2x4_ASAP7_75t_SL g16242 ( 
.A(n_16030),
.B(n_2607),
.Y(n_16242)
);

AND2x2_ASAP7_75t_L g16243 ( 
.A(n_16096),
.B(n_2608),
.Y(n_16243)
);

OR2x6_ASAP7_75t_L g16244 ( 
.A(n_16090),
.B(n_2608),
.Y(n_16244)
);

AOI211xp5_ASAP7_75t_L g16245 ( 
.A1(n_16016),
.A2(n_2611),
.B(n_2609),
.C(n_2610),
.Y(n_16245)
);

INVx1_ASAP7_75t_L g16246 ( 
.A(n_16037),
.Y(n_16246)
);

INVx1_ASAP7_75t_L g16247 ( 
.A(n_16037),
.Y(n_16247)
);

AND2x4_ASAP7_75t_L g16248 ( 
.A(n_16090),
.B(n_2610),
.Y(n_16248)
);

INVx1_ASAP7_75t_L g16249 ( 
.A(n_16037),
.Y(n_16249)
);

NAND2xp5_ASAP7_75t_SL g16250 ( 
.A(n_16062),
.B(n_2612),
.Y(n_16250)
);

INVx1_ASAP7_75t_L g16251 ( 
.A(n_16037),
.Y(n_16251)
);

INVxp67_ASAP7_75t_SL g16252 ( 
.A(n_16061),
.Y(n_16252)
);

HB1xp67_ASAP7_75t_L g16253 ( 
.A(n_16062),
.Y(n_16253)
);

AND2x4_ASAP7_75t_L g16254 ( 
.A(n_16090),
.B(n_2612),
.Y(n_16254)
);

INVx1_ASAP7_75t_L g16255 ( 
.A(n_16037),
.Y(n_16255)
);

INVx2_ASAP7_75t_L g16256 ( 
.A(n_16061),
.Y(n_16256)
);

AND2x2_ASAP7_75t_L g16257 ( 
.A(n_16090),
.B(n_2613),
.Y(n_16257)
);

INVx2_ASAP7_75t_SL g16258 ( 
.A(n_16138),
.Y(n_16258)
);

NOR2x1_ASAP7_75t_L g16259 ( 
.A(n_16140),
.B(n_2614),
.Y(n_16259)
);

INVxp67_ASAP7_75t_L g16260 ( 
.A(n_16252),
.Y(n_16260)
);

HB1xp67_ASAP7_75t_L g16261 ( 
.A(n_16244),
.Y(n_16261)
);

AND2x2_ASAP7_75t_L g16262 ( 
.A(n_16146),
.B(n_2614),
.Y(n_16262)
);

AND2x2_ASAP7_75t_L g16263 ( 
.A(n_16193),
.B(n_2615),
.Y(n_16263)
);

AND2x4_ASAP7_75t_SL g16264 ( 
.A(n_16159),
.B(n_2615),
.Y(n_16264)
);

OR2x2_ASAP7_75t_L g16265 ( 
.A(n_16148),
.B(n_2616),
.Y(n_16265)
);

NOR2xp33_ASAP7_75t_L g16266 ( 
.A(n_16181),
.B(n_2616),
.Y(n_16266)
);

INVx1_ASAP7_75t_L g16267 ( 
.A(n_16253),
.Y(n_16267)
);

OR2x2_ASAP7_75t_L g16268 ( 
.A(n_16244),
.B(n_2617),
.Y(n_16268)
);

INVx1_ASAP7_75t_L g16269 ( 
.A(n_16257),
.Y(n_16269)
);

INVx2_ASAP7_75t_L g16270 ( 
.A(n_16135),
.Y(n_16270)
);

INVx1_ASAP7_75t_L g16271 ( 
.A(n_16155),
.Y(n_16271)
);

OR2x2_ASAP7_75t_L g16272 ( 
.A(n_16219),
.B(n_2618),
.Y(n_16272)
);

HB1xp67_ASAP7_75t_L g16273 ( 
.A(n_16256),
.Y(n_16273)
);

INVx1_ASAP7_75t_L g16274 ( 
.A(n_16137),
.Y(n_16274)
);

AND2x4_ASAP7_75t_L g16275 ( 
.A(n_16141),
.B(n_2618),
.Y(n_16275)
);

INVx1_ASAP7_75t_L g16276 ( 
.A(n_16160),
.Y(n_16276)
);

AND2x2_ASAP7_75t_L g16277 ( 
.A(n_16145),
.B(n_2619),
.Y(n_16277)
);

AND2x2_ASAP7_75t_L g16278 ( 
.A(n_16132),
.B(n_2619),
.Y(n_16278)
);

HB1xp67_ASAP7_75t_L g16279 ( 
.A(n_16139),
.Y(n_16279)
);

NAND2xp5_ASAP7_75t_L g16280 ( 
.A(n_16248),
.B(n_2620),
.Y(n_16280)
);

INVx1_ASAP7_75t_L g16281 ( 
.A(n_16185),
.Y(n_16281)
);

INVx2_ASAP7_75t_L g16282 ( 
.A(n_16254),
.Y(n_16282)
);

AND2x2_ASAP7_75t_L g16283 ( 
.A(n_16144),
.B(n_2620),
.Y(n_16283)
);

AND2x4_ASAP7_75t_L g16284 ( 
.A(n_16156),
.B(n_2621),
.Y(n_16284)
);

AND2x4_ASAP7_75t_L g16285 ( 
.A(n_16246),
.B(n_2621),
.Y(n_16285)
);

AND2x2_ASAP7_75t_L g16286 ( 
.A(n_16247),
.B(n_2622),
.Y(n_16286)
);

INVx1_ASAP7_75t_L g16287 ( 
.A(n_16184),
.Y(n_16287)
);

INVx1_ASAP7_75t_L g16288 ( 
.A(n_16205),
.Y(n_16288)
);

INVx1_ASAP7_75t_L g16289 ( 
.A(n_16249),
.Y(n_16289)
);

INVx2_ASAP7_75t_L g16290 ( 
.A(n_16180),
.Y(n_16290)
);

INVx1_ASAP7_75t_L g16291 ( 
.A(n_16251),
.Y(n_16291)
);

INVx1_ASAP7_75t_L g16292 ( 
.A(n_16255),
.Y(n_16292)
);

INVxp67_ASAP7_75t_L g16293 ( 
.A(n_16136),
.Y(n_16293)
);

OR2x2_ASAP7_75t_L g16294 ( 
.A(n_16133),
.B(n_2622),
.Y(n_16294)
);

OR2x6_ASAP7_75t_L g16295 ( 
.A(n_16149),
.B(n_2623),
.Y(n_16295)
);

AND2x2_ASAP7_75t_L g16296 ( 
.A(n_16200),
.B(n_2623),
.Y(n_16296)
);

INVxp33_ASAP7_75t_L g16297 ( 
.A(n_16212),
.Y(n_16297)
);

BUFx2_ASAP7_75t_L g16298 ( 
.A(n_16166),
.Y(n_16298)
);

OR2x6_ASAP7_75t_L g16299 ( 
.A(n_16134),
.B(n_2624),
.Y(n_16299)
);

INVx1_ASAP7_75t_L g16300 ( 
.A(n_16151),
.Y(n_16300)
);

INVx2_ASAP7_75t_L g16301 ( 
.A(n_16175),
.Y(n_16301)
);

AND2x2_ASAP7_75t_L g16302 ( 
.A(n_16213),
.B(n_2624),
.Y(n_16302)
);

INVx2_ASAP7_75t_L g16303 ( 
.A(n_16183),
.Y(n_16303)
);

INVxp67_ASAP7_75t_L g16304 ( 
.A(n_16250),
.Y(n_16304)
);

AND2x2_ASAP7_75t_L g16305 ( 
.A(n_16215),
.B(n_2625),
.Y(n_16305)
);

NAND2xp5_ASAP7_75t_L g16306 ( 
.A(n_16242),
.B(n_2625),
.Y(n_16306)
);

INVx2_ASAP7_75t_L g16307 ( 
.A(n_16165),
.Y(n_16307)
);

OR2x2_ASAP7_75t_L g16308 ( 
.A(n_16186),
.B(n_16239),
.Y(n_16308)
);

AND2x2_ASAP7_75t_L g16309 ( 
.A(n_16176),
.B(n_2626),
.Y(n_16309)
);

INVx1_ASAP7_75t_L g16310 ( 
.A(n_16142),
.Y(n_16310)
);

INVx2_ASAP7_75t_L g16311 ( 
.A(n_16209),
.Y(n_16311)
);

AND2x2_ASAP7_75t_L g16312 ( 
.A(n_16150),
.B(n_2626),
.Y(n_16312)
);

OR2x2_ASAP7_75t_L g16313 ( 
.A(n_16177),
.B(n_2627),
.Y(n_16313)
);

AND2x2_ASAP7_75t_L g16314 ( 
.A(n_16182),
.B(n_2627),
.Y(n_16314)
);

AND2x2_ASAP7_75t_L g16315 ( 
.A(n_16157),
.B(n_2628),
.Y(n_16315)
);

NAND2xp5_ASAP7_75t_L g16316 ( 
.A(n_16147),
.B(n_2629),
.Y(n_16316)
);

AND2x4_ASAP7_75t_L g16317 ( 
.A(n_16154),
.B(n_2629),
.Y(n_16317)
);

NAND2xp5_ASAP7_75t_L g16318 ( 
.A(n_16203),
.B(n_2630),
.Y(n_16318)
);

AND2x2_ASAP7_75t_L g16319 ( 
.A(n_16174),
.B(n_2630),
.Y(n_16319)
);

INVx1_ASAP7_75t_SL g16320 ( 
.A(n_16208),
.Y(n_16320)
);

INVx1_ASAP7_75t_L g16321 ( 
.A(n_16158),
.Y(n_16321)
);

INVxp67_ASAP7_75t_L g16322 ( 
.A(n_16243),
.Y(n_16322)
);

AND2x2_ASAP7_75t_L g16323 ( 
.A(n_16168),
.B(n_2631),
.Y(n_16323)
);

INVx1_ASAP7_75t_L g16324 ( 
.A(n_16163),
.Y(n_16324)
);

AND2x2_ASAP7_75t_L g16325 ( 
.A(n_16172),
.B(n_2632),
.Y(n_16325)
);

AND2x2_ASAP7_75t_L g16326 ( 
.A(n_16179),
.B(n_2632),
.Y(n_16326)
);

INVx2_ASAP7_75t_L g16327 ( 
.A(n_16198),
.Y(n_16327)
);

OR2x2_ASAP7_75t_L g16328 ( 
.A(n_16173),
.B(n_2633),
.Y(n_16328)
);

INVx1_ASAP7_75t_L g16329 ( 
.A(n_16164),
.Y(n_16329)
);

OR2x2_ASAP7_75t_L g16330 ( 
.A(n_16153),
.B(n_2634),
.Y(n_16330)
);

NAND2xp5_ASAP7_75t_L g16331 ( 
.A(n_16143),
.B(n_2634),
.Y(n_16331)
);

INVx2_ASAP7_75t_L g16332 ( 
.A(n_16207),
.Y(n_16332)
);

INVx2_ASAP7_75t_L g16333 ( 
.A(n_16221),
.Y(n_16333)
);

INVx1_ASAP7_75t_L g16334 ( 
.A(n_16152),
.Y(n_16334)
);

NAND2xp5_ASAP7_75t_L g16335 ( 
.A(n_16199),
.B(n_16162),
.Y(n_16335)
);

INVx1_ASAP7_75t_L g16336 ( 
.A(n_16178),
.Y(n_16336)
);

NAND2xp5_ASAP7_75t_L g16337 ( 
.A(n_16187),
.B(n_2635),
.Y(n_16337)
);

NAND2xp5_ASAP7_75t_L g16338 ( 
.A(n_16194),
.B(n_2635),
.Y(n_16338)
);

INVx1_ASAP7_75t_L g16339 ( 
.A(n_16170),
.Y(n_16339)
);

INVx1_ASAP7_75t_L g16340 ( 
.A(n_16191),
.Y(n_16340)
);

INVx2_ASAP7_75t_L g16341 ( 
.A(n_16189),
.Y(n_16341)
);

AND2x2_ASAP7_75t_L g16342 ( 
.A(n_16222),
.B(n_2636),
.Y(n_16342)
);

NAND2x1_ASAP7_75t_SL g16343 ( 
.A(n_16233),
.B(n_2637),
.Y(n_16343)
);

AND2x4_ASAP7_75t_L g16344 ( 
.A(n_16195),
.B(n_2638),
.Y(n_16344)
);

NAND2xp5_ASAP7_75t_L g16345 ( 
.A(n_16204),
.B(n_2638),
.Y(n_16345)
);

INVx1_ASAP7_75t_L g16346 ( 
.A(n_16161),
.Y(n_16346)
);

NOR2x1p5_ASAP7_75t_L g16347 ( 
.A(n_16188),
.B(n_16223),
.Y(n_16347)
);

INVx1_ASAP7_75t_L g16348 ( 
.A(n_16169),
.Y(n_16348)
);

INVx2_ASAP7_75t_L g16349 ( 
.A(n_16216),
.Y(n_16349)
);

NAND2xp5_ASAP7_75t_L g16350 ( 
.A(n_16192),
.B(n_2639),
.Y(n_16350)
);

INVx1_ASAP7_75t_L g16351 ( 
.A(n_16171),
.Y(n_16351)
);

OR2x2_ASAP7_75t_L g16352 ( 
.A(n_16206),
.B(n_2639),
.Y(n_16352)
);

INVx1_ASAP7_75t_L g16353 ( 
.A(n_16235),
.Y(n_16353)
);

OR2x6_ASAP7_75t_L g16354 ( 
.A(n_16218),
.B(n_2640),
.Y(n_16354)
);

NOR2xp33_ASAP7_75t_L g16355 ( 
.A(n_16224),
.B(n_2640),
.Y(n_16355)
);

INVx1_ASAP7_75t_L g16356 ( 
.A(n_16197),
.Y(n_16356)
);

AND2x2_ASAP7_75t_L g16357 ( 
.A(n_16211),
.B(n_2641),
.Y(n_16357)
);

OR2x2_ASAP7_75t_L g16358 ( 
.A(n_16241),
.B(n_2641),
.Y(n_16358)
);

INVx1_ASAP7_75t_L g16359 ( 
.A(n_16210),
.Y(n_16359)
);

AND2x2_ASAP7_75t_L g16360 ( 
.A(n_16226),
.B(n_2642),
.Y(n_16360)
);

AND2x2_ASAP7_75t_L g16361 ( 
.A(n_16201),
.B(n_2642),
.Y(n_16361)
);

HB1xp67_ASAP7_75t_L g16362 ( 
.A(n_16167),
.Y(n_16362)
);

INVx1_ASAP7_75t_L g16363 ( 
.A(n_16225),
.Y(n_16363)
);

INVx1_ASAP7_75t_L g16364 ( 
.A(n_16220),
.Y(n_16364)
);

AND2x2_ASAP7_75t_L g16365 ( 
.A(n_16236),
.B(n_2643),
.Y(n_16365)
);

INVx1_ASAP7_75t_L g16366 ( 
.A(n_16227),
.Y(n_16366)
);

AND2x2_ASAP7_75t_L g16367 ( 
.A(n_16240),
.B(n_2643),
.Y(n_16367)
);

NAND2xp5_ASAP7_75t_L g16368 ( 
.A(n_16230),
.B(n_2644),
.Y(n_16368)
);

AND2x2_ASAP7_75t_L g16369 ( 
.A(n_16217),
.B(n_2644),
.Y(n_16369)
);

OR2x2_ASAP7_75t_L g16370 ( 
.A(n_16196),
.B(n_2645),
.Y(n_16370)
);

INVx1_ASAP7_75t_L g16371 ( 
.A(n_16202),
.Y(n_16371)
);

NAND2x1p5_ASAP7_75t_L g16372 ( 
.A(n_16229),
.B(n_2645),
.Y(n_16372)
);

AND2x2_ASAP7_75t_L g16373 ( 
.A(n_16214),
.B(n_2646),
.Y(n_16373)
);

INVx2_ASAP7_75t_L g16374 ( 
.A(n_16232),
.Y(n_16374)
);

INVx1_ASAP7_75t_L g16375 ( 
.A(n_16231),
.Y(n_16375)
);

NAND2xp5_ASAP7_75t_L g16376 ( 
.A(n_16245),
.B(n_2646),
.Y(n_16376)
);

OR2x2_ASAP7_75t_L g16377 ( 
.A(n_16238),
.B(n_2647),
.Y(n_16377)
);

INVx1_ASAP7_75t_L g16378 ( 
.A(n_16190),
.Y(n_16378)
);

HB1xp67_ASAP7_75t_L g16379 ( 
.A(n_16237),
.Y(n_16379)
);

INVx1_ASAP7_75t_L g16380 ( 
.A(n_16234),
.Y(n_16380)
);

INVx3_ASAP7_75t_L g16381 ( 
.A(n_16228),
.Y(n_16381)
);

AND2x2_ASAP7_75t_L g16382 ( 
.A(n_16138),
.B(n_2647),
.Y(n_16382)
);

NAND3xp33_ASAP7_75t_L g16383 ( 
.A(n_16140),
.B(n_2648),
.C(n_2649),
.Y(n_16383)
);

INVx1_ASAP7_75t_L g16384 ( 
.A(n_16181),
.Y(n_16384)
);

INVx1_ASAP7_75t_L g16385 ( 
.A(n_16181),
.Y(n_16385)
);

INVx2_ASAP7_75t_L g16386 ( 
.A(n_16135),
.Y(n_16386)
);

INVx1_ASAP7_75t_L g16387 ( 
.A(n_16181),
.Y(n_16387)
);

INVx2_ASAP7_75t_SL g16388 ( 
.A(n_16138),
.Y(n_16388)
);

INVx1_ASAP7_75t_L g16389 ( 
.A(n_16181),
.Y(n_16389)
);

INVx1_ASAP7_75t_L g16390 ( 
.A(n_16181),
.Y(n_16390)
);

INVx1_ASAP7_75t_L g16391 ( 
.A(n_16181),
.Y(n_16391)
);

AND2x2_ASAP7_75t_L g16392 ( 
.A(n_16138),
.B(n_2650),
.Y(n_16392)
);

INVx1_ASAP7_75t_L g16393 ( 
.A(n_16181),
.Y(n_16393)
);

NAND2xp5_ASAP7_75t_L g16394 ( 
.A(n_16252),
.B(n_2651),
.Y(n_16394)
);

NAND2xp5_ASAP7_75t_L g16395 ( 
.A(n_16252),
.B(n_2651),
.Y(n_16395)
);

NOR2x1_ASAP7_75t_SL g16396 ( 
.A(n_16244),
.B(n_2652),
.Y(n_16396)
);

NAND2xp5_ASAP7_75t_L g16397 ( 
.A(n_16252),
.B(n_2652),
.Y(n_16397)
);

AND2x2_ASAP7_75t_L g16398 ( 
.A(n_16138),
.B(n_2653),
.Y(n_16398)
);

INVx3_ASAP7_75t_L g16399 ( 
.A(n_16138),
.Y(n_16399)
);

NAND2xp5_ASAP7_75t_L g16400 ( 
.A(n_16252),
.B(n_2654),
.Y(n_16400)
);

AND2x2_ASAP7_75t_L g16401 ( 
.A(n_16138),
.B(n_2654),
.Y(n_16401)
);

NAND2x1_ASAP7_75t_SL g16402 ( 
.A(n_16253),
.B(n_2655),
.Y(n_16402)
);

AND2x2_ASAP7_75t_L g16403 ( 
.A(n_16138),
.B(n_2655),
.Y(n_16403)
);

INVx1_ASAP7_75t_L g16404 ( 
.A(n_16181),
.Y(n_16404)
);

INVx1_ASAP7_75t_L g16405 ( 
.A(n_16181),
.Y(n_16405)
);

NOR2xp33_ASAP7_75t_L g16406 ( 
.A(n_16148),
.B(n_2656),
.Y(n_16406)
);

OR2x2_ASAP7_75t_L g16407 ( 
.A(n_16148),
.B(n_2656),
.Y(n_16407)
);

AND2x2_ASAP7_75t_L g16408 ( 
.A(n_16138),
.B(n_2657),
.Y(n_16408)
);

INVx2_ASAP7_75t_L g16409 ( 
.A(n_16135),
.Y(n_16409)
);

INVx1_ASAP7_75t_L g16410 ( 
.A(n_16402),
.Y(n_16410)
);

INVx2_ASAP7_75t_SL g16411 ( 
.A(n_16264),
.Y(n_16411)
);

INVx2_ASAP7_75t_L g16412 ( 
.A(n_16399),
.Y(n_16412)
);

INVx1_ASAP7_75t_L g16413 ( 
.A(n_16396),
.Y(n_16413)
);

NOR2x1p5_ASAP7_75t_SL g16414 ( 
.A(n_16308),
.B(n_2657),
.Y(n_16414)
);

AND2x2_ASAP7_75t_L g16415 ( 
.A(n_16258),
.B(n_2658),
.Y(n_16415)
);

AOI22xp5_ASAP7_75t_L g16416 ( 
.A1(n_16388),
.A2(n_16260),
.B1(n_16271),
.B2(n_16347),
.Y(n_16416)
);

INVx1_ASAP7_75t_L g16417 ( 
.A(n_16261),
.Y(n_16417)
);

INVx1_ASAP7_75t_L g16418 ( 
.A(n_16279),
.Y(n_16418)
);

INVx1_ASAP7_75t_L g16419 ( 
.A(n_16273),
.Y(n_16419)
);

INVx1_ASAP7_75t_L g16420 ( 
.A(n_16382),
.Y(n_16420)
);

INVx1_ASAP7_75t_L g16421 ( 
.A(n_16392),
.Y(n_16421)
);

INVxp67_ASAP7_75t_L g16422 ( 
.A(n_16259),
.Y(n_16422)
);

NAND2xp5_ASAP7_75t_SL g16423 ( 
.A(n_16287),
.B(n_2658),
.Y(n_16423)
);

OR2x2_ASAP7_75t_L g16424 ( 
.A(n_16306),
.B(n_2659),
.Y(n_16424)
);

NAND2xp5_ASAP7_75t_L g16425 ( 
.A(n_16398),
.B(n_2659),
.Y(n_16425)
);

INVx2_ASAP7_75t_L g16426 ( 
.A(n_16401),
.Y(n_16426)
);

BUFx2_ASAP7_75t_L g16427 ( 
.A(n_16299),
.Y(n_16427)
);

INVx1_ASAP7_75t_L g16428 ( 
.A(n_16403),
.Y(n_16428)
);

HB1xp67_ASAP7_75t_L g16429 ( 
.A(n_16299),
.Y(n_16429)
);

INVx1_ASAP7_75t_L g16430 ( 
.A(n_16408),
.Y(n_16430)
);

NAND2xp5_ASAP7_75t_L g16431 ( 
.A(n_16262),
.B(n_2660),
.Y(n_16431)
);

NAND2xp5_ASAP7_75t_SL g16432 ( 
.A(n_16297),
.B(n_2660),
.Y(n_16432)
);

OR2x2_ASAP7_75t_L g16433 ( 
.A(n_16298),
.B(n_2661),
.Y(n_16433)
);

OR2x2_ASAP7_75t_L g16434 ( 
.A(n_16294),
.B(n_16272),
.Y(n_16434)
);

INVx1_ASAP7_75t_L g16435 ( 
.A(n_16268),
.Y(n_16435)
);

AND2x2_ASAP7_75t_L g16436 ( 
.A(n_16282),
.B(n_2662),
.Y(n_16436)
);

INVx1_ASAP7_75t_L g16437 ( 
.A(n_16263),
.Y(n_16437)
);

INVx1_ASAP7_75t_L g16438 ( 
.A(n_16394),
.Y(n_16438)
);

OR2x2_ASAP7_75t_L g16439 ( 
.A(n_16395),
.B(n_2663),
.Y(n_16439)
);

OR2x6_ASAP7_75t_L g16440 ( 
.A(n_16332),
.B(n_2663),
.Y(n_16440)
);

AND2x2_ASAP7_75t_L g16441 ( 
.A(n_16296),
.B(n_2664),
.Y(n_16441)
);

OR2x2_ASAP7_75t_L g16442 ( 
.A(n_16397),
.B(n_2664),
.Y(n_16442)
);

INVx1_ASAP7_75t_L g16443 ( 
.A(n_16400),
.Y(n_16443)
);

INVx2_ASAP7_75t_L g16444 ( 
.A(n_16372),
.Y(n_16444)
);

NOR2x1_ASAP7_75t_L g16445 ( 
.A(n_16383),
.B(n_2665),
.Y(n_16445)
);

NOR3xp33_ASAP7_75t_L g16446 ( 
.A(n_16322),
.B(n_2665),
.C(n_2666),
.Y(n_16446)
);

INVx1_ASAP7_75t_L g16447 ( 
.A(n_16267),
.Y(n_16447)
);

AOI22xp5_ASAP7_75t_L g16448 ( 
.A1(n_16349),
.A2(n_2668),
.B1(n_2666),
.B2(n_2667),
.Y(n_16448)
);

AND2x2_ASAP7_75t_L g16449 ( 
.A(n_16270),
.B(n_2667),
.Y(n_16449)
);

INVx1_ASAP7_75t_L g16450 ( 
.A(n_16277),
.Y(n_16450)
);

NAND2xp5_ASAP7_75t_SL g16451 ( 
.A(n_16281),
.B(n_16275),
.Y(n_16451)
);

NAND2xp5_ASAP7_75t_L g16452 ( 
.A(n_16320),
.B(n_2668),
.Y(n_16452)
);

INVx1_ASAP7_75t_L g16453 ( 
.A(n_16302),
.Y(n_16453)
);

INVx1_ASAP7_75t_L g16454 ( 
.A(n_16305),
.Y(n_16454)
);

AND2x2_ASAP7_75t_L g16455 ( 
.A(n_16386),
.B(n_2669),
.Y(n_16455)
);

NAND2xp5_ASAP7_75t_L g16456 ( 
.A(n_16288),
.B(n_2669),
.Y(n_16456)
);

OR2x2_ASAP7_75t_L g16457 ( 
.A(n_16409),
.B(n_2670),
.Y(n_16457)
);

AND2x2_ASAP7_75t_L g16458 ( 
.A(n_16269),
.B(n_16301),
.Y(n_16458)
);

INVx1_ASAP7_75t_L g16459 ( 
.A(n_16265),
.Y(n_16459)
);

AOI222xp33_ASAP7_75t_L g16460 ( 
.A1(n_16384),
.A2(n_2672),
.B1(n_2674),
.B2(n_2670),
.C1(n_2671),
.C2(n_2673),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_16407),
.Y(n_16461)
);

INVx1_ASAP7_75t_L g16462 ( 
.A(n_16343),
.Y(n_16462)
);

INVx3_ASAP7_75t_L g16463 ( 
.A(n_16285),
.Y(n_16463)
);

AND2x4_ASAP7_75t_L g16464 ( 
.A(n_16307),
.B(n_2671),
.Y(n_16464)
);

NOR2xp33_ASAP7_75t_L g16465 ( 
.A(n_16293),
.B(n_2672),
.Y(n_16465)
);

INVx1_ASAP7_75t_L g16466 ( 
.A(n_16278),
.Y(n_16466)
);

INVx2_ASAP7_75t_L g16467 ( 
.A(n_16354),
.Y(n_16467)
);

NAND2xp5_ASAP7_75t_L g16468 ( 
.A(n_16344),
.B(n_2674),
.Y(n_16468)
);

INVx1_ASAP7_75t_L g16469 ( 
.A(n_16283),
.Y(n_16469)
);

INVx2_ASAP7_75t_L g16470 ( 
.A(n_16354),
.Y(n_16470)
);

INVx1_ASAP7_75t_L g16471 ( 
.A(n_16286),
.Y(n_16471)
);

OR2x2_ASAP7_75t_L g16472 ( 
.A(n_16358),
.B(n_2675),
.Y(n_16472)
);

NOR2xp67_ASAP7_75t_L g16473 ( 
.A(n_16304),
.B(n_2675),
.Y(n_16473)
);

NAND2xp5_ASAP7_75t_L g16474 ( 
.A(n_16284),
.B(n_2676),
.Y(n_16474)
);

INVxp67_ASAP7_75t_SL g16475 ( 
.A(n_16266),
.Y(n_16475)
);

AND2x2_ASAP7_75t_L g16476 ( 
.A(n_16303),
.B(n_2676),
.Y(n_16476)
);

AND2x2_ASAP7_75t_L g16477 ( 
.A(n_16311),
.B(n_2677),
.Y(n_16477)
);

INVx3_ASAP7_75t_L g16478 ( 
.A(n_16317),
.Y(n_16478)
);

INVx1_ASAP7_75t_L g16479 ( 
.A(n_16312),
.Y(n_16479)
);

NAND2xp5_ASAP7_75t_L g16480 ( 
.A(n_16314),
.B(n_16315),
.Y(n_16480)
);

OR2x6_ASAP7_75t_L g16481 ( 
.A(n_16290),
.B(n_16385),
.Y(n_16481)
);

AND2x2_ASAP7_75t_L g16482 ( 
.A(n_16276),
.B(n_2677),
.Y(n_16482)
);

INVxp67_ASAP7_75t_L g16483 ( 
.A(n_16406),
.Y(n_16483)
);

OR2x6_ASAP7_75t_L g16484 ( 
.A(n_16387),
.B(n_16389),
.Y(n_16484)
);

AND2x2_ASAP7_75t_L g16485 ( 
.A(n_16360),
.B(n_2678),
.Y(n_16485)
);

INVx2_ASAP7_75t_L g16486 ( 
.A(n_16295),
.Y(n_16486)
);

AND2x2_ASAP7_75t_L g16487 ( 
.A(n_16327),
.B(n_2679),
.Y(n_16487)
);

OAI211xp5_ASAP7_75t_L g16488 ( 
.A1(n_16390),
.A2(n_2681),
.B(n_2679),
.C(n_2680),
.Y(n_16488)
);

INVx1_ASAP7_75t_L g16489 ( 
.A(n_16323),
.Y(n_16489)
);

OAI21xp33_ASAP7_75t_L g16490 ( 
.A1(n_16289),
.A2(n_2680),
.B(n_2681),
.Y(n_16490)
);

INVx1_ASAP7_75t_L g16491 ( 
.A(n_16325),
.Y(n_16491)
);

INVx1_ASAP7_75t_L g16492 ( 
.A(n_16326),
.Y(n_16492)
);

AND2x2_ASAP7_75t_L g16493 ( 
.A(n_16324),
.B(n_2682),
.Y(n_16493)
);

INVxp67_ASAP7_75t_SL g16494 ( 
.A(n_16280),
.Y(n_16494)
);

INVx1_ASAP7_75t_L g16495 ( 
.A(n_16319),
.Y(n_16495)
);

NAND2xp5_ASAP7_75t_L g16496 ( 
.A(n_16361),
.B(n_2682),
.Y(n_16496)
);

INVx1_ASAP7_75t_L g16497 ( 
.A(n_16357),
.Y(n_16497)
);

INVx2_ASAP7_75t_L g16498 ( 
.A(n_16295),
.Y(n_16498)
);

INVx1_ASAP7_75t_L g16499 ( 
.A(n_16313),
.Y(n_16499)
);

INVx1_ASAP7_75t_L g16500 ( 
.A(n_16342),
.Y(n_16500)
);

OR2x2_ASAP7_75t_SL g16501 ( 
.A(n_16362),
.B(n_2683),
.Y(n_16501)
);

INVx1_ASAP7_75t_L g16502 ( 
.A(n_16365),
.Y(n_16502)
);

NAND2xp5_ASAP7_75t_L g16503 ( 
.A(n_16391),
.B(n_2683),
.Y(n_16503)
);

OR2x6_ASAP7_75t_L g16504 ( 
.A(n_16393),
.B(n_2684),
.Y(n_16504)
);

NAND2xp5_ASAP7_75t_L g16505 ( 
.A(n_16404),
.B(n_16405),
.Y(n_16505)
);

AND2x2_ASAP7_75t_L g16506 ( 
.A(n_16329),
.B(n_2684),
.Y(n_16506)
);

INVx1_ASAP7_75t_L g16507 ( 
.A(n_16367),
.Y(n_16507)
);

AND2x2_ASAP7_75t_L g16508 ( 
.A(n_16341),
.B(n_2685),
.Y(n_16508)
);

INVx1_ASAP7_75t_L g16509 ( 
.A(n_16369),
.Y(n_16509)
);

AND2x2_ASAP7_75t_L g16510 ( 
.A(n_16291),
.B(n_2685),
.Y(n_16510)
);

INVx1_ASAP7_75t_L g16511 ( 
.A(n_16328),
.Y(n_16511)
);

INVx2_ASAP7_75t_L g16512 ( 
.A(n_16352),
.Y(n_16512)
);

INVx2_ASAP7_75t_SL g16513 ( 
.A(n_16309),
.Y(n_16513)
);

INVx1_ASAP7_75t_L g16514 ( 
.A(n_16338),
.Y(n_16514)
);

AND2x2_ASAP7_75t_L g16515 ( 
.A(n_16292),
.B(n_2686),
.Y(n_16515)
);

OR2x2_ASAP7_75t_L g16516 ( 
.A(n_16377),
.B(n_2686),
.Y(n_16516)
);

NAND2xp5_ASAP7_75t_L g16517 ( 
.A(n_16300),
.B(n_2687),
.Y(n_16517)
);

INVx1_ASAP7_75t_L g16518 ( 
.A(n_16318),
.Y(n_16518)
);

NOR2xp33_ASAP7_75t_L g16519 ( 
.A(n_16353),
.B(n_2687),
.Y(n_16519)
);

AND2x2_ASAP7_75t_L g16520 ( 
.A(n_16359),
.B(n_16363),
.Y(n_16520)
);

INVx1_ASAP7_75t_L g16521 ( 
.A(n_16337),
.Y(n_16521)
);

INVx1_ASAP7_75t_L g16522 ( 
.A(n_16370),
.Y(n_16522)
);

OR2x2_ASAP7_75t_L g16523 ( 
.A(n_16335),
.B(n_2688),
.Y(n_16523)
);

NAND2xp5_ASAP7_75t_L g16524 ( 
.A(n_16364),
.B(n_16366),
.Y(n_16524)
);

A2O1A1Ixp33_ASAP7_75t_L g16525 ( 
.A1(n_16355),
.A2(n_2690),
.B(n_2688),
.C(n_2689),
.Y(n_16525)
);

INVx1_ASAP7_75t_L g16526 ( 
.A(n_16316),
.Y(n_16526)
);

INVx2_ASAP7_75t_L g16527 ( 
.A(n_16330),
.Y(n_16527)
);

INVx1_ASAP7_75t_SL g16528 ( 
.A(n_16373),
.Y(n_16528)
);

INVx1_ASAP7_75t_L g16529 ( 
.A(n_16331),
.Y(n_16529)
);

AOI22xp5_ASAP7_75t_L g16530 ( 
.A1(n_16378),
.A2(n_2693),
.B1(n_2690),
.B2(n_2691),
.Y(n_16530)
);

INVx1_ASAP7_75t_L g16531 ( 
.A(n_16350),
.Y(n_16531)
);

OR2x2_ASAP7_75t_L g16532 ( 
.A(n_16345),
.B(n_2691),
.Y(n_16532)
);

NOR2xp33_ASAP7_75t_L g16533 ( 
.A(n_16336),
.B(n_2693),
.Y(n_16533)
);

OR2x6_ASAP7_75t_L g16534 ( 
.A(n_16333),
.B(n_2694),
.Y(n_16534)
);

INVx2_ASAP7_75t_SL g16535 ( 
.A(n_16374),
.Y(n_16535)
);

INVx1_ASAP7_75t_L g16536 ( 
.A(n_16368),
.Y(n_16536)
);

INVx1_ASAP7_75t_L g16537 ( 
.A(n_16379),
.Y(n_16537)
);

OAI322xp33_ASAP7_75t_L g16538 ( 
.A1(n_16375),
.A2(n_2699),
.A3(n_2698),
.B1(n_2696),
.B2(n_2694),
.C1(n_2695),
.C2(n_2697),
.Y(n_16538)
);

NAND2xp5_ASAP7_75t_L g16539 ( 
.A(n_16339),
.B(n_2695),
.Y(n_16539)
);

INVx2_ASAP7_75t_L g16540 ( 
.A(n_16381),
.Y(n_16540)
);

INVxp67_ASAP7_75t_L g16541 ( 
.A(n_16376),
.Y(n_16541)
);

AND2x2_ASAP7_75t_L g16542 ( 
.A(n_16274),
.B(n_2696),
.Y(n_16542)
);

OR2x2_ASAP7_75t_L g16543 ( 
.A(n_16321),
.B(n_2698),
.Y(n_16543)
);

NAND2xp5_ASAP7_75t_L g16544 ( 
.A(n_16346),
.B(n_2699),
.Y(n_16544)
);

OAI22xp5_ASAP7_75t_L g16545 ( 
.A1(n_16310),
.A2(n_2702),
.B1(n_2700),
.B2(n_2701),
.Y(n_16545)
);

BUFx2_ASAP7_75t_L g16546 ( 
.A(n_16380),
.Y(n_16546)
);

NAND2xp5_ASAP7_75t_L g16547 ( 
.A(n_16348),
.B(n_2702),
.Y(n_16547)
);

AND2x2_ASAP7_75t_L g16548 ( 
.A(n_16351),
.B(n_2703),
.Y(n_16548)
);

OR2x2_ASAP7_75t_L g16549 ( 
.A(n_16340),
.B(n_2703),
.Y(n_16549)
);

AOI22xp5_ASAP7_75t_L g16550 ( 
.A1(n_16356),
.A2(n_16334),
.B1(n_16371),
.B2(n_2706),
.Y(n_16550)
);

AOI22xp5_ASAP7_75t_L g16551 ( 
.A1(n_16258),
.A2(n_2707),
.B1(n_2704),
.B2(n_2705),
.Y(n_16551)
);

AND2x2_ASAP7_75t_L g16552 ( 
.A(n_16399),
.B(n_2705),
.Y(n_16552)
);

INVx1_ASAP7_75t_L g16553 ( 
.A(n_16402),
.Y(n_16553)
);

OAI211xp5_ASAP7_75t_L g16554 ( 
.A1(n_16260),
.A2(n_2710),
.B(n_2707),
.C(n_2709),
.Y(n_16554)
);

INVx1_ASAP7_75t_L g16555 ( 
.A(n_16414),
.Y(n_16555)
);

OAI22xp5_ASAP7_75t_L g16556 ( 
.A1(n_16416),
.A2(n_2713),
.B1(n_2711),
.B2(n_2712),
.Y(n_16556)
);

NAND4xp25_ASAP7_75t_L g16557 ( 
.A(n_16412),
.B(n_2715),
.C(n_2712),
.D(n_2714),
.Y(n_16557)
);

INVx1_ASAP7_75t_L g16558 ( 
.A(n_16552),
.Y(n_16558)
);

OAI22xp5_ASAP7_75t_L g16559 ( 
.A1(n_16417),
.A2(n_2716),
.B1(n_2714),
.B2(n_2715),
.Y(n_16559)
);

NOR2xp33_ASAP7_75t_L g16560 ( 
.A(n_16422),
.B(n_2716),
.Y(n_16560)
);

HB1xp67_ASAP7_75t_L g16561 ( 
.A(n_16473),
.Y(n_16561)
);

INVx1_ASAP7_75t_L g16562 ( 
.A(n_16429),
.Y(n_16562)
);

OAI32xp33_ASAP7_75t_L g16563 ( 
.A1(n_16410),
.A2(n_2719),
.A3(n_2717),
.B1(n_2718),
.B2(n_2720),
.Y(n_16563)
);

INVx1_ASAP7_75t_L g16564 ( 
.A(n_16413),
.Y(n_16564)
);

INVx2_ASAP7_75t_L g16565 ( 
.A(n_16501),
.Y(n_16565)
);

A2O1A1Ixp33_ASAP7_75t_L g16566 ( 
.A1(n_16553),
.A2(n_16465),
.B(n_16419),
.C(n_16418),
.Y(n_16566)
);

INVx1_ASAP7_75t_SL g16567 ( 
.A(n_16427),
.Y(n_16567)
);

O2A1O1Ixp5_ASAP7_75t_SL g16568 ( 
.A1(n_16451),
.A2(n_2720),
.B(n_2717),
.C(n_2718),
.Y(n_16568)
);

INVx2_ASAP7_75t_SL g16569 ( 
.A(n_16415),
.Y(n_16569)
);

OAI21xp5_ASAP7_75t_L g16570 ( 
.A1(n_16505),
.A2(n_2721),
.B(n_2722),
.Y(n_16570)
);

INVx2_ASAP7_75t_L g16571 ( 
.A(n_16440),
.Y(n_16571)
);

INVx1_ASAP7_75t_L g16572 ( 
.A(n_16433),
.Y(n_16572)
);

INVx1_ASAP7_75t_L g16573 ( 
.A(n_16440),
.Y(n_16573)
);

OAI21xp5_ASAP7_75t_L g16574 ( 
.A1(n_16447),
.A2(n_2721),
.B(n_2722),
.Y(n_16574)
);

AOI22xp5_ASAP7_75t_L g16575 ( 
.A1(n_16411),
.A2(n_2725),
.B1(n_2723),
.B2(n_2724),
.Y(n_16575)
);

NAND2x1p5_ASAP7_75t_L g16576 ( 
.A(n_16463),
.B(n_2723),
.Y(n_16576)
);

OAI22xp5_ASAP7_75t_L g16577 ( 
.A1(n_16484),
.A2(n_2728),
.B1(n_2725),
.B2(n_2727),
.Y(n_16577)
);

INVx2_ASAP7_75t_L g16578 ( 
.A(n_16534),
.Y(n_16578)
);

NAND2x1p5_ASAP7_75t_L g16579 ( 
.A(n_16478),
.B(n_2727),
.Y(n_16579)
);

NAND2xp5_ASAP7_75t_L g16580 ( 
.A(n_16464),
.B(n_2729),
.Y(n_16580)
);

INVxp67_ASAP7_75t_L g16581 ( 
.A(n_16519),
.Y(n_16581)
);

INVx1_ASAP7_75t_L g16582 ( 
.A(n_16441),
.Y(n_16582)
);

INVx1_ASAP7_75t_L g16583 ( 
.A(n_16485),
.Y(n_16583)
);

AND2x2_ASAP7_75t_L g16584 ( 
.A(n_16426),
.B(n_2729),
.Y(n_16584)
);

NAND2xp5_ASAP7_75t_L g16585 ( 
.A(n_16436),
.B(n_2730),
.Y(n_16585)
);

AND2x2_ASAP7_75t_L g16586 ( 
.A(n_16481),
.B(n_2730),
.Y(n_16586)
);

INVx2_ASAP7_75t_L g16587 ( 
.A(n_16534),
.Y(n_16587)
);

NOR2xp67_ASAP7_75t_L g16588 ( 
.A(n_16462),
.B(n_2731),
.Y(n_16588)
);

INVx1_ASAP7_75t_L g16589 ( 
.A(n_16477),
.Y(n_16589)
);

INVx1_ASAP7_75t_L g16590 ( 
.A(n_16449),
.Y(n_16590)
);

INVx2_ASAP7_75t_L g16591 ( 
.A(n_16504),
.Y(n_16591)
);

AOI22xp33_ASAP7_75t_SL g16592 ( 
.A1(n_16546),
.A2(n_2734),
.B1(n_2732),
.B2(n_2733),
.Y(n_16592)
);

NAND2xp5_ASAP7_75t_L g16593 ( 
.A(n_16420),
.B(n_2732),
.Y(n_16593)
);

OAI21xp5_ASAP7_75t_L g16594 ( 
.A1(n_16445),
.A2(n_2733),
.B(n_2734),
.Y(n_16594)
);

INVx1_ASAP7_75t_L g16595 ( 
.A(n_16455),
.Y(n_16595)
);

INVx1_ASAP7_75t_L g16596 ( 
.A(n_16424),
.Y(n_16596)
);

OR2x2_ASAP7_75t_L g16597 ( 
.A(n_16481),
.B(n_2735),
.Y(n_16597)
);

OR2x2_ASAP7_75t_L g16598 ( 
.A(n_16484),
.B(n_2735),
.Y(n_16598)
);

INVx1_ASAP7_75t_L g16599 ( 
.A(n_16482),
.Y(n_16599)
);

INVx1_ASAP7_75t_SL g16600 ( 
.A(n_16472),
.Y(n_16600)
);

INVx1_ASAP7_75t_SL g16601 ( 
.A(n_16516),
.Y(n_16601)
);

AOI22xp5_ASAP7_75t_L g16602 ( 
.A1(n_16540),
.A2(n_2738),
.B1(n_2736),
.B2(n_2737),
.Y(n_16602)
);

INVx1_ASAP7_75t_L g16603 ( 
.A(n_16431),
.Y(n_16603)
);

INVx4_ASAP7_75t_L g16604 ( 
.A(n_16458),
.Y(n_16604)
);

AND2x2_ASAP7_75t_L g16605 ( 
.A(n_16421),
.B(n_2737),
.Y(n_16605)
);

INVx1_ASAP7_75t_L g16606 ( 
.A(n_16476),
.Y(n_16606)
);

AOI22xp5_ASAP7_75t_L g16607 ( 
.A1(n_16428),
.A2(n_2740),
.B1(n_2738),
.B2(n_2739),
.Y(n_16607)
);

AOI222xp33_ASAP7_75t_L g16608 ( 
.A1(n_16537),
.A2(n_2742),
.B1(n_2744),
.B2(n_2740),
.C1(n_2741),
.C2(n_2743),
.Y(n_16608)
);

NAND2xp5_ASAP7_75t_L g16609 ( 
.A(n_16430),
.B(n_2741),
.Y(n_16609)
);

INVx1_ASAP7_75t_L g16610 ( 
.A(n_16425),
.Y(n_16610)
);

INVx1_ASAP7_75t_L g16611 ( 
.A(n_16504),
.Y(n_16611)
);

AND2x2_ASAP7_75t_L g16612 ( 
.A(n_16520),
.B(n_2742),
.Y(n_16612)
);

INVx1_ASAP7_75t_L g16613 ( 
.A(n_16510),
.Y(n_16613)
);

NAND2xp5_ASAP7_75t_L g16614 ( 
.A(n_16467),
.B(n_2743),
.Y(n_16614)
);

NAND2xp5_ASAP7_75t_L g16615 ( 
.A(n_16470),
.B(n_2744),
.Y(n_16615)
);

NAND2xp5_ASAP7_75t_L g16616 ( 
.A(n_16515),
.B(n_2745),
.Y(n_16616)
);

INVx1_ASAP7_75t_L g16617 ( 
.A(n_16493),
.Y(n_16617)
);

OAI21xp33_ASAP7_75t_L g16618 ( 
.A1(n_16524),
.A2(n_2745),
.B(n_2746),
.Y(n_16618)
);

AND2x2_ASAP7_75t_L g16619 ( 
.A(n_16487),
.B(n_2746),
.Y(n_16619)
);

INVxp67_ASAP7_75t_SL g16620 ( 
.A(n_16474),
.Y(n_16620)
);

NAND2x1_ASAP7_75t_L g16621 ( 
.A(n_16444),
.B(n_2747),
.Y(n_16621)
);

INVx1_ASAP7_75t_SL g16622 ( 
.A(n_16434),
.Y(n_16622)
);

AND2x2_ASAP7_75t_L g16623 ( 
.A(n_16450),
.B(n_2747),
.Y(n_16623)
);

AOI21xp5_ASAP7_75t_L g16624 ( 
.A1(n_16432),
.A2(n_2748),
.B(n_2749),
.Y(n_16624)
);

INVx1_ASAP7_75t_L g16625 ( 
.A(n_16506),
.Y(n_16625)
);

INVx1_ASAP7_75t_L g16626 ( 
.A(n_16457),
.Y(n_16626)
);

NAND2xp5_ASAP7_75t_L g16627 ( 
.A(n_16486),
.B(n_2748),
.Y(n_16627)
);

INVx1_ASAP7_75t_L g16628 ( 
.A(n_16508),
.Y(n_16628)
);

XOR2x2_ASAP7_75t_L g16629 ( 
.A(n_16480),
.B(n_2749),
.Y(n_16629)
);

OR2x2_ASAP7_75t_L g16630 ( 
.A(n_16498),
.B(n_2750),
.Y(n_16630)
);

AND2x2_ASAP7_75t_L g16631 ( 
.A(n_16437),
.B(n_2750),
.Y(n_16631)
);

INVx2_ASAP7_75t_L g16632 ( 
.A(n_16543),
.Y(n_16632)
);

XNOR2xp5_ASAP7_75t_L g16633 ( 
.A(n_16528),
.B(n_2751),
.Y(n_16633)
);

INVx2_ASAP7_75t_SL g16634 ( 
.A(n_16513),
.Y(n_16634)
);

AND2x2_ASAP7_75t_L g16635 ( 
.A(n_16502),
.B(n_2751),
.Y(n_16635)
);

INVx2_ASAP7_75t_L g16636 ( 
.A(n_16549),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_16452),
.Y(n_16637)
);

NAND2x1p5_ASAP7_75t_L g16638 ( 
.A(n_16535),
.B(n_2752),
.Y(n_16638)
);

INVx1_ASAP7_75t_L g16639 ( 
.A(n_16496),
.Y(n_16639)
);

OR2x2_ASAP7_75t_L g16640 ( 
.A(n_16523),
.B(n_2752),
.Y(n_16640)
);

OAI32xp33_ASAP7_75t_L g16641 ( 
.A1(n_16503),
.A2(n_2755),
.A3(n_2753),
.B1(n_2754),
.B2(n_2756),
.Y(n_16641)
);

INVx1_ASAP7_75t_L g16642 ( 
.A(n_16468),
.Y(n_16642)
);

NAND2xp5_ASAP7_75t_L g16643 ( 
.A(n_16507),
.B(n_2754),
.Y(n_16643)
);

OR2x2_ASAP7_75t_L g16644 ( 
.A(n_16495),
.B(n_2755),
.Y(n_16644)
);

INVx1_ASAP7_75t_L g16645 ( 
.A(n_16542),
.Y(n_16645)
);

INVx1_ASAP7_75t_L g16646 ( 
.A(n_16456),
.Y(n_16646)
);

INVx1_ASAP7_75t_L g16647 ( 
.A(n_16517),
.Y(n_16647)
);

AND2x2_ASAP7_75t_L g16648 ( 
.A(n_16466),
.B(n_2756),
.Y(n_16648)
);

INVx2_ASAP7_75t_SL g16649 ( 
.A(n_16512),
.Y(n_16649)
);

INVx1_ASAP7_75t_SL g16650 ( 
.A(n_16439),
.Y(n_16650)
);

AOI21xp5_ASAP7_75t_L g16651 ( 
.A1(n_16423),
.A2(n_2757),
.B(n_2758),
.Y(n_16651)
);

NAND2xp5_ASAP7_75t_L g16652 ( 
.A(n_16460),
.B(n_16469),
.Y(n_16652)
);

OR2x2_ASAP7_75t_L g16653 ( 
.A(n_16442),
.B(n_2759),
.Y(n_16653)
);

INVx1_ASAP7_75t_L g16654 ( 
.A(n_16548),
.Y(n_16654)
);

INVx1_ASAP7_75t_L g16655 ( 
.A(n_16539),
.Y(n_16655)
);

AOI21xp33_ASAP7_75t_L g16656 ( 
.A1(n_16475),
.A2(n_2759),
.B(n_2760),
.Y(n_16656)
);

INVxp67_ASAP7_75t_L g16657 ( 
.A(n_16533),
.Y(n_16657)
);

AOI22xp5_ASAP7_75t_L g16658 ( 
.A1(n_16471),
.A2(n_2762),
.B1(n_2760),
.B2(n_2761),
.Y(n_16658)
);

NAND2xp5_ASAP7_75t_L g16659 ( 
.A(n_16479),
.B(n_2761),
.Y(n_16659)
);

NAND4xp75_ASAP7_75t_SL g16660 ( 
.A(n_16483),
.B(n_2764),
.C(n_2762),
.D(n_2763),
.Y(n_16660)
);

HB1xp67_ASAP7_75t_L g16661 ( 
.A(n_16499),
.Y(n_16661)
);

AOI22xp33_ASAP7_75t_L g16662 ( 
.A1(n_16489),
.A2(n_2767),
.B1(n_2765),
.B2(n_2766),
.Y(n_16662)
);

OAI22xp5_ASAP7_75t_L g16663 ( 
.A1(n_16491),
.A2(n_16497),
.B1(n_16492),
.B2(n_16509),
.Y(n_16663)
);

INVx1_ASAP7_75t_SL g16664 ( 
.A(n_16532),
.Y(n_16664)
);

NAND2xp5_ASAP7_75t_L g16665 ( 
.A(n_16453),
.B(n_2765),
.Y(n_16665)
);

AOI22xp33_ASAP7_75t_SL g16666 ( 
.A1(n_16435),
.A2(n_2769),
.B1(n_2767),
.B2(n_2768),
.Y(n_16666)
);

OAI22xp5_ASAP7_75t_L g16667 ( 
.A1(n_16550),
.A2(n_2771),
.B1(n_2768),
.B2(n_2769),
.Y(n_16667)
);

INVx2_ASAP7_75t_L g16668 ( 
.A(n_16454),
.Y(n_16668)
);

OR2x2_ASAP7_75t_L g16669 ( 
.A(n_16500),
.B(n_2771),
.Y(n_16669)
);

AND2x2_ASAP7_75t_L g16670 ( 
.A(n_16522),
.B(n_2772),
.Y(n_16670)
);

NAND2xp5_ASAP7_75t_L g16671 ( 
.A(n_16551),
.B(n_2772),
.Y(n_16671)
);

AOI22xp5_ASAP7_75t_L g16672 ( 
.A1(n_16541),
.A2(n_2775),
.B1(n_2773),
.B2(n_2774),
.Y(n_16672)
);

AOI21xp33_ASAP7_75t_SL g16673 ( 
.A1(n_16446),
.A2(n_2773),
.B(n_2774),
.Y(n_16673)
);

NAND2xp5_ASAP7_75t_L g16674 ( 
.A(n_16459),
.B(n_2775),
.Y(n_16674)
);

OAI31xp33_ASAP7_75t_L g16675 ( 
.A1(n_16554),
.A2(n_2778),
.A3(n_2776),
.B(n_2777),
.Y(n_16675)
);

AOI31xp33_ASAP7_75t_L g16676 ( 
.A1(n_16461),
.A2(n_2779),
.A3(n_2777),
.B(n_2778),
.Y(n_16676)
);

INVx1_ASAP7_75t_L g16677 ( 
.A(n_16488),
.Y(n_16677)
);

AND2x4_ASAP7_75t_L g16678 ( 
.A(n_16527),
.B(n_2779),
.Y(n_16678)
);

AOI22xp5_ASAP7_75t_L g16679 ( 
.A1(n_16438),
.A2(n_2782),
.B1(n_2780),
.B2(n_2781),
.Y(n_16679)
);

INVx1_ASAP7_75t_L g16680 ( 
.A(n_16544),
.Y(n_16680)
);

INVxp67_ASAP7_75t_L g16681 ( 
.A(n_16547),
.Y(n_16681)
);

NOR2xp33_ASAP7_75t_L g16682 ( 
.A(n_16490),
.B(n_2780),
.Y(n_16682)
);

OR2x2_ASAP7_75t_L g16683 ( 
.A(n_16511),
.B(n_2781),
.Y(n_16683)
);

INVx2_ASAP7_75t_L g16684 ( 
.A(n_16443),
.Y(n_16684)
);

OR2x2_ASAP7_75t_L g16685 ( 
.A(n_16494),
.B(n_2783),
.Y(n_16685)
);

NAND2xp5_ASAP7_75t_SL g16686 ( 
.A(n_16530),
.B(n_2784),
.Y(n_16686)
);

OAI22xp5_ASAP7_75t_L g16687 ( 
.A1(n_16448),
.A2(n_2788),
.B1(n_2785),
.B2(n_2786),
.Y(n_16687)
);

INVx2_ASAP7_75t_L g16688 ( 
.A(n_16514),
.Y(n_16688)
);

INVx1_ASAP7_75t_L g16689 ( 
.A(n_16525),
.Y(n_16689)
);

NAND2xp5_ASAP7_75t_L g16690 ( 
.A(n_16521),
.B(n_2786),
.Y(n_16690)
);

OAI22xp5_ASAP7_75t_L g16691 ( 
.A1(n_16567),
.A2(n_16562),
.B1(n_16622),
.B2(n_16564),
.Y(n_16691)
);

INVx2_ASAP7_75t_L g16692 ( 
.A(n_16597),
.Y(n_16692)
);

NAND4xp25_ASAP7_75t_L g16693 ( 
.A(n_16566),
.B(n_16536),
.C(n_16518),
.D(n_16529),
.Y(n_16693)
);

AOI22xp33_ASAP7_75t_SL g16694 ( 
.A1(n_16604),
.A2(n_16526),
.B1(n_16531),
.B2(n_16545),
.Y(n_16694)
);

INVx2_ASAP7_75t_SL g16695 ( 
.A(n_16598),
.Y(n_16695)
);

INVx1_ASAP7_75t_L g16696 ( 
.A(n_16586),
.Y(n_16696)
);

INVx1_ASAP7_75t_SL g16697 ( 
.A(n_16660),
.Y(n_16697)
);

OR2x2_ASAP7_75t_L g16698 ( 
.A(n_16555),
.B(n_16638),
.Y(n_16698)
);

AND2x4_ASAP7_75t_L g16699 ( 
.A(n_16588),
.B(n_16538),
.Y(n_16699)
);

INVx1_ASAP7_75t_L g16700 ( 
.A(n_16576),
.Y(n_16700)
);

NAND2xp5_ASAP7_75t_L g16701 ( 
.A(n_16612),
.B(n_2788),
.Y(n_16701)
);

INVx1_ASAP7_75t_L g16702 ( 
.A(n_16579),
.Y(n_16702)
);

NAND2xp5_ASAP7_75t_L g16703 ( 
.A(n_16605),
.B(n_2789),
.Y(n_16703)
);

INVx1_ASAP7_75t_L g16704 ( 
.A(n_16633),
.Y(n_16704)
);

OAI22xp33_ASAP7_75t_L g16705 ( 
.A1(n_16649),
.A2(n_2791),
.B1(n_2789),
.B2(n_2790),
.Y(n_16705)
);

INVx1_ASAP7_75t_L g16706 ( 
.A(n_16561),
.Y(n_16706)
);

AND2x2_ASAP7_75t_L g16707 ( 
.A(n_16569),
.B(n_2791),
.Y(n_16707)
);

AOI221x1_ASAP7_75t_L g16708 ( 
.A1(n_16663),
.A2(n_2794),
.B1(n_2792),
.B2(n_2793),
.C(n_2795),
.Y(n_16708)
);

INVx2_ASAP7_75t_SL g16709 ( 
.A(n_16621),
.Y(n_16709)
);

OAI21xp33_ASAP7_75t_L g16710 ( 
.A1(n_16634),
.A2(n_2793),
.B(n_2794),
.Y(n_16710)
);

INVx1_ASAP7_75t_L g16711 ( 
.A(n_16661),
.Y(n_16711)
);

INVx1_ASAP7_75t_L g16712 ( 
.A(n_16623),
.Y(n_16712)
);

OAI21xp33_ASAP7_75t_SL g16713 ( 
.A1(n_16573),
.A2(n_2795),
.B(n_2796),
.Y(n_16713)
);

NAND3xp33_ASAP7_75t_L g16714 ( 
.A(n_16675),
.B(n_2796),
.C(n_2797),
.Y(n_16714)
);

NAND2xp5_ASAP7_75t_L g16715 ( 
.A(n_16635),
.B(n_2797),
.Y(n_16715)
);

NAND2xp5_ASAP7_75t_L g16716 ( 
.A(n_16678),
.B(n_2798),
.Y(n_16716)
);

INVx2_ASAP7_75t_L g16717 ( 
.A(n_16678),
.Y(n_16717)
);

INVx1_ASAP7_75t_L g16718 ( 
.A(n_16619),
.Y(n_16718)
);

INVx1_ASAP7_75t_SL g16719 ( 
.A(n_16670),
.Y(n_16719)
);

INVx1_ASAP7_75t_L g16720 ( 
.A(n_16644),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_16631),
.Y(n_16721)
);

OR2x2_ASAP7_75t_L g16722 ( 
.A(n_16571),
.B(n_2798),
.Y(n_16722)
);

INVx2_ASAP7_75t_SL g16723 ( 
.A(n_16578),
.Y(n_16723)
);

AND2x2_ASAP7_75t_L g16724 ( 
.A(n_16565),
.B(n_2799),
.Y(n_16724)
);

AND2x2_ASAP7_75t_L g16725 ( 
.A(n_16582),
.B(n_2800),
.Y(n_16725)
);

OAI22xp33_ASAP7_75t_SL g16726 ( 
.A1(n_16685),
.A2(n_16611),
.B1(n_16677),
.B2(n_16558),
.Y(n_16726)
);

INVx1_ASAP7_75t_L g16727 ( 
.A(n_16630),
.Y(n_16727)
);

INVxp67_ASAP7_75t_L g16728 ( 
.A(n_16560),
.Y(n_16728)
);

INVx3_ASAP7_75t_L g16729 ( 
.A(n_16591),
.Y(n_16729)
);

OR2x2_ASAP7_75t_L g16730 ( 
.A(n_16587),
.B(n_2800),
.Y(n_16730)
);

NOR2xp33_ASAP7_75t_L g16731 ( 
.A(n_16557),
.B(n_2802),
.Y(n_16731)
);

AND2x2_ASAP7_75t_L g16732 ( 
.A(n_16583),
.B(n_2802),
.Y(n_16732)
);

INVx1_ASAP7_75t_L g16733 ( 
.A(n_16648),
.Y(n_16733)
);

AOI211xp5_ASAP7_75t_L g16734 ( 
.A1(n_16673),
.A2(n_2805),
.B(n_2803),
.C(n_2804),
.Y(n_16734)
);

NOR2xp33_ASAP7_75t_SL g16735 ( 
.A(n_16600),
.B(n_2803),
.Y(n_16735)
);

NAND2xp5_ASAP7_75t_L g16736 ( 
.A(n_16592),
.B(n_2805),
.Y(n_16736)
);

INVx2_ASAP7_75t_L g16737 ( 
.A(n_16669),
.Y(n_16737)
);

INVx1_ASAP7_75t_L g16738 ( 
.A(n_16683),
.Y(n_16738)
);

INVx1_ASAP7_75t_SL g16739 ( 
.A(n_16640),
.Y(n_16739)
);

OAI22xp5_ASAP7_75t_L g16740 ( 
.A1(n_16668),
.A2(n_2808),
.B1(n_2806),
.B2(n_2807),
.Y(n_16740)
);

NOR2xp67_ASAP7_75t_L g16741 ( 
.A(n_16572),
.B(n_2806),
.Y(n_16741)
);

NAND2xp5_ASAP7_75t_SL g16742 ( 
.A(n_16594),
.B(n_2807),
.Y(n_16742)
);

INVx1_ASAP7_75t_L g16743 ( 
.A(n_16584),
.Y(n_16743)
);

INVx2_ASAP7_75t_L g16744 ( 
.A(n_16653),
.Y(n_16744)
);

AND2x2_ASAP7_75t_L g16745 ( 
.A(n_16599),
.B(n_2809),
.Y(n_16745)
);

AOI221xp5_ASAP7_75t_L g16746 ( 
.A1(n_16689),
.A2(n_2811),
.B1(n_2809),
.B2(n_2810),
.C(n_2812),
.Y(n_16746)
);

INVx1_ASAP7_75t_L g16747 ( 
.A(n_16676),
.Y(n_16747)
);

NAND2xp5_ASAP7_75t_L g16748 ( 
.A(n_16666),
.B(n_2810),
.Y(n_16748)
);

AOI31xp33_ASAP7_75t_L g16749 ( 
.A1(n_16601),
.A2(n_16625),
.A3(n_16617),
.B(n_16652),
.Y(n_16749)
);

INVx1_ASAP7_75t_SL g16750 ( 
.A(n_16629),
.Y(n_16750)
);

AND2x4_ASAP7_75t_L g16751 ( 
.A(n_16589),
.B(n_2811),
.Y(n_16751)
);

AOI22xp5_ASAP7_75t_L g16752 ( 
.A1(n_16613),
.A2(n_2814),
.B1(n_2812),
.B2(n_2813),
.Y(n_16752)
);

INVx1_ASAP7_75t_L g16753 ( 
.A(n_16580),
.Y(n_16753)
);

INVxp33_ASAP7_75t_L g16754 ( 
.A(n_16682),
.Y(n_16754)
);

OAI211xp5_ASAP7_75t_L g16755 ( 
.A1(n_16593),
.A2(n_16609),
.B(n_16643),
.C(n_16665),
.Y(n_16755)
);

INVxp67_ASAP7_75t_L g16756 ( 
.A(n_16585),
.Y(n_16756)
);

AND2x2_ASAP7_75t_L g16757 ( 
.A(n_16645),
.B(n_2813),
.Y(n_16757)
);

INVxp67_ASAP7_75t_L g16758 ( 
.A(n_16616),
.Y(n_16758)
);

AND2x2_ASAP7_75t_L g16759 ( 
.A(n_16654),
.B(n_2814),
.Y(n_16759)
);

AND2x2_ASAP7_75t_L g16760 ( 
.A(n_16606),
.B(n_2815),
.Y(n_16760)
);

NAND2xp5_ASAP7_75t_L g16761 ( 
.A(n_16575),
.B(n_2815),
.Y(n_16761)
);

OAI22xp5_ASAP7_75t_SL g16762 ( 
.A1(n_16628),
.A2(n_2818),
.B1(n_2816),
.B2(n_2817),
.Y(n_16762)
);

NAND2xp5_ASAP7_75t_L g16763 ( 
.A(n_16608),
.B(n_2816),
.Y(n_16763)
);

AOI21xp33_ASAP7_75t_L g16764 ( 
.A1(n_16614),
.A2(n_2817),
.B(n_2818),
.Y(n_16764)
);

INVxp67_ASAP7_75t_L g16765 ( 
.A(n_16615),
.Y(n_16765)
);

INVx1_ASAP7_75t_L g16766 ( 
.A(n_16627),
.Y(n_16766)
);

AND2x2_ASAP7_75t_L g16767 ( 
.A(n_16590),
.B(n_2819),
.Y(n_16767)
);

INVx1_ASAP7_75t_L g16768 ( 
.A(n_16659),
.Y(n_16768)
);

INVx1_ASAP7_75t_L g16769 ( 
.A(n_16674),
.Y(n_16769)
);

INVx1_ASAP7_75t_L g16770 ( 
.A(n_16671),
.Y(n_16770)
);

AOI21xp5_ASAP7_75t_L g16771 ( 
.A1(n_16651),
.A2(n_2819),
.B(n_2820),
.Y(n_16771)
);

INVx1_ASAP7_75t_L g16772 ( 
.A(n_16556),
.Y(n_16772)
);

INVxp67_ASAP7_75t_L g16773 ( 
.A(n_16577),
.Y(n_16773)
);

INVx1_ASAP7_75t_L g16774 ( 
.A(n_16690),
.Y(n_16774)
);

NOR2xp33_ASAP7_75t_L g16775 ( 
.A(n_16618),
.B(n_2821),
.Y(n_16775)
);

INVxp67_ASAP7_75t_L g16776 ( 
.A(n_16559),
.Y(n_16776)
);

OAI21xp33_ASAP7_75t_SL g16777 ( 
.A1(n_16568),
.A2(n_2821),
.B(n_2822),
.Y(n_16777)
);

NAND2xp5_ASAP7_75t_L g16778 ( 
.A(n_16595),
.B(n_2822),
.Y(n_16778)
);

OAI22xp5_ASAP7_75t_L g16779 ( 
.A1(n_16581),
.A2(n_2825),
.B1(n_2823),
.B2(n_2824),
.Y(n_16779)
);

AOI22xp5_ASAP7_75t_L g16780 ( 
.A1(n_16650),
.A2(n_2825),
.B1(n_2823),
.B2(n_2824),
.Y(n_16780)
);

INVx1_ASAP7_75t_L g16781 ( 
.A(n_16632),
.Y(n_16781)
);

OR2x2_ASAP7_75t_L g16782 ( 
.A(n_16636),
.B(n_2826),
.Y(n_16782)
);

NAND2xp5_ASAP7_75t_L g16783 ( 
.A(n_16662),
.B(n_2826),
.Y(n_16783)
);

AO21x1_ASAP7_75t_L g16784 ( 
.A1(n_16686),
.A2(n_2827),
.B(n_2828),
.Y(n_16784)
);

AOI21xp5_ASAP7_75t_L g16785 ( 
.A1(n_16624),
.A2(n_2827),
.B(n_2828),
.Y(n_16785)
);

INVx2_ASAP7_75t_L g16786 ( 
.A(n_16626),
.Y(n_16786)
);

INVx1_ASAP7_75t_L g16787 ( 
.A(n_16574),
.Y(n_16787)
);

NAND2xp5_ASAP7_75t_L g16788 ( 
.A(n_16607),
.B(n_2829),
.Y(n_16788)
);

INVx1_ASAP7_75t_L g16789 ( 
.A(n_16667),
.Y(n_16789)
);

AND2x2_ASAP7_75t_L g16790 ( 
.A(n_16664),
.B(n_2829),
.Y(n_16790)
);

NAND2xp5_ASAP7_75t_L g16791 ( 
.A(n_16672),
.B(n_2830),
.Y(n_16791)
);

INVx1_ASAP7_75t_L g16792 ( 
.A(n_16570),
.Y(n_16792)
);

NAND5xp2_ASAP7_75t_L g16793 ( 
.A(n_16610),
.B(n_2832),
.C(n_2830),
.D(n_2831),
.E(n_2833),
.Y(n_16793)
);

NAND2xp5_ASAP7_75t_L g16794 ( 
.A(n_16596),
.B(n_2831),
.Y(n_16794)
);

AOI222xp33_ASAP7_75t_L g16795 ( 
.A1(n_16657),
.A2(n_2835),
.B1(n_2837),
.B2(n_2832),
.C1(n_2834),
.C2(n_2836),
.Y(n_16795)
);

OAI21xp33_ASAP7_75t_L g16796 ( 
.A1(n_16639),
.A2(n_16603),
.B(n_16620),
.Y(n_16796)
);

INVx2_ASAP7_75t_L g16797 ( 
.A(n_16637),
.Y(n_16797)
);

NAND3xp33_ASAP7_75t_L g16798 ( 
.A(n_16688),
.B(n_2835),
.C(n_2837),
.Y(n_16798)
);

O2A1O1Ixp33_ASAP7_75t_SL g16799 ( 
.A1(n_16563),
.A2(n_2840),
.B(n_2838),
.C(n_2839),
.Y(n_16799)
);

AOI322xp5_ASAP7_75t_L g16800 ( 
.A1(n_16642),
.A2(n_2844),
.A3(n_2843),
.B1(n_2841),
.B2(n_2838),
.C1(n_2839),
.C2(n_2842),
.Y(n_16800)
);

INVx1_ASAP7_75t_L g16801 ( 
.A(n_16687),
.Y(n_16801)
);

AND2x2_ASAP7_75t_L g16802 ( 
.A(n_16684),
.B(n_2841),
.Y(n_16802)
);

OAI211xp5_ASAP7_75t_L g16803 ( 
.A1(n_16656),
.A2(n_2847),
.B(n_2842),
.C(n_2845),
.Y(n_16803)
);

OAI31xp33_ASAP7_75t_L g16804 ( 
.A1(n_16646),
.A2(n_2849),
.A3(n_2845),
.B(n_2848),
.Y(n_16804)
);

OR2x2_ASAP7_75t_L g16805 ( 
.A(n_16655),
.B(n_2848),
.Y(n_16805)
);

AND2x2_ASAP7_75t_L g16806 ( 
.A(n_16647),
.B(n_2849),
.Y(n_16806)
);

NOR2xp33_ASAP7_75t_SL g16807 ( 
.A(n_16641),
.B(n_2850),
.Y(n_16807)
);

OAI22xp5_ASAP7_75t_L g16808 ( 
.A1(n_16681),
.A2(n_2852),
.B1(n_2850),
.B2(n_2851),
.Y(n_16808)
);

OAI22xp5_ASAP7_75t_L g16809 ( 
.A1(n_16680),
.A2(n_2854),
.B1(n_2852),
.B2(n_2853),
.Y(n_16809)
);

INVx2_ASAP7_75t_L g16810 ( 
.A(n_16658),
.Y(n_16810)
);

AOI22xp5_ASAP7_75t_L g16811 ( 
.A1(n_16602),
.A2(n_2855),
.B1(n_2853),
.B2(n_2854),
.Y(n_16811)
);

INVx1_ASAP7_75t_L g16812 ( 
.A(n_16679),
.Y(n_16812)
);

CKINVDCx14_ASAP7_75t_R g16813 ( 
.A(n_16555),
.Y(n_16813)
);

INVxp67_ASAP7_75t_L g16814 ( 
.A(n_16555),
.Y(n_16814)
);

OAI32xp33_ASAP7_75t_L g16815 ( 
.A1(n_16567),
.A2(n_2857),
.A3(n_2855),
.B1(n_2856),
.B2(n_2858),
.Y(n_16815)
);

OR2x2_ASAP7_75t_L g16816 ( 
.A(n_16555),
.B(n_2856),
.Y(n_16816)
);

BUFx2_ASAP7_75t_L g16817 ( 
.A(n_16555),
.Y(n_16817)
);

OAI222xp33_ASAP7_75t_L g16818 ( 
.A1(n_16697),
.A2(n_16814),
.B1(n_16711),
.B2(n_16691),
.C1(n_16709),
.C2(n_16813),
.Y(n_16818)
);

OAI21xp33_ASAP7_75t_L g16819 ( 
.A1(n_16807),
.A2(n_2857),
.B(n_2858),
.Y(n_16819)
);

AOI21xp5_ASAP7_75t_L g16820 ( 
.A1(n_16742),
.A2(n_2859),
.B(n_2860),
.Y(n_16820)
);

INVx1_ASAP7_75t_L g16821 ( 
.A(n_16816),
.Y(n_16821)
);

INVx2_ASAP7_75t_L g16822 ( 
.A(n_16751),
.Y(n_16822)
);

AOI21xp33_ASAP7_75t_SL g16823 ( 
.A1(n_16698),
.A2(n_2860),
.B(n_2861),
.Y(n_16823)
);

OA21x2_ASAP7_75t_L g16824 ( 
.A1(n_16817),
.A2(n_2861),
.B(n_2862),
.Y(n_16824)
);

AOI21x1_ASAP7_75t_L g16825 ( 
.A1(n_16741),
.A2(n_2862),
.B(n_2863),
.Y(n_16825)
);

OAI221xp5_ASAP7_75t_L g16826 ( 
.A1(n_16713),
.A2(n_2865),
.B1(n_2863),
.B2(n_2864),
.C(n_2866),
.Y(n_16826)
);

OAI221xp5_ASAP7_75t_L g16827 ( 
.A1(n_16694),
.A2(n_2866),
.B1(n_2864),
.B2(n_2865),
.C(n_2867),
.Y(n_16827)
);

A2O1A1Ixp33_ASAP7_75t_L g16828 ( 
.A1(n_16777),
.A2(n_16804),
.B(n_16731),
.C(n_16775),
.Y(n_16828)
);

AOI22xp33_ASAP7_75t_L g16829 ( 
.A1(n_16729),
.A2(n_2869),
.B1(n_2867),
.B2(n_2868),
.Y(n_16829)
);

OAI21xp5_ASAP7_75t_L g16830 ( 
.A1(n_16714),
.A2(n_2868),
.B(n_2869),
.Y(n_16830)
);

OAI21xp33_ASAP7_75t_L g16831 ( 
.A1(n_16723),
.A2(n_2870),
.B(n_2871),
.Y(n_16831)
);

INVx1_ASAP7_75t_L g16832 ( 
.A(n_16725),
.Y(n_16832)
);

OAI22xp5_ASAP7_75t_L g16833 ( 
.A1(n_16706),
.A2(n_2872),
.B1(n_2870),
.B2(n_2871),
.Y(n_16833)
);

AOI22xp33_ASAP7_75t_L g16834 ( 
.A1(n_16699),
.A2(n_2874),
.B1(n_2872),
.B2(n_2873),
.Y(n_16834)
);

AOI22xp5_ASAP7_75t_L g16835 ( 
.A1(n_16699),
.A2(n_2876),
.B1(n_2874),
.B2(n_2875),
.Y(n_16835)
);

INVx1_ASAP7_75t_L g16836 ( 
.A(n_16732),
.Y(n_16836)
);

OAI21xp33_ASAP7_75t_L g16837 ( 
.A1(n_16749),
.A2(n_2875),
.B(n_2877),
.Y(n_16837)
);

OAI21xp5_ASAP7_75t_SL g16838 ( 
.A1(n_16773),
.A2(n_2878),
.B(n_2879),
.Y(n_16838)
);

OAI322xp33_ASAP7_75t_L g16839 ( 
.A1(n_16776),
.A2(n_16750),
.A3(n_16747),
.B1(n_16781),
.B2(n_16772),
.C1(n_16719),
.C2(n_16704),
.Y(n_16839)
);

OAI21xp5_ASAP7_75t_L g16840 ( 
.A1(n_16785),
.A2(n_2878),
.B(n_2879),
.Y(n_16840)
);

O2A1O1Ixp33_ASAP7_75t_L g16841 ( 
.A1(n_16799),
.A2(n_16726),
.B(n_16702),
.C(n_16700),
.Y(n_16841)
);

OAI22xp5_ASAP7_75t_L g16842 ( 
.A1(n_16811),
.A2(n_2882),
.B1(n_2880),
.B2(n_2881),
.Y(n_16842)
);

AOI31xp33_ASAP7_75t_L g16843 ( 
.A1(n_16784),
.A2(n_16734),
.A3(n_16754),
.B(n_16763),
.Y(n_16843)
);

XOR2x2_ASAP7_75t_L g16844 ( 
.A(n_16798),
.B(n_2880),
.Y(n_16844)
);

AOI211xp5_ASAP7_75t_L g16845 ( 
.A1(n_16803),
.A2(n_2884),
.B(n_2882),
.C(n_2883),
.Y(n_16845)
);

A2O1A1Ixp33_ASAP7_75t_L g16846 ( 
.A1(n_16710),
.A2(n_2885),
.B(n_2883),
.C(n_2884),
.Y(n_16846)
);

OAI22xp5_ASAP7_75t_L g16847 ( 
.A1(n_16786),
.A2(n_2887),
.B1(n_2885),
.B2(n_2886),
.Y(n_16847)
);

AND2x2_ASAP7_75t_L g16848 ( 
.A(n_16707),
.B(n_16790),
.Y(n_16848)
);

AOI21xp5_ASAP7_75t_L g16849 ( 
.A1(n_16716),
.A2(n_2886),
.B(n_2887),
.Y(n_16849)
);

INVx1_ASAP7_75t_L g16850 ( 
.A(n_16751),
.Y(n_16850)
);

INVx2_ASAP7_75t_SL g16851 ( 
.A(n_16717),
.Y(n_16851)
);

A2O1A1Ixp33_ASAP7_75t_L g16852 ( 
.A1(n_16771),
.A2(n_2890),
.B(n_2888),
.C(n_2889),
.Y(n_16852)
);

NAND2xp5_ASAP7_75t_L g16853 ( 
.A(n_16745),
.B(n_2888),
.Y(n_16853)
);

NOR2xp33_ASAP7_75t_SL g16854 ( 
.A(n_16735),
.B(n_2889),
.Y(n_16854)
);

AOI21xp33_ASAP7_75t_L g16855 ( 
.A1(n_16695),
.A2(n_2890),
.B(n_2891),
.Y(n_16855)
);

NAND2xp5_ASAP7_75t_L g16856 ( 
.A(n_16757),
.B(n_2891),
.Y(n_16856)
);

OAI21xp33_ASAP7_75t_L g16857 ( 
.A1(n_16693),
.A2(n_2892),
.B(n_2893),
.Y(n_16857)
);

OAI21xp33_ASAP7_75t_SL g16858 ( 
.A1(n_16718),
.A2(n_2892),
.B(n_2893),
.Y(n_16858)
);

INVxp67_ASAP7_75t_L g16859 ( 
.A(n_16793),
.Y(n_16859)
);

AOI22xp5_ASAP7_75t_L g16860 ( 
.A1(n_16739),
.A2(n_2896),
.B1(n_2894),
.B2(n_2895),
.Y(n_16860)
);

INVx1_ASAP7_75t_L g16861 ( 
.A(n_16759),
.Y(n_16861)
);

NAND2xp5_ASAP7_75t_L g16862 ( 
.A(n_16760),
.B(n_2894),
.Y(n_16862)
);

INVxp67_ASAP7_75t_L g16863 ( 
.A(n_16767),
.Y(n_16863)
);

AOI22xp5_ASAP7_75t_L g16864 ( 
.A1(n_16696),
.A2(n_2897),
.B1(n_2895),
.B2(n_2896),
.Y(n_16864)
);

OAI32xp33_ASAP7_75t_L g16865 ( 
.A1(n_16778),
.A2(n_2899),
.A3(n_2897),
.B1(n_2898),
.B2(n_2900),
.Y(n_16865)
);

NAND2x1_ASAP7_75t_L g16866 ( 
.A(n_16802),
.B(n_2898),
.Y(n_16866)
);

INVx1_ASAP7_75t_L g16867 ( 
.A(n_16722),
.Y(n_16867)
);

OAI32xp33_ASAP7_75t_L g16868 ( 
.A1(n_16748),
.A2(n_2901),
.A3(n_2899),
.B1(n_2900),
.B2(n_2902),
.Y(n_16868)
);

INVx1_ASAP7_75t_L g16869 ( 
.A(n_16730),
.Y(n_16869)
);

AO21x1_ASAP7_75t_L g16870 ( 
.A1(n_16736),
.A2(n_16794),
.B(n_16788),
.Y(n_16870)
);

A2O1A1Ixp33_ASAP7_75t_L g16871 ( 
.A1(n_16796),
.A2(n_2903),
.B(n_2901),
.C(n_2902),
.Y(n_16871)
);

OAI22xp5_ASAP7_75t_L g16872 ( 
.A1(n_16783),
.A2(n_2905),
.B1(n_2903),
.B2(n_2904),
.Y(n_16872)
);

AOI22xp5_ASAP7_75t_L g16873 ( 
.A1(n_16712),
.A2(n_2906),
.B1(n_2904),
.B2(n_2905),
.Y(n_16873)
);

OAI21xp33_ASAP7_75t_L g16874 ( 
.A1(n_16801),
.A2(n_2906),
.B(n_2907),
.Y(n_16874)
);

INVx1_ASAP7_75t_L g16875 ( 
.A(n_16724),
.Y(n_16875)
);

OAI211xp5_ASAP7_75t_L g16876 ( 
.A1(n_16708),
.A2(n_2909),
.B(n_2907),
.C(n_2908),
.Y(n_16876)
);

AOI22xp5_ASAP7_75t_L g16877 ( 
.A1(n_16721),
.A2(n_2910),
.B1(n_2908),
.B2(n_2909),
.Y(n_16877)
);

AO22x1_ASAP7_75t_L g16878 ( 
.A1(n_16733),
.A2(n_2912),
.B1(n_2910),
.B2(n_2911),
.Y(n_16878)
);

INVxp67_ASAP7_75t_L g16879 ( 
.A(n_16782),
.Y(n_16879)
);

INVx1_ASAP7_75t_L g16880 ( 
.A(n_16805),
.Y(n_16880)
);

INVx1_ASAP7_75t_SL g16881 ( 
.A(n_16806),
.Y(n_16881)
);

AOI22xp5_ASAP7_75t_L g16882 ( 
.A1(n_16812),
.A2(n_16792),
.B1(n_16787),
.B2(n_16789),
.Y(n_16882)
);

OAI221xp5_ASAP7_75t_SL g16883 ( 
.A1(n_16728),
.A2(n_2915),
.B1(n_2913),
.B2(n_2914),
.C(n_2916),
.Y(n_16883)
);

INVx1_ASAP7_75t_L g16884 ( 
.A(n_16701),
.Y(n_16884)
);

OAI21xp33_ASAP7_75t_SL g16885 ( 
.A1(n_16743),
.A2(n_2913),
.B(n_2914),
.Y(n_16885)
);

INVx1_ASAP7_75t_SL g16886 ( 
.A(n_16762),
.Y(n_16886)
);

NAND4xp25_ASAP7_75t_L g16887 ( 
.A(n_16810),
.B(n_16727),
.C(n_16720),
.D(n_16770),
.Y(n_16887)
);

AOI32xp33_ASAP7_75t_L g16888 ( 
.A1(n_16738),
.A2(n_2918),
.A3(n_2915),
.B1(n_2917),
.B2(n_2919),
.Y(n_16888)
);

NAND4xp25_ASAP7_75t_L g16889 ( 
.A(n_16755),
.B(n_2921),
.C(n_2918),
.D(n_2920),
.Y(n_16889)
);

NAND2xp5_ASAP7_75t_L g16890 ( 
.A(n_16705),
.B(n_2920),
.Y(n_16890)
);

AOI222xp33_ASAP7_75t_L g16891 ( 
.A1(n_16765),
.A2(n_2923),
.B1(n_2925),
.B2(n_2921),
.C1(n_2922),
.C2(n_2924),
.Y(n_16891)
);

OAI22xp5_ASAP7_75t_L g16892 ( 
.A1(n_16703),
.A2(n_2924),
.B1(n_2922),
.B2(n_2923),
.Y(n_16892)
);

OAI21xp5_ASAP7_75t_L g16893 ( 
.A1(n_16758),
.A2(n_16756),
.B(n_16797),
.Y(n_16893)
);

NAND3xp33_ASAP7_75t_SL g16894 ( 
.A(n_16795),
.B(n_16744),
.C(n_16737),
.Y(n_16894)
);

OAI21xp5_ASAP7_75t_L g16895 ( 
.A1(n_16692),
.A2(n_2925),
.B(n_2926),
.Y(n_16895)
);

NOR4xp25_ASAP7_75t_L g16896 ( 
.A(n_16753),
.B(n_2928),
.C(n_2926),
.D(n_2927),
.Y(n_16896)
);

INVx1_ASAP7_75t_L g16897 ( 
.A(n_16715),
.Y(n_16897)
);

AOI21xp5_ASAP7_75t_L g16898 ( 
.A1(n_16761),
.A2(n_2928),
.B(n_2929),
.Y(n_16898)
);

AOI21xp33_ASAP7_75t_L g16899 ( 
.A1(n_16766),
.A2(n_2929),
.B(n_2930),
.Y(n_16899)
);

AOI22xp33_ASAP7_75t_SL g16900 ( 
.A1(n_16768),
.A2(n_2932),
.B1(n_2930),
.B2(n_2931),
.Y(n_16900)
);

INVx1_ASAP7_75t_L g16901 ( 
.A(n_16791),
.Y(n_16901)
);

OAI21xp5_ASAP7_75t_SL g16902 ( 
.A1(n_16769),
.A2(n_2931),
.B(n_2933),
.Y(n_16902)
);

AOI22xp5_ASAP7_75t_L g16903 ( 
.A1(n_16774),
.A2(n_2936),
.B1(n_2934),
.B2(n_2935),
.Y(n_16903)
);

NAND3xp33_ASAP7_75t_L g16904 ( 
.A(n_16746),
.B(n_2934),
.C(n_2935),
.Y(n_16904)
);

AOI21xp33_ASAP7_75t_L g16905 ( 
.A1(n_16815),
.A2(n_16764),
.B(n_16808),
.Y(n_16905)
);

INVx1_ASAP7_75t_L g16906 ( 
.A(n_16780),
.Y(n_16906)
);

NAND2xp5_ASAP7_75t_L g16907 ( 
.A(n_16752),
.B(n_2936),
.Y(n_16907)
);

NOR2xp67_ASAP7_75t_SL g16908 ( 
.A(n_16800),
.B(n_2937),
.Y(n_16908)
);

A2O1A1Ixp33_ASAP7_75t_L g16909 ( 
.A1(n_16779),
.A2(n_2939),
.B(n_2937),
.C(n_2938),
.Y(n_16909)
);

AOI22xp5_ASAP7_75t_L g16910 ( 
.A1(n_16740),
.A2(n_2941),
.B1(n_2939),
.B2(n_2940),
.Y(n_16910)
);

INVx1_ASAP7_75t_L g16911 ( 
.A(n_16809),
.Y(n_16911)
);

AOI21xp33_ASAP7_75t_L g16912 ( 
.A1(n_16691),
.A2(n_2940),
.B(n_2941),
.Y(n_16912)
);

INVx2_ASAP7_75t_L g16913 ( 
.A(n_16816),
.Y(n_16913)
);

INVx1_ASAP7_75t_L g16914 ( 
.A(n_16816),
.Y(n_16914)
);

OAI22xp5_ASAP7_75t_L g16915 ( 
.A1(n_16813),
.A2(n_2944),
.B1(n_2942),
.B2(n_2943),
.Y(n_16915)
);

INVx1_ASAP7_75t_L g16916 ( 
.A(n_16816),
.Y(n_16916)
);

OAI32xp33_ASAP7_75t_L g16917 ( 
.A1(n_16777),
.A2(n_2946),
.A3(n_2944),
.B1(n_2945),
.B2(n_2947),
.Y(n_16917)
);

AOI21xp33_ASAP7_75t_SL g16918 ( 
.A1(n_16709),
.A2(n_2945),
.B(n_2946),
.Y(n_16918)
);

NAND3xp33_ASAP7_75t_SL g16919 ( 
.A(n_16784),
.B(n_2948),
.C(n_2949),
.Y(n_16919)
);

OR2x2_ASAP7_75t_L g16920 ( 
.A(n_16709),
.B(n_2948),
.Y(n_16920)
);

A2O1A1Ixp33_ASAP7_75t_L g16921 ( 
.A1(n_16741),
.A2(n_2951),
.B(n_2949),
.C(n_2950),
.Y(n_16921)
);

CKINVDCx16_ASAP7_75t_R g16922 ( 
.A(n_16691),
.Y(n_16922)
);

AOI22xp5_ASAP7_75t_L g16923 ( 
.A1(n_16691),
.A2(n_2952),
.B1(n_2950),
.B2(n_2951),
.Y(n_16923)
);

OAI22xp5_ASAP7_75t_L g16924 ( 
.A1(n_16813),
.A2(n_2954),
.B1(n_2952),
.B2(n_2953),
.Y(n_16924)
);

OAI22xp33_ASAP7_75t_L g16925 ( 
.A1(n_16735),
.A2(n_2955),
.B1(n_2953),
.B2(n_2954),
.Y(n_16925)
);

INVxp67_ASAP7_75t_L g16926 ( 
.A(n_16735),
.Y(n_16926)
);

OAI21xp5_ASAP7_75t_L g16927 ( 
.A1(n_16691),
.A2(n_2955),
.B(n_2956),
.Y(n_16927)
);

HB1xp67_ASAP7_75t_L g16928 ( 
.A(n_16741),
.Y(n_16928)
);

A2O1A1Ixp33_ASAP7_75t_L g16929 ( 
.A1(n_16741),
.A2(n_2958),
.B(n_2956),
.C(n_2957),
.Y(n_16929)
);

OAI22xp5_ASAP7_75t_L g16930 ( 
.A1(n_16813),
.A2(n_2959),
.B1(n_2957),
.B2(n_2958),
.Y(n_16930)
);

INVx1_ASAP7_75t_L g16931 ( 
.A(n_16816),
.Y(n_16931)
);

OAI22xp5_ASAP7_75t_L g16932 ( 
.A1(n_16813),
.A2(n_2962),
.B1(n_2960),
.B2(n_2961),
.Y(n_16932)
);

OAI21xp33_ASAP7_75t_L g16933 ( 
.A1(n_16807),
.A2(n_2960),
.B(n_2962),
.Y(n_16933)
);

OAI22xp5_ASAP7_75t_L g16934 ( 
.A1(n_16813),
.A2(n_2965),
.B1(n_2963),
.B2(n_2964),
.Y(n_16934)
);

INVx1_ASAP7_75t_L g16935 ( 
.A(n_16816),
.Y(n_16935)
);

OAI222xp33_ASAP7_75t_L g16936 ( 
.A1(n_16697),
.A2(n_2966),
.B1(n_2968),
.B2(n_2964),
.C1(n_2965),
.C2(n_2967),
.Y(n_16936)
);

INVx1_ASAP7_75t_L g16937 ( 
.A(n_16816),
.Y(n_16937)
);

INVxp67_ASAP7_75t_L g16938 ( 
.A(n_16735),
.Y(n_16938)
);

O2A1O1Ixp33_ASAP7_75t_L g16939 ( 
.A1(n_16713),
.A2(n_2968),
.B(n_2966),
.C(n_2967),
.Y(n_16939)
);

AOI211xp5_ASAP7_75t_L g16940 ( 
.A1(n_16691),
.A2(n_2972),
.B(n_2969),
.C(n_2970),
.Y(n_16940)
);

AOI32xp33_ASAP7_75t_L g16941 ( 
.A1(n_16711),
.A2(n_2972),
.A3(n_2969),
.B1(n_2970),
.B2(n_2973),
.Y(n_16941)
);

NOR2xp33_ASAP7_75t_L g16942 ( 
.A(n_16793),
.B(n_2973),
.Y(n_16942)
);

OAI31xp33_ASAP7_75t_L g16943 ( 
.A1(n_16691),
.A2(n_2976),
.A3(n_2974),
.B(n_2975),
.Y(n_16943)
);

INVx1_ASAP7_75t_SL g16944 ( 
.A(n_16698),
.Y(n_16944)
);

OAI211xp5_ASAP7_75t_L g16945 ( 
.A1(n_16713),
.A2(n_2976),
.B(n_2974),
.C(n_2975),
.Y(n_16945)
);

O2A1O1Ixp33_ASAP7_75t_L g16946 ( 
.A1(n_16713),
.A2(n_2979),
.B(n_2977),
.C(n_2978),
.Y(n_16946)
);

O2A1O1Ixp33_ASAP7_75t_L g16947 ( 
.A1(n_16713),
.A2(n_2980),
.B(n_2977),
.C(n_2978),
.Y(n_16947)
);

O2A1O1Ixp33_ASAP7_75t_L g16948 ( 
.A1(n_16713),
.A2(n_2983),
.B(n_2981),
.C(n_2982),
.Y(n_16948)
);

OAI221xp5_ASAP7_75t_SL g16949 ( 
.A1(n_16837),
.A2(n_2983),
.B1(n_2981),
.B2(n_2982),
.C(n_2984),
.Y(n_16949)
);

NAND2xp5_ASAP7_75t_L g16950 ( 
.A(n_16878),
.B(n_2984),
.Y(n_16950)
);

AND2x2_ASAP7_75t_L g16951 ( 
.A(n_16848),
.B(n_2985),
.Y(n_16951)
);

OAI22xp33_ASAP7_75t_SL g16952 ( 
.A1(n_16922),
.A2(n_2987),
.B1(n_2985),
.B2(n_2986),
.Y(n_16952)
);

NAND3xp33_ASAP7_75t_SL g16953 ( 
.A(n_16854),
.B(n_2986),
.C(n_2987),
.Y(n_16953)
);

INVxp67_ASAP7_75t_L g16954 ( 
.A(n_16942),
.Y(n_16954)
);

AOI32xp33_ASAP7_75t_L g16955 ( 
.A1(n_16944),
.A2(n_2990),
.A3(n_2988),
.B1(n_2989),
.B2(n_2991),
.Y(n_16955)
);

AOI32xp33_ASAP7_75t_L g16956 ( 
.A1(n_16886),
.A2(n_2992),
.A3(n_2989),
.B1(n_2991),
.B2(n_2993),
.Y(n_16956)
);

AND2x2_ASAP7_75t_L g16957 ( 
.A(n_16851),
.B(n_2992),
.Y(n_16957)
);

A2O1A1Ixp33_ASAP7_75t_L g16958 ( 
.A1(n_16841),
.A2(n_2996),
.B(n_2994),
.C(n_2995),
.Y(n_16958)
);

NAND2xp5_ASAP7_75t_L g16959 ( 
.A(n_16896),
.B(n_2994),
.Y(n_16959)
);

AO22x1_ASAP7_75t_L g16960 ( 
.A1(n_16850),
.A2(n_2997),
.B1(n_2995),
.B2(n_2996),
.Y(n_16960)
);

OAI21xp33_ASAP7_75t_SL g16961 ( 
.A1(n_16943),
.A2(n_2997),
.B(n_2998),
.Y(n_16961)
);

INVx2_ASAP7_75t_L g16962 ( 
.A(n_16824),
.Y(n_16962)
);

AOI322xp5_ASAP7_75t_L g16963 ( 
.A1(n_16894),
.A2(n_3003),
.A3(n_3002),
.B1(n_3000),
.B2(n_2998),
.C1(n_2999),
.C2(n_3001),
.Y(n_16963)
);

INVx3_ASAP7_75t_L g16964 ( 
.A(n_16866),
.Y(n_16964)
);

NOR2xp33_ASAP7_75t_L g16965 ( 
.A(n_16818),
.B(n_2999),
.Y(n_16965)
);

INVx1_ASAP7_75t_L g16966 ( 
.A(n_16825),
.Y(n_16966)
);

NAND2xp5_ASAP7_75t_SL g16967 ( 
.A(n_16918),
.B(n_3000),
.Y(n_16967)
);

NAND2x1p5_ASAP7_75t_L g16968 ( 
.A(n_16822),
.B(n_3001),
.Y(n_16968)
);

AOI21xp33_ASAP7_75t_L g16969 ( 
.A1(n_16939),
.A2(n_3002),
.B(n_3003),
.Y(n_16969)
);

AO21x1_ASAP7_75t_L g16970 ( 
.A1(n_16843),
.A2(n_3004),
.B(n_3005),
.Y(n_16970)
);

OAI321xp33_ASAP7_75t_L g16971 ( 
.A1(n_16887),
.A2(n_3007),
.A3(n_3009),
.B1(n_3005),
.B2(n_3006),
.C(n_3008),
.Y(n_16971)
);

OAI21xp33_ASAP7_75t_L g16972 ( 
.A1(n_16882),
.A2(n_16933),
.B(n_16819),
.Y(n_16972)
);

NAND2xp5_ASAP7_75t_L g16973 ( 
.A(n_16834),
.B(n_3006),
.Y(n_16973)
);

INVx1_ASAP7_75t_SL g16974 ( 
.A(n_16920),
.Y(n_16974)
);

OAI21xp33_ASAP7_75t_L g16975 ( 
.A1(n_16857),
.A2(n_16859),
.B(n_16926),
.Y(n_16975)
);

INVx1_ASAP7_75t_L g16976 ( 
.A(n_16824),
.Y(n_16976)
);

INVx2_ASAP7_75t_SL g16977 ( 
.A(n_16928),
.Y(n_16977)
);

NAND4xp25_ASAP7_75t_L g16978 ( 
.A(n_16828),
.B(n_3011),
.C(n_3008),
.D(n_3010),
.Y(n_16978)
);

AND2x2_ASAP7_75t_L g16979 ( 
.A(n_16832),
.B(n_3011),
.Y(n_16979)
);

AND2x2_ASAP7_75t_L g16980 ( 
.A(n_16836),
.B(n_16861),
.Y(n_16980)
);

INVx1_ASAP7_75t_L g16981 ( 
.A(n_16853),
.Y(n_16981)
);

OAI21xp33_ASAP7_75t_L g16982 ( 
.A1(n_16938),
.A2(n_3012),
.B(n_3013),
.Y(n_16982)
);

NAND2xp5_ASAP7_75t_L g16983 ( 
.A(n_16823),
.B(n_3012),
.Y(n_16983)
);

OAI222xp33_ASAP7_75t_L g16984 ( 
.A1(n_16908),
.A2(n_3015),
.B1(n_3017),
.B2(n_3013),
.C1(n_3014),
.C2(n_3016),
.Y(n_16984)
);

AOI22xp33_ASAP7_75t_L g16985 ( 
.A1(n_16919),
.A2(n_3016),
.B1(n_3014),
.B2(n_3015),
.Y(n_16985)
);

AND2x2_ASAP7_75t_L g16986 ( 
.A(n_16913),
.B(n_3017),
.Y(n_16986)
);

AND2x2_ASAP7_75t_L g16987 ( 
.A(n_16881),
.B(n_3018),
.Y(n_16987)
);

INVx1_ASAP7_75t_L g16988 ( 
.A(n_16856),
.Y(n_16988)
);

OAI21xp33_ASAP7_75t_L g16989 ( 
.A1(n_16906),
.A2(n_3019),
.B(n_3020),
.Y(n_16989)
);

NAND2xp5_ASAP7_75t_L g16990 ( 
.A(n_16900),
.B(n_3021),
.Y(n_16990)
);

AND2x2_ASAP7_75t_L g16991 ( 
.A(n_16875),
.B(n_3021),
.Y(n_16991)
);

AND2x4_ASAP7_75t_L g16992 ( 
.A(n_16821),
.B(n_3022),
.Y(n_16992)
);

INVx2_ASAP7_75t_L g16993 ( 
.A(n_16844),
.Y(n_16993)
);

NAND2xp5_ASAP7_75t_L g16994 ( 
.A(n_16941),
.B(n_3022),
.Y(n_16994)
);

INVxp67_ASAP7_75t_SL g16995 ( 
.A(n_16946),
.Y(n_16995)
);

NAND2xp5_ASAP7_75t_L g16996 ( 
.A(n_16888),
.B(n_3023),
.Y(n_16996)
);

OAI321xp33_ASAP7_75t_L g16997 ( 
.A1(n_16893),
.A2(n_3026),
.A3(n_3028),
.B1(n_3023),
.B2(n_3025),
.C(n_3027),
.Y(n_16997)
);

OAI21xp33_ASAP7_75t_L g16998 ( 
.A1(n_16911),
.A2(n_3026),
.B(n_3027),
.Y(n_16998)
);

NAND2xp5_ASAP7_75t_L g16999 ( 
.A(n_16921),
.B(n_3029),
.Y(n_16999)
);

OAI211xp5_ASAP7_75t_L g17000 ( 
.A1(n_16858),
.A2(n_3031),
.B(n_3029),
.C(n_3030),
.Y(n_17000)
);

INVx1_ASAP7_75t_L g17001 ( 
.A(n_16862),
.Y(n_17001)
);

OAI21xp33_ASAP7_75t_SL g17002 ( 
.A1(n_16912),
.A2(n_3030),
.B(n_3031),
.Y(n_17002)
);

AOI221xp5_ASAP7_75t_L g17003 ( 
.A1(n_16917),
.A2(n_3034),
.B1(n_3032),
.B2(n_3033),
.C(n_3035),
.Y(n_17003)
);

AOI22xp5_ASAP7_75t_L g17004 ( 
.A1(n_16863),
.A2(n_3035),
.B1(n_3032),
.B2(n_3033),
.Y(n_17004)
);

INVx2_ASAP7_75t_L g17005 ( 
.A(n_16914),
.Y(n_17005)
);

HB1xp67_ASAP7_75t_L g17006 ( 
.A(n_16885),
.Y(n_17006)
);

AO22x1_ASAP7_75t_L g17007 ( 
.A1(n_16840),
.A2(n_3038),
.B1(n_3036),
.B2(n_3037),
.Y(n_17007)
);

AOI222xp33_ASAP7_75t_L g17008 ( 
.A1(n_16879),
.A2(n_16937),
.B1(n_16916),
.B2(n_16935),
.C1(n_16931),
.C2(n_16867),
.Y(n_17008)
);

AOI22xp5_ASAP7_75t_L g17009 ( 
.A1(n_16874),
.A2(n_3039),
.B1(n_3036),
.B2(n_3037),
.Y(n_17009)
);

HB1xp67_ASAP7_75t_L g17010 ( 
.A(n_16936),
.Y(n_17010)
);

AOI22xp5_ASAP7_75t_L g17011 ( 
.A1(n_16869),
.A2(n_3041),
.B1(n_3039),
.B2(n_3040),
.Y(n_17011)
);

AOI21xp33_ASAP7_75t_SL g17012 ( 
.A1(n_16925),
.A2(n_3040),
.B(n_3041),
.Y(n_17012)
);

AND2x2_ASAP7_75t_L g17013 ( 
.A(n_16927),
.B(n_3042),
.Y(n_17013)
);

OAI22xp5_ASAP7_75t_L g17014 ( 
.A1(n_16835),
.A2(n_3046),
.B1(n_3043),
.B2(n_3045),
.Y(n_17014)
);

NAND2xp5_ASAP7_75t_L g17015 ( 
.A(n_16929),
.B(n_3043),
.Y(n_17015)
);

INVx1_ASAP7_75t_L g17016 ( 
.A(n_16947),
.Y(n_17016)
);

OR2x2_ASAP7_75t_L g17017 ( 
.A(n_16890),
.B(n_3045),
.Y(n_17017)
);

AOI211xp5_ASAP7_75t_L g17018 ( 
.A1(n_16876),
.A2(n_3048),
.B(n_3046),
.C(n_3047),
.Y(n_17018)
);

OAI21xp33_ASAP7_75t_SL g17019 ( 
.A1(n_16905),
.A2(n_3047),
.B(n_3048),
.Y(n_17019)
);

INVx2_ASAP7_75t_SL g17020 ( 
.A(n_16880),
.Y(n_17020)
);

OAI21xp33_ASAP7_75t_L g17021 ( 
.A1(n_16830),
.A2(n_3049),
.B(n_3050),
.Y(n_17021)
);

NAND2xp5_ASAP7_75t_L g17022 ( 
.A(n_16940),
.B(n_3049),
.Y(n_17022)
);

OAI22xp5_ASAP7_75t_L g17023 ( 
.A1(n_16923),
.A2(n_3052),
.B1(n_3050),
.B2(n_3051),
.Y(n_17023)
);

INVx1_ASAP7_75t_L g17024 ( 
.A(n_16948),
.Y(n_17024)
);

AOI22xp5_ASAP7_75t_L g17025 ( 
.A1(n_16838),
.A2(n_3054),
.B1(n_3051),
.B2(n_3053),
.Y(n_17025)
);

AOI22xp5_ASAP7_75t_SL g17026 ( 
.A1(n_16915),
.A2(n_3055),
.B1(n_3053),
.B2(n_3054),
.Y(n_17026)
);

AOI22xp33_ASAP7_75t_SL g17027 ( 
.A1(n_16945),
.A2(n_3058),
.B1(n_3055),
.B2(n_3057),
.Y(n_17027)
);

OAI21xp5_ASAP7_75t_L g17028 ( 
.A1(n_16820),
.A2(n_3057),
.B(n_3059),
.Y(n_17028)
);

OAI21xp33_ASAP7_75t_L g17029 ( 
.A1(n_16884),
.A2(n_3059),
.B(n_3060),
.Y(n_17029)
);

AOI221xp5_ASAP7_75t_SL g17030 ( 
.A1(n_16839),
.A2(n_3063),
.B1(n_3061),
.B2(n_3062),
.C(n_3064),
.Y(n_17030)
);

A2O1A1Ixp33_ASAP7_75t_L g17031 ( 
.A1(n_16849),
.A2(n_3063),
.B(n_3061),
.C(n_3062),
.Y(n_17031)
);

NAND2xp5_ASAP7_75t_SL g17032 ( 
.A(n_16845),
.B(n_3064),
.Y(n_17032)
);

INVx1_ASAP7_75t_L g17033 ( 
.A(n_16826),
.Y(n_17033)
);

AOI31xp33_ASAP7_75t_L g17034 ( 
.A1(n_16870),
.A2(n_3067),
.A3(n_3065),
.B(n_3066),
.Y(n_17034)
);

INVx1_ASAP7_75t_L g17035 ( 
.A(n_16831),
.Y(n_17035)
);

O2A1O1Ixp33_ASAP7_75t_L g17036 ( 
.A1(n_16852),
.A2(n_3067),
.B(n_3065),
.C(n_3066),
.Y(n_17036)
);

OAI21xp33_ASAP7_75t_SL g17037 ( 
.A1(n_16907),
.A2(n_3068),
.B(n_3069),
.Y(n_17037)
);

NAND2xp5_ASAP7_75t_L g17038 ( 
.A(n_16871),
.B(n_3068),
.Y(n_17038)
);

NAND2xp5_ASAP7_75t_L g17039 ( 
.A(n_16902),
.B(n_3070),
.Y(n_17039)
);

INVx2_ASAP7_75t_L g17040 ( 
.A(n_16897),
.Y(n_17040)
);

OAI22xp5_ASAP7_75t_L g17041 ( 
.A1(n_16910),
.A2(n_3072),
.B1(n_3070),
.B2(n_3071),
.Y(n_17041)
);

NOR2xp33_ASAP7_75t_L g17042 ( 
.A(n_16889),
.B(n_3071),
.Y(n_17042)
);

OAI22xp5_ASAP7_75t_L g17043 ( 
.A1(n_16827),
.A2(n_3074),
.B1(n_3072),
.B2(n_3073),
.Y(n_17043)
);

OAI21xp5_ASAP7_75t_L g17044 ( 
.A1(n_16904),
.A2(n_3073),
.B(n_3074),
.Y(n_17044)
);

A2O1A1Ixp33_ASAP7_75t_L g17045 ( 
.A1(n_16898),
.A2(n_3077),
.B(n_3075),
.C(n_3076),
.Y(n_17045)
);

INVx2_ASAP7_75t_L g17046 ( 
.A(n_16901),
.Y(n_17046)
);

AOI222xp33_ASAP7_75t_L g17047 ( 
.A1(n_16842),
.A2(n_3077),
.B1(n_3079),
.B2(n_3075),
.C1(n_3076),
.C2(n_3078),
.Y(n_17047)
);

OAI31xp33_ASAP7_75t_L g17048 ( 
.A1(n_16846),
.A2(n_3081),
.A3(n_3079),
.B(n_3080),
.Y(n_17048)
);

OR2x2_ASAP7_75t_L g17049 ( 
.A(n_16909),
.B(n_3080),
.Y(n_17049)
);

OR2x2_ASAP7_75t_L g17050 ( 
.A(n_16872),
.B(n_3081),
.Y(n_17050)
);

OAI21xp33_ASAP7_75t_L g17051 ( 
.A1(n_16868),
.A2(n_3082),
.B(n_3083),
.Y(n_17051)
);

NAND2xp33_ASAP7_75t_SL g17052 ( 
.A(n_16924),
.B(n_3082),
.Y(n_17052)
);

INVx1_ASAP7_75t_L g17053 ( 
.A(n_16895),
.Y(n_17053)
);

AOI22xp5_ASAP7_75t_L g17054 ( 
.A1(n_16930),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.Y(n_17054)
);

INVx1_ASAP7_75t_SL g17055 ( 
.A(n_16855),
.Y(n_17055)
);

AOI22xp5_ASAP7_75t_L g17056 ( 
.A1(n_16932),
.A2(n_3086),
.B1(n_3084),
.B2(n_3085),
.Y(n_17056)
);

INVx1_ASAP7_75t_L g17057 ( 
.A(n_16934),
.Y(n_17057)
);

INVxp33_ASAP7_75t_L g17058 ( 
.A(n_16860),
.Y(n_17058)
);

AOI21xp33_ASAP7_75t_L g17059 ( 
.A1(n_16891),
.A2(n_3086),
.B(n_3087),
.Y(n_17059)
);

AOI221xp5_ASAP7_75t_L g17060 ( 
.A1(n_16865),
.A2(n_3089),
.B1(n_3087),
.B2(n_3088),
.C(n_3090),
.Y(n_17060)
);

NAND2xp33_ASAP7_75t_L g17061 ( 
.A(n_16829),
.B(n_3088),
.Y(n_17061)
);

AND2x2_ASAP7_75t_L g17062 ( 
.A(n_16899),
.B(n_3089),
.Y(n_17062)
);

INVx1_ASAP7_75t_L g17063 ( 
.A(n_16892),
.Y(n_17063)
);

NAND2xp5_ASAP7_75t_L g17064 ( 
.A(n_16873),
.B(n_3090),
.Y(n_17064)
);

OR2x2_ASAP7_75t_L g17065 ( 
.A(n_16883),
.B(n_3091),
.Y(n_17065)
);

INVx1_ASAP7_75t_L g17066 ( 
.A(n_16847),
.Y(n_17066)
);

INVx1_ASAP7_75t_L g17067 ( 
.A(n_16833),
.Y(n_17067)
);

INVx1_ASAP7_75t_L g17068 ( 
.A(n_16877),
.Y(n_17068)
);

AOI22xp5_ASAP7_75t_L g17069 ( 
.A1(n_16965),
.A2(n_16864),
.B1(n_16903),
.B2(n_3093),
.Y(n_17069)
);

AND4x1_ASAP7_75t_L g17070 ( 
.A(n_17008),
.B(n_3094),
.C(n_3091),
.D(n_3092),
.Y(n_17070)
);

XOR2x2_ASAP7_75t_L g17071 ( 
.A(n_17030),
.B(n_17018),
.Y(n_17071)
);

NOR2xp33_ASAP7_75t_L g17072 ( 
.A(n_16984),
.B(n_3092),
.Y(n_17072)
);

NAND3xp33_ASAP7_75t_SL g17073 ( 
.A(n_16963),
.B(n_3094),
.C(n_3095),
.Y(n_17073)
);

OAI21xp33_ASAP7_75t_SL g17074 ( 
.A1(n_16976),
.A2(n_3095),
.B(n_3096),
.Y(n_17074)
);

NAND2xp5_ASAP7_75t_L g17075 ( 
.A(n_16951),
.B(n_3096),
.Y(n_17075)
);

OAI211xp5_ASAP7_75t_L g17076 ( 
.A1(n_17027),
.A2(n_3099),
.B(n_3097),
.C(n_3098),
.Y(n_17076)
);

NOR3xp33_ASAP7_75t_L g17077 ( 
.A(n_16975),
.B(n_3097),
.C(n_3100),
.Y(n_17077)
);

OAI221xp5_ASAP7_75t_L g17078 ( 
.A1(n_16958),
.A2(n_3103),
.B1(n_3101),
.B2(n_3102),
.C(n_3104),
.Y(n_17078)
);

A2O1A1Ixp33_ASAP7_75t_L g17079 ( 
.A1(n_16956),
.A2(n_3106),
.B(n_3104),
.C(n_3105),
.Y(n_17079)
);

AOI222xp33_ASAP7_75t_L g17080 ( 
.A1(n_17019),
.A2(n_16961),
.B1(n_16966),
.B2(n_17061),
.C1(n_17052),
.C2(n_17002),
.Y(n_17080)
);

AOI222xp33_ASAP7_75t_L g17081 ( 
.A1(n_17051),
.A2(n_3109),
.B1(n_3111),
.B2(n_3107),
.C1(n_3108),
.C2(n_3110),
.Y(n_17081)
);

NAND2xp5_ASAP7_75t_L g17082 ( 
.A(n_16957),
.B(n_3107),
.Y(n_17082)
);

NAND2xp5_ASAP7_75t_L g17083 ( 
.A(n_16991),
.B(n_3108),
.Y(n_17083)
);

AOI21xp33_ASAP7_75t_SL g17084 ( 
.A1(n_17034),
.A2(n_3109),
.B(n_3110),
.Y(n_17084)
);

NOR2xp33_ASAP7_75t_L g17085 ( 
.A(n_16978),
.B(n_16964),
.Y(n_17085)
);

AOI221xp5_ASAP7_75t_L g17086 ( 
.A1(n_17012),
.A2(n_3114),
.B1(n_3111),
.B2(n_3112),
.C(n_3115),
.Y(n_17086)
);

AOI21xp5_ASAP7_75t_L g17087 ( 
.A1(n_17006),
.A2(n_3114),
.B(n_3115),
.Y(n_17087)
);

NAND2xp5_ASAP7_75t_L g17088 ( 
.A(n_16964),
.B(n_3116),
.Y(n_17088)
);

AOI32xp33_ASAP7_75t_L g17089 ( 
.A1(n_17058),
.A2(n_3118),
.A3(n_3116),
.B1(n_3117),
.B2(n_3119),
.Y(n_17089)
);

AOI211x1_ASAP7_75t_L g17090 ( 
.A1(n_16970),
.A2(n_17059),
.B(n_17000),
.C(n_16969),
.Y(n_17090)
);

OAI22xp5_ASAP7_75t_L g17091 ( 
.A1(n_16985),
.A2(n_3121),
.B1(n_3119),
.B2(n_3120),
.Y(n_17091)
);

OAI22xp33_ASAP7_75t_SL g17092 ( 
.A1(n_16962),
.A2(n_3122),
.B1(n_3120),
.B2(n_3121),
.Y(n_17092)
);

AOI211xp5_ASAP7_75t_L g17093 ( 
.A1(n_17043),
.A2(n_3124),
.B(n_3122),
.C(n_3123),
.Y(n_17093)
);

NAND3xp33_ASAP7_75t_L g17094 ( 
.A(n_17060),
.B(n_3123),
.C(n_3124),
.Y(n_17094)
);

NOR2xp33_ASAP7_75t_L g17095 ( 
.A(n_16982),
.B(n_3125),
.Y(n_17095)
);

OAI22xp33_ASAP7_75t_L g17096 ( 
.A1(n_17025),
.A2(n_3127),
.B1(n_3125),
.B2(n_3126),
.Y(n_17096)
);

INVx2_ASAP7_75t_L g17097 ( 
.A(n_16968),
.Y(n_17097)
);

AOI21xp5_ASAP7_75t_L g17098 ( 
.A1(n_16967),
.A2(n_3126),
.B(n_3127),
.Y(n_17098)
);

NOR3xp33_ASAP7_75t_L g17099 ( 
.A(n_16972),
.B(n_3128),
.C(n_3129),
.Y(n_17099)
);

A2O1A1Ixp33_ASAP7_75t_L g17100 ( 
.A1(n_17036),
.A2(n_3131),
.B(n_3129),
.C(n_3130),
.Y(n_17100)
);

AOI21xp5_ASAP7_75t_L g17101 ( 
.A1(n_16959),
.A2(n_3130),
.B(n_3131),
.Y(n_17101)
);

OAI21xp33_ASAP7_75t_L g17102 ( 
.A1(n_17020),
.A2(n_3132),
.B(n_3133),
.Y(n_17102)
);

AOI322xp5_ASAP7_75t_L g17103 ( 
.A1(n_16977),
.A2(n_3137),
.A3(n_3136),
.B1(n_3134),
.B2(n_3132),
.C1(n_3133),
.C2(n_3135),
.Y(n_17103)
);

NAND2xp5_ASAP7_75t_L g17104 ( 
.A(n_16979),
.B(n_3134),
.Y(n_17104)
);

OAI22xp5_ASAP7_75t_L g17105 ( 
.A1(n_17009),
.A2(n_3138),
.B1(n_3136),
.B2(n_3137),
.Y(n_17105)
);

OAI31xp33_ASAP7_75t_L g17106 ( 
.A1(n_16952),
.A2(n_3141),
.A3(n_3138),
.B(n_3139),
.Y(n_17106)
);

AOI221xp5_ASAP7_75t_L g17107 ( 
.A1(n_16995),
.A2(n_3142),
.B1(n_3139),
.B2(n_3141),
.C(n_3143),
.Y(n_17107)
);

INVx1_ASAP7_75t_SL g17108 ( 
.A(n_16986),
.Y(n_17108)
);

AOI21xp33_ASAP7_75t_L g17109 ( 
.A1(n_17065),
.A2(n_3143),
.B(n_3144),
.Y(n_17109)
);

OAI22xp5_ASAP7_75t_L g17110 ( 
.A1(n_17054),
.A2(n_3146),
.B1(n_3144),
.B2(n_3145),
.Y(n_17110)
);

NOR2xp33_ASAP7_75t_L g17111 ( 
.A(n_16998),
.B(n_3146),
.Y(n_17111)
);

OAI211xp5_ASAP7_75t_L g17112 ( 
.A1(n_17003),
.A2(n_3149),
.B(n_3147),
.C(n_3148),
.Y(n_17112)
);

INVx2_ASAP7_75t_L g17113 ( 
.A(n_16992),
.Y(n_17113)
);

NAND3xp33_ASAP7_75t_L g17114 ( 
.A(n_17047),
.B(n_16955),
.C(n_17031),
.Y(n_17114)
);

NAND2xp5_ASAP7_75t_L g17115 ( 
.A(n_17007),
.B(n_3147),
.Y(n_17115)
);

NAND2xp5_ASAP7_75t_L g17116 ( 
.A(n_17026),
.B(n_3148),
.Y(n_17116)
);

NAND2x1_ASAP7_75t_SL g17117 ( 
.A(n_17010),
.B(n_3149),
.Y(n_17117)
);

OAI32xp33_ASAP7_75t_L g17118 ( 
.A1(n_16950),
.A2(n_3152),
.A3(n_3150),
.B1(n_3151),
.B2(n_3153),
.Y(n_17118)
);

OAI22xp33_ASAP7_75t_L g17119 ( 
.A1(n_17056),
.A2(n_16983),
.B1(n_16990),
.B2(n_16973),
.Y(n_17119)
);

NAND2xp5_ASAP7_75t_L g17120 ( 
.A(n_16987),
.B(n_3150),
.Y(n_17120)
);

AOI22xp5_ASAP7_75t_L g17121 ( 
.A1(n_17042),
.A2(n_3153),
.B1(n_3151),
.B2(n_3152),
.Y(n_17121)
);

AOI22xp5_ASAP7_75t_L g17122 ( 
.A1(n_17005),
.A2(n_3156),
.B1(n_3154),
.B2(n_3155),
.Y(n_17122)
);

NAND3xp33_ASAP7_75t_SL g17123 ( 
.A(n_16974),
.B(n_3155),
.C(n_3157),
.Y(n_17123)
);

O2A1O1Ixp33_ASAP7_75t_L g17124 ( 
.A1(n_17045),
.A2(n_3159),
.B(n_3157),
.C(n_3158),
.Y(n_17124)
);

OAI22xp33_ASAP7_75t_L g17125 ( 
.A1(n_17038),
.A2(n_3161),
.B1(n_3158),
.B2(n_3159),
.Y(n_17125)
);

NAND2xp5_ASAP7_75t_SL g17126 ( 
.A(n_16971),
.B(n_3161),
.Y(n_17126)
);

OAI22xp5_ASAP7_75t_L g17127 ( 
.A1(n_16949),
.A2(n_3164),
.B1(n_3162),
.B2(n_3163),
.Y(n_17127)
);

AOI22xp5_ASAP7_75t_L g17128 ( 
.A1(n_16980),
.A2(n_3167),
.B1(n_3165),
.B2(n_3166),
.Y(n_17128)
);

AOI21xp33_ASAP7_75t_L g17129 ( 
.A1(n_17037),
.A2(n_3165),
.B(n_3167),
.Y(n_17129)
);

AO22x2_ASAP7_75t_L g17130 ( 
.A1(n_17057),
.A2(n_3170),
.B1(n_3168),
.B2(n_3169),
.Y(n_17130)
);

NOR2x1_ASAP7_75t_SL g17131 ( 
.A(n_16953),
.B(n_3168),
.Y(n_17131)
);

AOI21xp33_ASAP7_75t_L g17132 ( 
.A1(n_16994),
.A2(n_3169),
.B(n_3172),
.Y(n_17132)
);

NOR3xp33_ASAP7_75t_L g17133 ( 
.A(n_17016),
.B(n_3172),
.C(n_3173),
.Y(n_17133)
);

INVx1_ASAP7_75t_L g17134 ( 
.A(n_16992),
.Y(n_17134)
);

NAND2xp5_ASAP7_75t_L g17135 ( 
.A(n_16960),
.B(n_3173),
.Y(n_17135)
);

AOI22xp5_ASAP7_75t_L g17136 ( 
.A1(n_16954),
.A2(n_3176),
.B1(n_3174),
.B2(n_3175),
.Y(n_17136)
);

NAND4xp25_ASAP7_75t_L g17137 ( 
.A(n_17048),
.B(n_3177),
.C(n_3174),
.D(n_3175),
.Y(n_17137)
);

AOI322xp5_ASAP7_75t_L g17138 ( 
.A1(n_17055),
.A2(n_17024),
.A3(n_17067),
.B1(n_17035),
.B2(n_17033),
.C1(n_17066),
.C2(n_17068),
.Y(n_17138)
);

OAI22xp5_ASAP7_75t_L g17139 ( 
.A1(n_16996),
.A2(n_3179),
.B1(n_3177),
.B2(n_3178),
.Y(n_17139)
);

OAI22xp5_ASAP7_75t_L g17140 ( 
.A1(n_17039),
.A2(n_3180),
.B1(n_3178),
.B2(n_3179),
.Y(n_17140)
);

AOI21xp5_ASAP7_75t_L g17141 ( 
.A1(n_17032),
.A2(n_17015),
.B(n_16999),
.Y(n_17141)
);

OAI21xp5_ASAP7_75t_L g17142 ( 
.A1(n_17044),
.A2(n_3180),
.B(n_3181),
.Y(n_17142)
);

AOI221xp5_ASAP7_75t_L g17143 ( 
.A1(n_17021),
.A2(n_3183),
.B1(n_3181),
.B2(n_3182),
.C(n_3184),
.Y(n_17143)
);

OAI21xp5_ASAP7_75t_SL g17144 ( 
.A1(n_17013),
.A2(n_3182),
.B(n_3183),
.Y(n_17144)
);

AOI221x1_ASAP7_75t_L g17145 ( 
.A1(n_17063),
.A2(n_3186),
.B1(n_3184),
.B2(n_3185),
.C(n_3187),
.Y(n_17145)
);

AND2x2_ASAP7_75t_L g17146 ( 
.A(n_17062),
.B(n_3185),
.Y(n_17146)
);

INVx1_ASAP7_75t_L g17147 ( 
.A(n_17022),
.Y(n_17147)
);

OAI21xp5_ASAP7_75t_L g17148 ( 
.A1(n_17028),
.A2(n_3186),
.B(n_3188),
.Y(n_17148)
);

AND2x2_ASAP7_75t_L g17149 ( 
.A(n_17053),
.B(n_3188),
.Y(n_17149)
);

NAND2xp5_ASAP7_75t_SL g17150 ( 
.A(n_16997),
.B(n_3189),
.Y(n_17150)
);

AOI21xp33_ASAP7_75t_L g17151 ( 
.A1(n_17017),
.A2(n_3189),
.B(n_3190),
.Y(n_17151)
);

OAI32xp33_ASAP7_75t_L g17152 ( 
.A1(n_17049),
.A2(n_3192),
.A3(n_3190),
.B1(n_3191),
.B2(n_3193),
.Y(n_17152)
);

OAI21xp33_ASAP7_75t_L g17153 ( 
.A1(n_16993),
.A2(n_3191),
.B(n_3192),
.Y(n_17153)
);

OAI22xp5_ASAP7_75t_L g17154 ( 
.A1(n_17040),
.A2(n_3195),
.B1(n_3193),
.B2(n_3194),
.Y(n_17154)
);

AOI22xp33_ASAP7_75t_L g17155 ( 
.A1(n_17046),
.A2(n_3196),
.B1(n_3194),
.B2(n_3195),
.Y(n_17155)
);

OAI21xp33_ASAP7_75t_L g17156 ( 
.A1(n_16981),
.A2(n_3196),
.B(n_3197),
.Y(n_17156)
);

AOI221xp5_ASAP7_75t_L g17157 ( 
.A1(n_17023),
.A2(n_3200),
.B1(n_3198),
.B2(n_3199),
.C(n_3201),
.Y(n_17157)
);

NAND3xp33_ASAP7_75t_SL g17158 ( 
.A(n_17050),
.B(n_3198),
.C(n_3199),
.Y(n_17158)
);

OR2x2_ASAP7_75t_L g17159 ( 
.A(n_17064),
.B(n_3202),
.Y(n_17159)
);

OAI221xp5_ASAP7_75t_L g17160 ( 
.A1(n_16989),
.A2(n_3204),
.B1(n_3202),
.B2(n_3203),
.C(n_3205),
.Y(n_17160)
);

OAI221xp5_ASAP7_75t_L g17161 ( 
.A1(n_17029),
.A2(n_3205),
.B1(n_3203),
.B2(n_3204),
.C(n_3206),
.Y(n_17161)
);

NAND2xp5_ASAP7_75t_L g17162 ( 
.A(n_17004),
.B(n_3207),
.Y(n_17162)
);

NOR2xp33_ASAP7_75t_L g17163 ( 
.A(n_17014),
.B(n_17041),
.Y(n_17163)
);

AND2x2_ASAP7_75t_L g17164 ( 
.A(n_16988),
.B(n_3207),
.Y(n_17164)
);

INVx1_ASAP7_75t_L g17165 ( 
.A(n_17001),
.Y(n_17165)
);

AOI21xp33_ASAP7_75t_L g17166 ( 
.A1(n_17011),
.A2(n_3208),
.B(n_3209),
.Y(n_17166)
);

AOI21xp5_ASAP7_75t_L g17167 ( 
.A1(n_17006),
.A2(n_3208),
.B(n_3209),
.Y(n_17167)
);

AOI211xp5_ASAP7_75t_L g17168 ( 
.A1(n_16984),
.A2(n_3212),
.B(n_3210),
.C(n_3211),
.Y(n_17168)
);

NAND2xp5_ASAP7_75t_L g17169 ( 
.A(n_16951),
.B(n_3210),
.Y(n_17169)
);

INVx1_ASAP7_75t_L g17170 ( 
.A(n_16976),
.Y(n_17170)
);

NAND2xp5_ASAP7_75t_L g17171 ( 
.A(n_16951),
.B(n_3211),
.Y(n_17171)
);

OAI22xp33_ASAP7_75t_L g17172 ( 
.A1(n_17034),
.A2(n_3214),
.B1(n_3212),
.B2(n_3213),
.Y(n_17172)
);

AOI21xp33_ASAP7_75t_SL g17173 ( 
.A1(n_17034),
.A2(n_3213),
.B(n_3214),
.Y(n_17173)
);

AOI22xp5_ASAP7_75t_L g17174 ( 
.A1(n_16965),
.A2(n_3217),
.B1(n_3215),
.B2(n_3216),
.Y(n_17174)
);

NAND3xp33_ASAP7_75t_SL g17175 ( 
.A(n_16963),
.B(n_3215),
.C(n_3216),
.Y(n_17175)
);

NOR3xp33_ASAP7_75t_L g17176 ( 
.A(n_16975),
.B(n_3217),
.C(n_3218),
.Y(n_17176)
);

OR2x2_ASAP7_75t_L g17177 ( 
.A(n_16964),
.B(n_3219),
.Y(n_17177)
);

OAI21xp33_ASAP7_75t_L g17178 ( 
.A1(n_16975),
.A2(n_3219),
.B(n_3220),
.Y(n_17178)
);

AO22x2_ASAP7_75t_L g17179 ( 
.A1(n_16976),
.A2(n_3222),
.B1(n_3220),
.B2(n_3221),
.Y(n_17179)
);

AOI21xp5_ASAP7_75t_L g17180 ( 
.A1(n_17006),
.A2(n_3221),
.B(n_3222),
.Y(n_17180)
);

AOI221xp5_ASAP7_75t_L g17181 ( 
.A1(n_17012),
.A2(n_3225),
.B1(n_3223),
.B2(n_3224),
.C(n_3226),
.Y(n_17181)
);

OAI21xp33_ASAP7_75t_L g17182 ( 
.A1(n_16975),
.A2(n_3223),
.B(n_3224),
.Y(n_17182)
);

AOI21xp5_ASAP7_75t_L g17183 ( 
.A1(n_17088),
.A2(n_3226),
.B(n_3227),
.Y(n_17183)
);

NAND3xp33_ASAP7_75t_SL g17184 ( 
.A(n_17070),
.B(n_3227),
.C(n_3229),
.Y(n_17184)
);

OAI22xp5_ASAP7_75t_L g17185 ( 
.A1(n_17174),
.A2(n_3231),
.B1(n_3229),
.B2(n_3230),
.Y(n_17185)
);

INVx1_ASAP7_75t_L g17186 ( 
.A(n_17149),
.Y(n_17186)
);

NOR2xp67_ASAP7_75t_L g17187 ( 
.A(n_17123),
.B(n_3231),
.Y(n_17187)
);

AOI221xp5_ASAP7_75t_L g17188 ( 
.A1(n_17084),
.A2(n_3234),
.B1(n_3232),
.B2(n_3233),
.C(n_3235),
.Y(n_17188)
);

INVx1_ASAP7_75t_L g17189 ( 
.A(n_17135),
.Y(n_17189)
);

INVx1_ASAP7_75t_L g17190 ( 
.A(n_17117),
.Y(n_17190)
);

AOI322xp5_ASAP7_75t_L g17191 ( 
.A1(n_17085),
.A2(n_3237),
.A3(n_3236),
.B1(n_3234),
.B2(n_3232),
.C1(n_3233),
.C2(n_3235),
.Y(n_17191)
);

AOI22xp5_ASAP7_75t_L g17192 ( 
.A1(n_17077),
.A2(n_3238),
.B1(n_3236),
.B2(n_3237),
.Y(n_17192)
);

AOI21xp33_ASAP7_75t_SL g17193 ( 
.A1(n_17172),
.A2(n_3238),
.B(n_3239),
.Y(n_17193)
);

NAND4xp25_ASAP7_75t_L g17194 ( 
.A(n_17138),
.B(n_3241),
.C(n_3239),
.D(n_3240),
.Y(n_17194)
);

AOI22xp5_ASAP7_75t_L g17195 ( 
.A1(n_17176),
.A2(n_3243),
.B1(n_3240),
.B2(n_3242),
.Y(n_17195)
);

OA21x2_ASAP7_75t_L g17196 ( 
.A1(n_17170),
.A2(n_3242),
.B(n_3244),
.Y(n_17196)
);

AO22x1_ASAP7_75t_L g17197 ( 
.A1(n_17133),
.A2(n_3246),
.B1(n_3244),
.B2(n_3245),
.Y(n_17197)
);

NOR3xp33_ASAP7_75t_SL g17198 ( 
.A(n_17073),
.B(n_17175),
.C(n_17158),
.Y(n_17198)
);

AOI221xp5_ASAP7_75t_L g17199 ( 
.A1(n_17173),
.A2(n_3247),
.B1(n_3245),
.B2(n_3246),
.C(n_3248),
.Y(n_17199)
);

OAI21xp33_ASAP7_75t_L g17200 ( 
.A1(n_17072),
.A2(n_3247),
.B(n_3248),
.Y(n_17200)
);

NOR3xp33_ASAP7_75t_L g17201 ( 
.A(n_17109),
.B(n_3249),
.C(n_3250),
.Y(n_17201)
);

O2A1O1Ixp33_ASAP7_75t_L g17202 ( 
.A1(n_17074),
.A2(n_3251),
.B(n_3249),
.C(n_3250),
.Y(n_17202)
);

AOI33xp33_ASAP7_75t_L g17203 ( 
.A1(n_17119),
.A2(n_3253),
.A3(n_3255),
.B1(n_3251),
.B2(n_3252),
.B3(n_3254),
.Y(n_17203)
);

AND2x2_ASAP7_75t_L g17204 ( 
.A(n_17146),
.B(n_3252),
.Y(n_17204)
);

AOI21xp5_ASAP7_75t_L g17205 ( 
.A1(n_17129),
.A2(n_3253),
.B(n_3255),
.Y(n_17205)
);

AOI222xp33_ASAP7_75t_L g17206 ( 
.A1(n_17150),
.A2(n_3258),
.B1(n_3260),
.B2(n_3256),
.C1(n_3257),
.C2(n_3259),
.Y(n_17206)
);

AOI221xp5_ASAP7_75t_L g17207 ( 
.A1(n_17132),
.A2(n_3260),
.B1(n_3257),
.B2(n_3259),
.C(n_3261),
.Y(n_17207)
);

NOR3xp33_ASAP7_75t_L g17208 ( 
.A(n_17139),
.B(n_3261),
.C(n_3262),
.Y(n_17208)
);

AOI21xp5_ASAP7_75t_L g17209 ( 
.A1(n_17101),
.A2(n_3262),
.B(n_3263),
.Y(n_17209)
);

AOI322xp5_ASAP7_75t_L g17210 ( 
.A1(n_17126),
.A2(n_3269),
.A3(n_3268),
.B1(n_3266),
.B2(n_3264),
.C1(n_3265),
.C2(n_3267),
.Y(n_17210)
);

OAI221xp5_ASAP7_75t_L g17211 ( 
.A1(n_17106),
.A2(n_3266),
.B1(n_3264),
.B2(n_3265),
.C(n_3267),
.Y(n_17211)
);

AOI21xp33_ASAP7_75t_L g17212 ( 
.A1(n_17080),
.A2(n_3268),
.B(n_3269),
.Y(n_17212)
);

OAI211xp5_ASAP7_75t_SL g17213 ( 
.A1(n_17069),
.A2(n_3272),
.B(n_3270),
.C(n_3271),
.Y(n_17213)
);

OAI211xp5_ASAP7_75t_L g17214 ( 
.A1(n_17081),
.A2(n_3272),
.B(n_3270),
.C(n_3271),
.Y(n_17214)
);

NOR2xp33_ASAP7_75t_L g17215 ( 
.A(n_17178),
.B(n_3273),
.Y(n_17215)
);

AOI221xp5_ASAP7_75t_L g17216 ( 
.A1(n_17127),
.A2(n_3275),
.B1(n_3273),
.B2(n_3274),
.C(n_3276),
.Y(n_17216)
);

NAND4xp25_ASAP7_75t_L g17217 ( 
.A(n_17168),
.B(n_3276),
.C(n_3274),
.D(n_3275),
.Y(n_17217)
);

AOI21xp5_ASAP7_75t_L g17218 ( 
.A1(n_17087),
.A2(n_17180),
.B(n_17167),
.Y(n_17218)
);

AOI221xp5_ASAP7_75t_L g17219 ( 
.A1(n_17090),
.A2(n_3279),
.B1(n_3277),
.B2(n_3278),
.C(n_3280),
.Y(n_17219)
);

AOI221xp5_ASAP7_75t_L g17220 ( 
.A1(n_17166),
.A2(n_3280),
.B1(n_3277),
.B2(n_3278),
.C(n_3281),
.Y(n_17220)
);

AOI21xp5_ASAP7_75t_L g17221 ( 
.A1(n_17115),
.A2(n_3281),
.B(n_3282),
.Y(n_17221)
);

AOI22xp5_ASAP7_75t_L g17222 ( 
.A1(n_17099),
.A2(n_3284),
.B1(n_3282),
.B2(n_3283),
.Y(n_17222)
);

AOI221xp5_ASAP7_75t_L g17223 ( 
.A1(n_17137),
.A2(n_17124),
.B1(n_17094),
.B2(n_17112),
.C(n_17079),
.Y(n_17223)
);

INVx1_ASAP7_75t_L g17224 ( 
.A(n_17075),
.Y(n_17224)
);

OAI22xp5_ASAP7_75t_L g17225 ( 
.A1(n_17121),
.A2(n_17160),
.B1(n_17161),
.B2(n_17114),
.Y(n_17225)
);

OAI22xp5_ASAP7_75t_L g17226 ( 
.A1(n_17169),
.A2(n_3285),
.B1(n_3283),
.B2(n_3284),
.Y(n_17226)
);

NAND4xp25_ASAP7_75t_L g17227 ( 
.A(n_17163),
.B(n_3287),
.C(n_3285),
.D(n_3286),
.Y(n_17227)
);

OAI22xp33_ASAP7_75t_L g17228 ( 
.A1(n_17116),
.A2(n_3288),
.B1(n_3286),
.B2(n_3287),
.Y(n_17228)
);

AND2x2_ASAP7_75t_L g17229 ( 
.A(n_17113),
.B(n_3288),
.Y(n_17229)
);

AOI21xp33_ASAP7_75t_L g17230 ( 
.A1(n_17159),
.A2(n_3289),
.B(n_3290),
.Y(n_17230)
);

AOI221xp5_ASAP7_75t_L g17231 ( 
.A1(n_17091),
.A2(n_3291),
.B1(n_3289),
.B2(n_3290),
.C(n_3292),
.Y(n_17231)
);

AOI21xp5_ASAP7_75t_L g17232 ( 
.A1(n_17098),
.A2(n_3291),
.B(n_3292),
.Y(n_17232)
);

AND5x1_ASAP7_75t_L g17233 ( 
.A(n_17141),
.B(n_17111),
.C(n_17095),
.D(n_17181),
.E(n_17086),
.Y(n_17233)
);

AOI221xp5_ASAP7_75t_L g17234 ( 
.A1(n_17076),
.A2(n_3295),
.B1(n_3293),
.B2(n_3294),
.C(n_3296),
.Y(n_17234)
);

OAI21xp5_ASAP7_75t_SL g17235 ( 
.A1(n_17144),
.A2(n_17108),
.B(n_17142),
.Y(n_17235)
);

OAI22xp33_ASAP7_75t_L g17236 ( 
.A1(n_17171),
.A2(n_3296),
.B1(n_3294),
.B2(n_3295),
.Y(n_17236)
);

AOI211x1_ASAP7_75t_L g17237 ( 
.A1(n_17148),
.A2(n_3299),
.B(n_3297),
.C(n_3298),
.Y(n_17237)
);

AOI221x1_ASAP7_75t_SL g17238 ( 
.A1(n_17134),
.A2(n_3299),
.B1(n_3297),
.B2(n_3298),
.C(n_3300),
.Y(n_17238)
);

AOI221x1_ASAP7_75t_L g17239 ( 
.A1(n_17182),
.A2(n_17165),
.B1(n_17097),
.B2(n_17092),
.C(n_17120),
.Y(n_17239)
);

AOI22xp5_ASAP7_75t_L g17240 ( 
.A1(n_17105),
.A2(n_17110),
.B1(n_17071),
.B2(n_17143),
.Y(n_17240)
);

AOI222xp33_ASAP7_75t_L g17241 ( 
.A1(n_17131),
.A2(n_3302),
.B1(n_3304),
.B2(n_3300),
.C1(n_3301),
.C2(n_3303),
.Y(n_17241)
);

NOR2xp33_ASAP7_75t_L g17242 ( 
.A(n_17102),
.B(n_3303),
.Y(n_17242)
);

AO21x1_ASAP7_75t_L g17243 ( 
.A1(n_17082),
.A2(n_3304),
.B(n_3305),
.Y(n_17243)
);

INVx1_ASAP7_75t_L g17244 ( 
.A(n_17177),
.Y(n_17244)
);

OA21x2_ASAP7_75t_L g17245 ( 
.A1(n_17083),
.A2(n_3305),
.B(n_3306),
.Y(n_17245)
);

INVx1_ASAP7_75t_SL g17246 ( 
.A(n_17164),
.Y(n_17246)
);

AOI21xp5_ASAP7_75t_L g17247 ( 
.A1(n_17100),
.A2(n_17104),
.B(n_17162),
.Y(n_17247)
);

AOI21xp5_ASAP7_75t_SL g17248 ( 
.A1(n_17145),
.A2(n_3306),
.B(n_3307),
.Y(n_17248)
);

O2A1O1Ixp5_ASAP7_75t_L g17249 ( 
.A1(n_17147),
.A2(n_3309),
.B(n_3307),
.C(n_3308),
.Y(n_17249)
);

OAI221xp5_ASAP7_75t_L g17250 ( 
.A1(n_17093),
.A2(n_3311),
.B1(n_3308),
.B2(n_3309),
.C(n_3312),
.Y(n_17250)
);

OAI211xp5_ASAP7_75t_SL g17251 ( 
.A1(n_17157),
.A2(n_3313),
.B(n_3311),
.C(n_3312),
.Y(n_17251)
);

NOR2xp33_ASAP7_75t_L g17252 ( 
.A(n_17153),
.B(n_3314),
.Y(n_17252)
);

INVx1_ASAP7_75t_L g17253 ( 
.A(n_17179),
.Y(n_17253)
);

AOI211xp5_ASAP7_75t_L g17254 ( 
.A1(n_17096),
.A2(n_3316),
.B(n_3314),
.C(n_3315),
.Y(n_17254)
);

OAI211xp5_ASAP7_75t_L g17255 ( 
.A1(n_17118),
.A2(n_3317),
.B(n_3315),
.C(n_3316),
.Y(n_17255)
);

OAI21xp33_ASAP7_75t_L g17256 ( 
.A1(n_17089),
.A2(n_3317),
.B(n_3318),
.Y(n_17256)
);

NAND2xp5_ASAP7_75t_SL g17257 ( 
.A(n_17125),
.B(n_3318),
.Y(n_17257)
);

INVx1_ASAP7_75t_L g17258 ( 
.A(n_17179),
.Y(n_17258)
);

AOI22xp5_ASAP7_75t_L g17259 ( 
.A1(n_17078),
.A2(n_3321),
.B1(n_3319),
.B2(n_3320),
.Y(n_17259)
);

OAI21xp33_ASAP7_75t_L g17260 ( 
.A1(n_17156),
.A2(n_3319),
.B(n_3320),
.Y(n_17260)
);

AOI21xp5_ASAP7_75t_L g17261 ( 
.A1(n_17152),
.A2(n_3321),
.B(n_3322),
.Y(n_17261)
);

AOI21xp5_ASAP7_75t_L g17262 ( 
.A1(n_17151),
.A2(n_3323),
.B(n_3324),
.Y(n_17262)
);

NOR2xp33_ASAP7_75t_L g17263 ( 
.A(n_17140),
.B(n_3323),
.Y(n_17263)
);

OAI21xp5_ASAP7_75t_L g17264 ( 
.A1(n_17107),
.A2(n_3324),
.B(n_3325),
.Y(n_17264)
);

O2A1O1Ixp33_ASAP7_75t_L g17265 ( 
.A1(n_17154),
.A2(n_3327),
.B(n_3325),
.C(n_3326),
.Y(n_17265)
);

AOI221xp5_ASAP7_75t_L g17266 ( 
.A1(n_17130),
.A2(n_3329),
.B1(n_3327),
.B2(n_3328),
.C(n_3330),
.Y(n_17266)
);

OAI32xp33_ASAP7_75t_L g17267 ( 
.A1(n_17155),
.A2(n_3330),
.A3(n_3328),
.B1(n_3329),
.B2(n_3331),
.Y(n_17267)
);

AOI21xp5_ASAP7_75t_L g17268 ( 
.A1(n_17130),
.A2(n_3332),
.B(n_3333),
.Y(n_17268)
);

INVx1_ASAP7_75t_L g17269 ( 
.A(n_17122),
.Y(n_17269)
);

AOI21xp5_ASAP7_75t_L g17270 ( 
.A1(n_17128),
.A2(n_3332),
.B(n_3333),
.Y(n_17270)
);

OAI22x1_ASAP7_75t_L g17271 ( 
.A1(n_17136),
.A2(n_3336),
.B1(n_3334),
.B2(n_3335),
.Y(n_17271)
);

NAND2xp5_ASAP7_75t_L g17272 ( 
.A(n_17103),
.B(n_3334),
.Y(n_17272)
);

OAI221xp5_ASAP7_75t_L g17273 ( 
.A1(n_17106),
.A2(n_3338),
.B1(n_3335),
.B2(n_3337),
.C(n_3339),
.Y(n_17273)
);

OAI211xp5_ASAP7_75t_SL g17274 ( 
.A1(n_17138),
.A2(n_3339),
.B(n_3337),
.C(n_3338),
.Y(n_17274)
);

OAI322xp33_ASAP7_75t_L g17275 ( 
.A1(n_17170),
.A2(n_3345),
.A3(n_3344),
.B1(n_3342),
.B2(n_3340),
.C1(n_3341),
.C2(n_3343),
.Y(n_17275)
);

AOI21xp5_ASAP7_75t_L g17276 ( 
.A1(n_17088),
.A2(n_3341),
.B(n_3342),
.Y(n_17276)
);

OAI321xp33_ASAP7_75t_L g17277 ( 
.A1(n_17073),
.A2(n_3345),
.A3(n_3347),
.B1(n_3343),
.B2(n_3344),
.C(n_3346),
.Y(n_17277)
);

AOI322xp5_ASAP7_75t_L g17278 ( 
.A1(n_17085),
.A2(n_3352),
.A3(n_3351),
.B1(n_3349),
.B2(n_3346),
.C1(n_3348),
.C2(n_3350),
.Y(n_17278)
);

NOR2xp33_ASAP7_75t_L g17279 ( 
.A(n_17178),
.B(n_3348),
.Y(n_17279)
);

NAND2xp5_ASAP7_75t_L g17280 ( 
.A(n_17149),
.B(n_3349),
.Y(n_17280)
);

OAI321xp33_ASAP7_75t_L g17281 ( 
.A1(n_17073),
.A2(n_3354),
.A3(n_3356),
.B1(n_3351),
.B2(n_3353),
.C(n_3355),
.Y(n_17281)
);

OAI211xp5_ASAP7_75t_SL g17282 ( 
.A1(n_17138),
.A2(n_3355),
.B(n_3353),
.C(n_3354),
.Y(n_17282)
);

A2O1A1Ixp33_ASAP7_75t_L g17283 ( 
.A1(n_17074),
.A2(n_3358),
.B(n_3356),
.C(n_3357),
.Y(n_17283)
);

AOI22xp5_ASAP7_75t_L g17284 ( 
.A1(n_17085),
.A2(n_3359),
.B1(n_3357),
.B2(n_3358),
.Y(n_17284)
);

AOI211x1_ASAP7_75t_L g17285 ( 
.A1(n_17087),
.A2(n_3361),
.B(n_3359),
.C(n_3360),
.Y(n_17285)
);

INVx1_ASAP7_75t_L g17286 ( 
.A(n_17149),
.Y(n_17286)
);

NAND3xp33_ASAP7_75t_SL g17287 ( 
.A(n_17070),
.B(n_3360),
.C(n_3361),
.Y(n_17287)
);

NOR2xp33_ASAP7_75t_L g17288 ( 
.A(n_17178),
.B(n_3362),
.Y(n_17288)
);

OAI21xp33_ASAP7_75t_SL g17289 ( 
.A1(n_17117),
.A2(n_3363),
.B(n_3364),
.Y(n_17289)
);

NOR4xp25_ASAP7_75t_L g17290 ( 
.A(n_17170),
.B(n_3365),
.C(n_3363),
.D(n_3364),
.Y(n_17290)
);

AND2x2_ASAP7_75t_L g17291 ( 
.A(n_17146),
.B(n_3365),
.Y(n_17291)
);

AOI211xp5_ASAP7_75t_L g17292 ( 
.A1(n_17172),
.A2(n_3368),
.B(n_3366),
.C(n_3367),
.Y(n_17292)
);

OAI221xp5_ASAP7_75t_SL g17293 ( 
.A1(n_17138),
.A2(n_3369),
.B1(n_3366),
.B2(n_3367),
.C(n_3370),
.Y(n_17293)
);

INVx1_ASAP7_75t_L g17294 ( 
.A(n_17149),
.Y(n_17294)
);

NAND3xp33_ASAP7_75t_SL g17295 ( 
.A(n_17070),
.B(n_3369),
.C(n_3370),
.Y(n_17295)
);

AOI21xp33_ASAP7_75t_L g17296 ( 
.A1(n_17088),
.A2(n_3371),
.B(n_3373),
.Y(n_17296)
);

AOI21xp5_ASAP7_75t_L g17297 ( 
.A1(n_17088),
.A2(n_3371),
.B(n_3373),
.Y(n_17297)
);

AOI21xp33_ASAP7_75t_L g17298 ( 
.A1(n_17088),
.A2(n_3374),
.B(n_3375),
.Y(n_17298)
);

AOI211xp5_ASAP7_75t_L g17299 ( 
.A1(n_17172),
.A2(n_3376),
.B(n_3374),
.C(n_3375),
.Y(n_17299)
);

AOI221xp5_ASAP7_75t_L g17300 ( 
.A1(n_17084),
.A2(n_3378),
.B1(n_3376),
.B2(n_3377),
.C(n_3380),
.Y(n_17300)
);

OAI21xp33_ASAP7_75t_L g17301 ( 
.A1(n_17138),
.A2(n_3377),
.B(n_3380),
.Y(n_17301)
);

AOI211xp5_ASAP7_75t_SL g17302 ( 
.A1(n_17109),
.A2(n_3383),
.B(n_3381),
.C(n_3382),
.Y(n_17302)
);

OAI21xp5_ASAP7_75t_SL g17303 ( 
.A1(n_17081),
.A2(n_3381),
.B(n_3382),
.Y(n_17303)
);

OAI22xp5_ASAP7_75t_L g17304 ( 
.A1(n_17174),
.A2(n_3387),
.B1(n_3385),
.B2(n_3386),
.Y(n_17304)
);

AOI21xp5_ASAP7_75t_L g17305 ( 
.A1(n_17088),
.A2(n_3385),
.B(n_3386),
.Y(n_17305)
);

NOR2xp33_ASAP7_75t_L g17306 ( 
.A(n_17178),
.B(n_3387),
.Y(n_17306)
);

NOR2xp33_ASAP7_75t_L g17307 ( 
.A(n_17178),
.B(n_3388),
.Y(n_17307)
);

AOI21xp5_ASAP7_75t_L g17308 ( 
.A1(n_17088),
.A2(n_3388),
.B(n_3389),
.Y(n_17308)
);

OAI21xp5_ASAP7_75t_SL g17309 ( 
.A1(n_17081),
.A2(n_3389),
.B(n_3390),
.Y(n_17309)
);

AOI211xp5_ASAP7_75t_L g17310 ( 
.A1(n_17172),
.A2(n_3392),
.B(n_3390),
.C(n_3391),
.Y(n_17310)
);

AOI22xp5_ASAP7_75t_L g17311 ( 
.A1(n_17085),
.A2(n_3394),
.B1(n_3391),
.B2(n_3393),
.Y(n_17311)
);

OAI221xp5_ASAP7_75t_L g17312 ( 
.A1(n_17106),
.A2(n_3395),
.B1(n_3393),
.B2(n_3394),
.C(n_3396),
.Y(n_17312)
);

INVx1_ASAP7_75t_L g17313 ( 
.A(n_17243),
.Y(n_17313)
);

OAI211xp5_ASAP7_75t_L g17314 ( 
.A1(n_17301),
.A2(n_3399),
.B(n_3396),
.C(n_3397),
.Y(n_17314)
);

INVx1_ASAP7_75t_L g17315 ( 
.A(n_17204),
.Y(n_17315)
);

NAND2xp5_ASAP7_75t_SL g17316 ( 
.A(n_17290),
.B(n_3397),
.Y(n_17316)
);

AOI211x1_ASAP7_75t_L g17317 ( 
.A1(n_17214),
.A2(n_3401),
.B(n_3399),
.C(n_3400),
.Y(n_17317)
);

NAND4xp25_ASAP7_75t_L g17318 ( 
.A(n_17239),
.B(n_3402),
.C(n_3400),
.D(n_3401),
.Y(n_17318)
);

INVx2_ASAP7_75t_L g17319 ( 
.A(n_17196),
.Y(n_17319)
);

AND4x1_ASAP7_75t_L g17320 ( 
.A(n_17302),
.B(n_3405),
.C(n_3403),
.D(n_3404),
.Y(n_17320)
);

INVx2_ASAP7_75t_L g17321 ( 
.A(n_17196),
.Y(n_17321)
);

NAND2xp5_ASAP7_75t_SL g17322 ( 
.A(n_17277),
.B(n_3405),
.Y(n_17322)
);

NOR3xp33_ASAP7_75t_SL g17323 ( 
.A(n_17194),
.B(n_3406),
.C(n_3407),
.Y(n_17323)
);

NAND2xp5_ASAP7_75t_L g17324 ( 
.A(n_17291),
.B(n_3406),
.Y(n_17324)
);

NOR2xp33_ASAP7_75t_L g17325 ( 
.A(n_17274),
.B(n_3407),
.Y(n_17325)
);

OAI21xp33_ASAP7_75t_L g17326 ( 
.A1(n_17198),
.A2(n_3408),
.B(n_3409),
.Y(n_17326)
);

AOI211xp5_ASAP7_75t_L g17327 ( 
.A1(n_17293),
.A2(n_3411),
.B(n_3408),
.C(n_3410),
.Y(n_17327)
);

AND2x2_ASAP7_75t_L g17328 ( 
.A(n_17246),
.B(n_3410),
.Y(n_17328)
);

INVxp67_ASAP7_75t_L g17329 ( 
.A(n_17229),
.Y(n_17329)
);

INVxp67_ASAP7_75t_L g17330 ( 
.A(n_17245),
.Y(n_17330)
);

NAND4xp25_ASAP7_75t_L g17331 ( 
.A(n_17223),
.B(n_3413),
.C(n_3411),
.D(n_3412),
.Y(n_17331)
);

OAI21xp33_ASAP7_75t_L g17332 ( 
.A1(n_17200),
.A2(n_3412),
.B(n_3413),
.Y(n_17332)
);

NAND2xp5_ASAP7_75t_SL g17333 ( 
.A(n_17281),
.B(n_17219),
.Y(n_17333)
);

NAND2xp5_ASAP7_75t_L g17334 ( 
.A(n_17197),
.B(n_3414),
.Y(n_17334)
);

NOR2xp33_ASAP7_75t_L g17335 ( 
.A(n_17282),
.B(n_3414),
.Y(n_17335)
);

NAND2xp5_ASAP7_75t_SL g17336 ( 
.A(n_17187),
.B(n_3415),
.Y(n_17336)
);

NAND3xp33_ASAP7_75t_L g17337 ( 
.A(n_17241),
.B(n_3415),
.C(n_3416),
.Y(n_17337)
);

NOR2xp67_ASAP7_75t_L g17338 ( 
.A(n_17289),
.B(n_3416),
.Y(n_17338)
);

NAND4xp25_ASAP7_75t_SL g17339 ( 
.A(n_17206),
.B(n_3419),
.C(n_3417),
.D(n_3418),
.Y(n_17339)
);

NOR4xp25_ASAP7_75t_L g17340 ( 
.A(n_17212),
.B(n_3420),
.C(n_3417),
.D(n_3418),
.Y(n_17340)
);

NAND2xp5_ASAP7_75t_SL g17341 ( 
.A(n_17234),
.B(n_3420),
.Y(n_17341)
);

BUFx2_ASAP7_75t_L g17342 ( 
.A(n_17245),
.Y(n_17342)
);

NAND2xp5_ASAP7_75t_L g17343 ( 
.A(n_17238),
.B(n_3421),
.Y(n_17343)
);

AOI21xp5_ASAP7_75t_L g17344 ( 
.A1(n_17248),
.A2(n_3421),
.B(n_3422),
.Y(n_17344)
);

NAND2xp5_ASAP7_75t_L g17345 ( 
.A(n_17210),
.B(n_3422),
.Y(n_17345)
);

AOI22xp5_ASAP7_75t_L g17346 ( 
.A1(n_17215),
.A2(n_3425),
.B1(n_3423),
.B2(n_3424),
.Y(n_17346)
);

AOI322xp5_ASAP7_75t_L g17347 ( 
.A1(n_17184),
.A2(n_3429),
.A3(n_3428),
.B1(n_3426),
.B2(n_3423),
.C1(n_3425),
.C2(n_3427),
.Y(n_17347)
);

NOR2xp33_ASAP7_75t_L g17348 ( 
.A(n_17217),
.B(n_3426),
.Y(n_17348)
);

AOI21xp33_ASAP7_75t_SL g17349 ( 
.A1(n_17228),
.A2(n_3427),
.B(n_3428),
.Y(n_17349)
);

NAND2xp5_ASAP7_75t_L g17350 ( 
.A(n_17283),
.B(n_17285),
.Y(n_17350)
);

HB1xp67_ASAP7_75t_L g17351 ( 
.A(n_17253),
.Y(n_17351)
);

NAND2xp5_ASAP7_75t_L g17352 ( 
.A(n_17203),
.B(n_17266),
.Y(n_17352)
);

NAND2xp5_ASAP7_75t_L g17353 ( 
.A(n_17268),
.B(n_3429),
.Y(n_17353)
);

AND2x2_ASAP7_75t_L g17354 ( 
.A(n_17244),
.B(n_3430),
.Y(n_17354)
);

INVx1_ASAP7_75t_L g17355 ( 
.A(n_17258),
.Y(n_17355)
);

AOI222xp33_ASAP7_75t_L g17356 ( 
.A1(n_17287),
.A2(n_3432),
.B1(n_3434),
.B2(n_3430),
.C1(n_3431),
.C2(n_3433),
.Y(n_17356)
);

NAND3xp33_ASAP7_75t_L g17357 ( 
.A(n_17216),
.B(n_3432),
.C(n_3433),
.Y(n_17357)
);

NAND4xp25_ASAP7_75t_L g17358 ( 
.A(n_17240),
.B(n_3436),
.C(n_3434),
.D(n_3435),
.Y(n_17358)
);

NAND2xp5_ASAP7_75t_L g17359 ( 
.A(n_17237),
.B(n_3436),
.Y(n_17359)
);

OAI21xp33_ASAP7_75t_L g17360 ( 
.A1(n_17256),
.A2(n_3437),
.B(n_3438),
.Y(n_17360)
);

INVx1_ASAP7_75t_L g17361 ( 
.A(n_17280),
.Y(n_17361)
);

NOR4xp25_ASAP7_75t_L g17362 ( 
.A(n_17235),
.B(n_3440),
.C(n_3437),
.D(n_3439),
.Y(n_17362)
);

AOI21xp5_ASAP7_75t_L g17363 ( 
.A1(n_17218),
.A2(n_3439),
.B(n_3440),
.Y(n_17363)
);

BUFx2_ASAP7_75t_L g17364 ( 
.A(n_17190),
.Y(n_17364)
);

NAND2xp5_ASAP7_75t_L g17365 ( 
.A(n_17188),
.B(n_3441),
.Y(n_17365)
);

OAI21xp5_ASAP7_75t_SL g17366 ( 
.A1(n_17303),
.A2(n_3442),
.B(n_3443),
.Y(n_17366)
);

INVx2_ASAP7_75t_L g17367 ( 
.A(n_17249),
.Y(n_17367)
);

NAND2xp33_ASAP7_75t_L g17368 ( 
.A(n_17201),
.B(n_3442),
.Y(n_17368)
);

HB1xp67_ASAP7_75t_L g17369 ( 
.A(n_17271),
.Y(n_17369)
);

NOR2xp33_ASAP7_75t_L g17370 ( 
.A(n_17211),
.B(n_3443),
.Y(n_17370)
);

NAND3xp33_ASAP7_75t_L g17371 ( 
.A(n_17292),
.B(n_3444),
.C(n_3445),
.Y(n_17371)
);

NOR3xp33_ASAP7_75t_L g17372 ( 
.A(n_17186),
.B(n_3444),
.C(n_3446),
.Y(n_17372)
);

NAND2xp5_ASAP7_75t_L g17373 ( 
.A(n_17199),
.B(n_3446),
.Y(n_17373)
);

NOR3xp33_ASAP7_75t_SL g17374 ( 
.A(n_17295),
.B(n_3447),
.C(n_3448),
.Y(n_17374)
);

INVx1_ASAP7_75t_L g17375 ( 
.A(n_17202),
.Y(n_17375)
);

XNOR2xp5_ASAP7_75t_L g17376 ( 
.A(n_17225),
.B(n_3447),
.Y(n_17376)
);

OAI211xp5_ASAP7_75t_SL g17377 ( 
.A1(n_17257),
.A2(n_3450),
.B(n_3448),
.C(n_3449),
.Y(n_17377)
);

NAND3xp33_ASAP7_75t_SL g17378 ( 
.A(n_17299),
.B(n_3450),
.C(n_3451),
.Y(n_17378)
);

INVx1_ASAP7_75t_L g17379 ( 
.A(n_17272),
.Y(n_17379)
);

AOI21xp5_ASAP7_75t_L g17380 ( 
.A1(n_17205),
.A2(n_17209),
.B(n_17221),
.Y(n_17380)
);

NOR2xp33_ASAP7_75t_L g17381 ( 
.A(n_17273),
.B(n_3451),
.Y(n_17381)
);

NOR2xp33_ASAP7_75t_L g17382 ( 
.A(n_17312),
.B(n_3452),
.Y(n_17382)
);

AND2x2_ASAP7_75t_L g17383 ( 
.A(n_17286),
.B(n_3453),
.Y(n_17383)
);

AOI221xp5_ASAP7_75t_L g17384 ( 
.A1(n_17193),
.A2(n_17251),
.B1(n_17309),
.B2(n_17261),
.C(n_17255),
.Y(n_17384)
);

NOR4xp25_ASAP7_75t_L g17385 ( 
.A(n_17269),
.B(n_3455),
.C(n_3453),
.D(n_3454),
.Y(n_17385)
);

INVx2_ASAP7_75t_L g17386 ( 
.A(n_17294),
.Y(n_17386)
);

INVx2_ASAP7_75t_L g17387 ( 
.A(n_17224),
.Y(n_17387)
);

OAI22xp5_ASAP7_75t_L g17388 ( 
.A1(n_17192),
.A2(n_3457),
.B1(n_3455),
.B2(n_3456),
.Y(n_17388)
);

INVx1_ASAP7_75t_L g17389 ( 
.A(n_17242),
.Y(n_17389)
);

NAND5xp2_ASAP7_75t_L g17390 ( 
.A(n_17247),
.B(n_3458),
.C(n_3456),
.D(n_3457),
.E(n_3459),
.Y(n_17390)
);

INVx1_ASAP7_75t_L g17391 ( 
.A(n_17252),
.Y(n_17391)
);

NAND2x1_ASAP7_75t_SL g17392 ( 
.A(n_17222),
.B(n_3458),
.Y(n_17392)
);

AO21x1_ASAP7_75t_L g17393 ( 
.A1(n_17279),
.A2(n_3459),
.B(n_3460),
.Y(n_17393)
);

NOR3xp33_ASAP7_75t_L g17394 ( 
.A(n_17189),
.B(n_3460),
.C(n_3461),
.Y(n_17394)
);

NOR3xp33_ASAP7_75t_L g17395 ( 
.A(n_17250),
.B(n_3461),
.C(n_3462),
.Y(n_17395)
);

INVx2_ASAP7_75t_L g17396 ( 
.A(n_17284),
.Y(n_17396)
);

AND2x2_ASAP7_75t_L g17397 ( 
.A(n_17288),
.B(n_3463),
.Y(n_17397)
);

NOR3xp33_ASAP7_75t_L g17398 ( 
.A(n_17213),
.B(n_3463),
.C(n_3464),
.Y(n_17398)
);

NAND2xp5_ASAP7_75t_L g17399 ( 
.A(n_17300),
.B(n_3464),
.Y(n_17399)
);

NOR4xp25_ASAP7_75t_L g17400 ( 
.A(n_17264),
.B(n_3467),
.C(n_3465),
.D(n_3466),
.Y(n_17400)
);

INVx1_ASAP7_75t_L g17401 ( 
.A(n_17306),
.Y(n_17401)
);

AOI211x1_ASAP7_75t_L g17402 ( 
.A1(n_17232),
.A2(n_3467),
.B(n_3465),
.C(n_3466),
.Y(n_17402)
);

NOR3xp33_ASAP7_75t_L g17403 ( 
.A(n_17207),
.B(n_3468),
.C(n_3469),
.Y(n_17403)
);

INVx2_ASAP7_75t_L g17404 ( 
.A(n_17311),
.Y(n_17404)
);

AOI21xp5_ASAP7_75t_L g17405 ( 
.A1(n_17262),
.A2(n_3468),
.B(n_3469),
.Y(n_17405)
);

NAND2xp5_ASAP7_75t_SL g17406 ( 
.A(n_17220),
.B(n_3470),
.Y(n_17406)
);

INVx1_ASAP7_75t_L g17407 ( 
.A(n_17307),
.Y(n_17407)
);

NOR2xp33_ASAP7_75t_L g17408 ( 
.A(n_17260),
.B(n_3470),
.Y(n_17408)
);

NAND4xp25_ASAP7_75t_SL g17409 ( 
.A(n_17310),
.B(n_3473),
.C(n_3471),
.D(n_3472),
.Y(n_17409)
);

NOR2xp33_ASAP7_75t_L g17410 ( 
.A(n_17230),
.B(n_3471),
.Y(n_17410)
);

OAI211xp5_ASAP7_75t_SL g17411 ( 
.A1(n_17263),
.A2(n_3474),
.B(n_3472),
.C(n_3473),
.Y(n_17411)
);

NAND2xp5_ASAP7_75t_L g17412 ( 
.A(n_17183),
.B(n_3474),
.Y(n_17412)
);

AOI211xp5_ASAP7_75t_SL g17413 ( 
.A1(n_17270),
.A2(n_3477),
.B(n_3475),
.C(n_3476),
.Y(n_17413)
);

INVx1_ASAP7_75t_L g17414 ( 
.A(n_17195),
.Y(n_17414)
);

NOR2x1_ASAP7_75t_L g17415 ( 
.A(n_17227),
.B(n_3475),
.Y(n_17415)
);

NAND4xp25_ASAP7_75t_L g17416 ( 
.A(n_17208),
.B(n_17254),
.C(n_17259),
.D(n_17265),
.Y(n_17416)
);

NOR2x1_ASAP7_75t_SL g17417 ( 
.A(n_17185),
.B(n_3476),
.Y(n_17417)
);

NAND2xp5_ASAP7_75t_L g17418 ( 
.A(n_17276),
.B(n_3477),
.Y(n_17418)
);

OR2x2_ASAP7_75t_L g17419 ( 
.A(n_17304),
.B(n_17297),
.Y(n_17419)
);

OAI21xp33_ASAP7_75t_SL g17420 ( 
.A1(n_17231),
.A2(n_3478),
.B(n_3479),
.Y(n_17420)
);

NOR2xp33_ASAP7_75t_SL g17421 ( 
.A(n_17275),
.B(n_3478),
.Y(n_17421)
);

NOR2x1_ASAP7_75t_SL g17422 ( 
.A(n_17226),
.B(n_3479),
.Y(n_17422)
);

NAND2xp5_ASAP7_75t_L g17423 ( 
.A(n_17305),
.B(n_3480),
.Y(n_17423)
);

AOI21xp5_ASAP7_75t_L g17424 ( 
.A1(n_17308),
.A2(n_3481),
.B(n_3482),
.Y(n_17424)
);

NAND4xp25_ASAP7_75t_SL g17425 ( 
.A(n_17296),
.B(n_3484),
.C(n_3482),
.D(n_3483),
.Y(n_17425)
);

INVx1_ASAP7_75t_L g17426 ( 
.A(n_17267),
.Y(n_17426)
);

INVx1_ASAP7_75t_L g17427 ( 
.A(n_17236),
.Y(n_17427)
);

AOI21xp33_ASAP7_75t_L g17428 ( 
.A1(n_17298),
.A2(n_3483),
.B(n_3484),
.Y(n_17428)
);

INVx1_ASAP7_75t_L g17429 ( 
.A(n_17233),
.Y(n_17429)
);

NOR3x1_ASAP7_75t_L g17430 ( 
.A(n_17191),
.B(n_3485),
.C(n_3486),
.Y(n_17430)
);

NAND2xp5_ASAP7_75t_L g17431 ( 
.A(n_17278),
.B(n_3485),
.Y(n_17431)
);

NAND2x1_ASAP7_75t_L g17432 ( 
.A(n_17248),
.B(n_3486),
.Y(n_17432)
);

AOI21xp5_ASAP7_75t_L g17433 ( 
.A1(n_17248),
.A2(n_3487),
.B(n_3488),
.Y(n_17433)
);

NAND4xp25_ASAP7_75t_SL g17434 ( 
.A(n_17206),
.B(n_3489),
.C(n_3487),
.D(n_3488),
.Y(n_17434)
);

NAND2xp5_ASAP7_75t_SL g17435 ( 
.A(n_17290),
.B(n_3489),
.Y(n_17435)
);

NOR3x1_ASAP7_75t_L g17436 ( 
.A(n_17194),
.B(n_3490),
.C(n_3491),
.Y(n_17436)
);

AND2x2_ASAP7_75t_L g17437 ( 
.A(n_17198),
.B(n_3492),
.Y(n_17437)
);

OR2x2_ASAP7_75t_L g17438 ( 
.A(n_17318),
.B(n_3493),
.Y(n_17438)
);

NAND2xp5_ASAP7_75t_SL g17439 ( 
.A(n_17362),
.B(n_3493),
.Y(n_17439)
);

INVx1_ASAP7_75t_L g17440 ( 
.A(n_17342),
.Y(n_17440)
);

AOI22xp5_ASAP7_75t_L g17441 ( 
.A1(n_17437),
.A2(n_3497),
.B1(n_3494),
.B2(n_3495),
.Y(n_17441)
);

INVx2_ASAP7_75t_L g17442 ( 
.A(n_17354),
.Y(n_17442)
);

AOI211xp5_ASAP7_75t_SL g17443 ( 
.A1(n_17351),
.A2(n_3497),
.B(n_3494),
.C(n_3495),
.Y(n_17443)
);

NOR2x1_ASAP7_75t_L g17444 ( 
.A(n_17319),
.B(n_3498),
.Y(n_17444)
);

NAND2xp5_ASAP7_75t_SL g17445 ( 
.A(n_17385),
.B(n_17340),
.Y(n_17445)
);

NOR4xp25_ASAP7_75t_L g17446 ( 
.A(n_17355),
.B(n_3500),
.C(n_3498),
.D(n_3499),
.Y(n_17446)
);

NOR2x1_ASAP7_75t_L g17447 ( 
.A(n_17321),
.B(n_3499),
.Y(n_17447)
);

OAI21xp33_ASAP7_75t_L g17448 ( 
.A1(n_17421),
.A2(n_3500),
.B(n_3501),
.Y(n_17448)
);

NAND2xp5_ASAP7_75t_L g17449 ( 
.A(n_17328),
.B(n_3501),
.Y(n_17449)
);

NOR3x1_ASAP7_75t_L g17450 ( 
.A(n_17366),
.B(n_3502),
.C(n_3503),
.Y(n_17450)
);

NOR3xp33_ASAP7_75t_L g17451 ( 
.A(n_17364),
.B(n_3502),
.C(n_3503),
.Y(n_17451)
);

INVx1_ASAP7_75t_SL g17452 ( 
.A(n_17383),
.Y(n_17452)
);

NAND4xp75_ASAP7_75t_L g17453 ( 
.A(n_17430),
.B(n_17436),
.C(n_17338),
.D(n_17393),
.Y(n_17453)
);

OAI22xp5_ASAP7_75t_L g17454 ( 
.A1(n_17346),
.A2(n_3506),
.B1(n_3504),
.B2(n_3505),
.Y(n_17454)
);

INVx1_ASAP7_75t_L g17455 ( 
.A(n_17334),
.Y(n_17455)
);

INVx1_ASAP7_75t_L g17456 ( 
.A(n_17343),
.Y(n_17456)
);

AND2x2_ASAP7_75t_L g17457 ( 
.A(n_17323),
.B(n_3504),
.Y(n_17457)
);

AND2x2_ASAP7_75t_L g17458 ( 
.A(n_17397),
.B(n_3505),
.Y(n_17458)
);

INVx1_ASAP7_75t_L g17459 ( 
.A(n_17324),
.Y(n_17459)
);

NAND5xp2_ASAP7_75t_L g17460 ( 
.A(n_17384),
.B(n_3508),
.C(n_3506),
.D(n_3507),
.E(n_3509),
.Y(n_17460)
);

INVx1_ASAP7_75t_L g17461 ( 
.A(n_17376),
.Y(n_17461)
);

NAND2xp5_ASAP7_75t_L g17462 ( 
.A(n_17347),
.B(n_3507),
.Y(n_17462)
);

NAND4xp25_ASAP7_75t_SL g17463 ( 
.A(n_17356),
.B(n_3510),
.C(n_3508),
.D(n_3509),
.Y(n_17463)
);

NAND2xp5_ASAP7_75t_L g17464 ( 
.A(n_17372),
.B(n_3511),
.Y(n_17464)
);

AOI21xp5_ASAP7_75t_L g17465 ( 
.A1(n_17336),
.A2(n_3511),
.B(n_3512),
.Y(n_17465)
);

INVx1_ASAP7_75t_L g17466 ( 
.A(n_17353),
.Y(n_17466)
);

OAI211xp5_ASAP7_75t_SL g17467 ( 
.A1(n_17368),
.A2(n_3514),
.B(n_3512),
.C(n_3513),
.Y(n_17467)
);

NOR3xp33_ASAP7_75t_L g17468 ( 
.A(n_17386),
.B(n_3514),
.C(n_3515),
.Y(n_17468)
);

NAND4xp25_ASAP7_75t_L g17469 ( 
.A(n_17327),
.B(n_3517),
.C(n_3515),
.D(n_3516),
.Y(n_17469)
);

INVx2_ASAP7_75t_L g17470 ( 
.A(n_17432),
.Y(n_17470)
);

NAND2xp5_ASAP7_75t_L g17471 ( 
.A(n_17394),
.B(n_3516),
.Y(n_17471)
);

INVx1_ASAP7_75t_L g17472 ( 
.A(n_17359),
.Y(n_17472)
);

AND2x2_ASAP7_75t_L g17473 ( 
.A(n_17374),
.B(n_3517),
.Y(n_17473)
);

NAND2xp5_ASAP7_75t_L g17474 ( 
.A(n_17326),
.B(n_3518),
.Y(n_17474)
);

NOR2xp33_ASAP7_75t_L g17475 ( 
.A(n_17411),
.B(n_3518),
.Y(n_17475)
);

NAND3xp33_ASAP7_75t_SL g17476 ( 
.A(n_17344),
.B(n_3519),
.C(n_3520),
.Y(n_17476)
);

NOR2x1_ASAP7_75t_L g17477 ( 
.A(n_17313),
.B(n_3519),
.Y(n_17477)
);

NOR2x1_ASAP7_75t_L g17478 ( 
.A(n_17358),
.B(n_3520),
.Y(n_17478)
);

NOR4xp25_ASAP7_75t_L g17479 ( 
.A(n_17330),
.B(n_3523),
.C(n_3521),
.D(n_3522),
.Y(n_17479)
);

XNOR2x1_ASAP7_75t_L g17480 ( 
.A(n_17415),
.B(n_3521),
.Y(n_17480)
);

NAND2xp5_ASAP7_75t_L g17481 ( 
.A(n_17413),
.B(n_17433),
.Y(n_17481)
);

INVx1_ASAP7_75t_L g17482 ( 
.A(n_17320),
.Y(n_17482)
);

NAND4xp25_ASAP7_75t_L g17483 ( 
.A(n_17325),
.B(n_17335),
.C(n_17317),
.D(n_17348),
.Y(n_17483)
);

NAND2xp5_ASAP7_75t_L g17484 ( 
.A(n_17363),
.B(n_3522),
.Y(n_17484)
);

A2O1A1Ixp33_ASAP7_75t_L g17485 ( 
.A1(n_17408),
.A2(n_3526),
.B(n_3523),
.C(n_3525),
.Y(n_17485)
);

NAND4xp25_ASAP7_75t_L g17486 ( 
.A(n_17402),
.B(n_3527),
.C(n_3525),
.D(n_3526),
.Y(n_17486)
);

AOI21xp5_ASAP7_75t_L g17487 ( 
.A1(n_17316),
.A2(n_3527),
.B(n_3528),
.Y(n_17487)
);

INVx1_ASAP7_75t_L g17488 ( 
.A(n_17431),
.Y(n_17488)
);

INVx1_ASAP7_75t_L g17489 ( 
.A(n_17369),
.Y(n_17489)
);

INVx3_ASAP7_75t_L g17490 ( 
.A(n_17367),
.Y(n_17490)
);

OR2x2_ASAP7_75t_L g17491 ( 
.A(n_17400),
.B(n_3528),
.Y(n_17491)
);

OR2x2_ASAP7_75t_L g17492 ( 
.A(n_17425),
.B(n_3529),
.Y(n_17492)
);

NAND4xp75_ASAP7_75t_SL g17493 ( 
.A(n_17370),
.B(n_3531),
.C(n_3529),
.D(n_3530),
.Y(n_17493)
);

INVxp67_ASAP7_75t_L g17494 ( 
.A(n_17390),
.Y(n_17494)
);

NAND5xp2_ASAP7_75t_L g17495 ( 
.A(n_17429),
.B(n_3532),
.C(n_3530),
.D(n_3531),
.E(n_3533),
.Y(n_17495)
);

INVx1_ASAP7_75t_L g17496 ( 
.A(n_17345),
.Y(n_17496)
);

NAND2xp5_ASAP7_75t_L g17497 ( 
.A(n_17398),
.B(n_3532),
.Y(n_17497)
);

OAI211xp5_ASAP7_75t_L g17498 ( 
.A1(n_17428),
.A2(n_17314),
.B(n_17360),
.C(n_17332),
.Y(n_17498)
);

OAI211xp5_ASAP7_75t_SL g17499 ( 
.A1(n_17420),
.A2(n_3535),
.B(n_3533),
.C(n_3534),
.Y(n_17499)
);

INVx1_ASAP7_75t_L g17500 ( 
.A(n_17435),
.Y(n_17500)
);

NAND2xp5_ASAP7_75t_L g17501 ( 
.A(n_17315),
.B(n_3534),
.Y(n_17501)
);

NAND2xp5_ASAP7_75t_L g17502 ( 
.A(n_17349),
.B(n_3535),
.Y(n_17502)
);

INVx1_ASAP7_75t_L g17503 ( 
.A(n_17422),
.Y(n_17503)
);

NAND2xp5_ASAP7_75t_SL g17504 ( 
.A(n_17387),
.B(n_3536),
.Y(n_17504)
);

INVx1_ASAP7_75t_L g17505 ( 
.A(n_17412),
.Y(n_17505)
);

NAND2x1_ASAP7_75t_SL g17506 ( 
.A(n_17375),
.B(n_3537),
.Y(n_17506)
);

NOR2xp33_ASAP7_75t_L g17507 ( 
.A(n_17377),
.B(n_3537),
.Y(n_17507)
);

NAND2xp5_ASAP7_75t_L g17508 ( 
.A(n_17424),
.B(n_3538),
.Y(n_17508)
);

AOI21xp5_ASAP7_75t_L g17509 ( 
.A1(n_17333),
.A2(n_3538),
.B(n_3539),
.Y(n_17509)
);

NAND3xp33_ASAP7_75t_L g17510 ( 
.A(n_17410),
.B(n_3539),
.C(n_3540),
.Y(n_17510)
);

NAND2xp5_ASAP7_75t_L g17511 ( 
.A(n_17405),
.B(n_3540),
.Y(n_17511)
);

NOR2x1_ASAP7_75t_L g17512 ( 
.A(n_17331),
.B(n_17409),
.Y(n_17512)
);

NOR3xp33_ASAP7_75t_L g17513 ( 
.A(n_17329),
.B(n_3541),
.C(n_3542),
.Y(n_17513)
);

NAND2xp5_ASAP7_75t_L g17514 ( 
.A(n_17381),
.B(n_3541),
.Y(n_17514)
);

INVx1_ASAP7_75t_L g17515 ( 
.A(n_17418),
.Y(n_17515)
);

NAND2xp5_ASAP7_75t_SL g17516 ( 
.A(n_17388),
.B(n_3542),
.Y(n_17516)
);

AOI211xp5_ASAP7_75t_SL g17517 ( 
.A1(n_17426),
.A2(n_3545),
.B(n_3543),
.C(n_3544),
.Y(n_17517)
);

NOR3xp33_ASAP7_75t_L g17518 ( 
.A(n_17427),
.B(n_3543),
.C(n_3544),
.Y(n_17518)
);

NAND4xp25_ASAP7_75t_L g17519 ( 
.A(n_17395),
.B(n_3548),
.C(n_3546),
.D(n_3547),
.Y(n_17519)
);

OAI211xp5_ASAP7_75t_SL g17520 ( 
.A1(n_17406),
.A2(n_3549),
.B(n_3546),
.C(n_3548),
.Y(n_17520)
);

NAND3xp33_ASAP7_75t_SL g17521 ( 
.A(n_17423),
.B(n_3549),
.C(n_3550),
.Y(n_17521)
);

INVx1_ASAP7_75t_L g17522 ( 
.A(n_17417),
.Y(n_17522)
);

NOR2xp67_ASAP7_75t_L g17523 ( 
.A(n_17339),
.B(n_3550),
.Y(n_17523)
);

NAND2xp5_ASAP7_75t_L g17524 ( 
.A(n_17382),
.B(n_3551),
.Y(n_17524)
);

NAND4xp25_ASAP7_75t_L g17525 ( 
.A(n_17371),
.B(n_3553),
.C(n_3551),
.D(n_3552),
.Y(n_17525)
);

NAND2xp5_ASAP7_75t_SL g17526 ( 
.A(n_17337),
.B(n_3553),
.Y(n_17526)
);

AND2x2_ASAP7_75t_L g17527 ( 
.A(n_17396),
.B(n_3554),
.Y(n_17527)
);

NAND2xp5_ASAP7_75t_L g17528 ( 
.A(n_17392),
.B(n_3554),
.Y(n_17528)
);

NOR3xp33_ASAP7_75t_L g17529 ( 
.A(n_17379),
.B(n_17391),
.C(n_17414),
.Y(n_17529)
);

NAND3xp33_ASAP7_75t_L g17530 ( 
.A(n_17403),
.B(n_3555),
.C(n_3556),
.Y(n_17530)
);

INVx1_ASAP7_75t_L g17531 ( 
.A(n_17350),
.Y(n_17531)
);

INVxp67_ASAP7_75t_SL g17532 ( 
.A(n_17322),
.Y(n_17532)
);

AOI21xp33_ASAP7_75t_SL g17533 ( 
.A1(n_17365),
.A2(n_3555),
.B(n_3556),
.Y(n_17533)
);

OAI21xp33_ASAP7_75t_L g17534 ( 
.A1(n_17352),
.A2(n_3557),
.B(n_3558),
.Y(n_17534)
);

NOR3xp33_ASAP7_75t_L g17535 ( 
.A(n_17389),
.B(n_17407),
.C(n_17401),
.Y(n_17535)
);

NAND4xp75_ASAP7_75t_L g17536 ( 
.A(n_17380),
.B(n_3560),
.C(n_3557),
.D(n_3559),
.Y(n_17536)
);

NAND3xp33_ASAP7_75t_L g17537 ( 
.A(n_17357),
.B(n_3559),
.C(n_3561),
.Y(n_17537)
);

HB1xp67_ASAP7_75t_L g17538 ( 
.A(n_17434),
.Y(n_17538)
);

NOR2xp33_ASAP7_75t_L g17539 ( 
.A(n_17378),
.B(n_3561),
.Y(n_17539)
);

OAI21xp5_ASAP7_75t_L g17540 ( 
.A1(n_17341),
.A2(n_3562),
.B(n_3563),
.Y(n_17540)
);

AOI221x1_ASAP7_75t_L g17541 ( 
.A1(n_17361),
.A2(n_3564),
.B1(n_3562),
.B2(n_3563),
.C(n_3565),
.Y(n_17541)
);

INVx1_ASAP7_75t_L g17542 ( 
.A(n_17373),
.Y(n_17542)
);

INVx1_ASAP7_75t_L g17543 ( 
.A(n_17399),
.Y(n_17543)
);

AOI31xp33_ASAP7_75t_L g17544 ( 
.A1(n_17419),
.A2(n_17404),
.A3(n_17416),
.B(n_3567),
.Y(n_17544)
);

NAND2xp5_ASAP7_75t_L g17545 ( 
.A(n_17328),
.B(n_3564),
.Y(n_17545)
);

INVxp67_ASAP7_75t_L g17546 ( 
.A(n_17390),
.Y(n_17546)
);

INVx2_ASAP7_75t_L g17547 ( 
.A(n_17354),
.Y(n_17547)
);

NAND3xp33_ASAP7_75t_L g17548 ( 
.A(n_17347),
.B(n_3566),
.C(n_3568),
.Y(n_17548)
);

INVx1_ASAP7_75t_SL g17549 ( 
.A(n_17354),
.Y(n_17549)
);

INVx1_ASAP7_75t_L g17550 ( 
.A(n_17342),
.Y(n_17550)
);

NAND2xp5_ASAP7_75t_L g17551 ( 
.A(n_17328),
.B(n_3568),
.Y(n_17551)
);

OAI22xp33_ASAP7_75t_SL g17552 ( 
.A1(n_17432),
.A2(n_3571),
.B1(n_3569),
.B2(n_3570),
.Y(n_17552)
);

INVx1_ASAP7_75t_L g17553 ( 
.A(n_17342),
.Y(n_17553)
);

INVx1_ASAP7_75t_L g17554 ( 
.A(n_17342),
.Y(n_17554)
);

INVx1_ASAP7_75t_L g17555 ( 
.A(n_17342),
.Y(n_17555)
);

AOI32xp33_ASAP7_75t_L g17556 ( 
.A1(n_17437),
.A2(n_3572),
.A3(n_3569),
.B1(n_3570),
.B2(n_3573),
.Y(n_17556)
);

INVx1_ASAP7_75t_L g17557 ( 
.A(n_17342),
.Y(n_17557)
);

NAND3xp33_ASAP7_75t_L g17558 ( 
.A(n_17347),
.B(n_3572),
.C(n_3573),
.Y(n_17558)
);

NOR2x1_ASAP7_75t_L g17559 ( 
.A(n_17444),
.B(n_3574),
.Y(n_17559)
);

NAND4xp75_ASAP7_75t_L g17560 ( 
.A(n_17477),
.B(n_3576),
.C(n_3574),
.D(n_3575),
.Y(n_17560)
);

OAI211xp5_ASAP7_75t_SL g17561 ( 
.A1(n_17448),
.A2(n_3577),
.B(n_3575),
.C(n_3576),
.Y(n_17561)
);

NAND2x1p5_ASAP7_75t_L g17562 ( 
.A(n_17447),
.B(n_3577),
.Y(n_17562)
);

NOR2x1_ASAP7_75t_L g17563 ( 
.A(n_17536),
.B(n_3578),
.Y(n_17563)
);

NOR2xp33_ASAP7_75t_L g17564 ( 
.A(n_17467),
.B(n_3578),
.Y(n_17564)
);

NOR3xp33_ASAP7_75t_L g17565 ( 
.A(n_17489),
.B(n_3579),
.C(n_3580),
.Y(n_17565)
);

OAI211xp5_ASAP7_75t_SL g17566 ( 
.A1(n_17440),
.A2(n_3581),
.B(n_3579),
.C(n_3580),
.Y(n_17566)
);

NOR2xp33_ASAP7_75t_L g17567 ( 
.A(n_17519),
.B(n_17499),
.Y(n_17567)
);

INVx1_ASAP7_75t_L g17568 ( 
.A(n_17506),
.Y(n_17568)
);

NAND5xp2_ASAP7_75t_L g17569 ( 
.A(n_17529),
.B(n_3584),
.C(n_3582),
.D(n_3583),
.E(n_3585),
.Y(n_17569)
);

NOR2x1_ASAP7_75t_SL g17570 ( 
.A(n_17476),
.B(n_3582),
.Y(n_17570)
);

NAND3xp33_ASAP7_75t_L g17571 ( 
.A(n_17556),
.B(n_3583),
.C(n_3584),
.Y(n_17571)
);

NOR2xp67_ASAP7_75t_L g17572 ( 
.A(n_17495),
.B(n_3585),
.Y(n_17572)
);

NAND2xp5_ASAP7_75t_L g17573 ( 
.A(n_17458),
.B(n_3586),
.Y(n_17573)
);

NAND2xp5_ASAP7_75t_L g17574 ( 
.A(n_17517),
.B(n_3586),
.Y(n_17574)
);

NAND2xp5_ASAP7_75t_L g17575 ( 
.A(n_17451),
.B(n_3587),
.Y(n_17575)
);

NAND2xp5_ASAP7_75t_L g17576 ( 
.A(n_17479),
.B(n_3587),
.Y(n_17576)
);

NOR3x1_ASAP7_75t_L g17577 ( 
.A(n_17453),
.B(n_3588),
.C(n_3589),
.Y(n_17577)
);

NAND3x1_ASAP7_75t_L g17578 ( 
.A(n_17528),
.B(n_3588),
.C(n_3589),
.Y(n_17578)
);

OR2x2_ASAP7_75t_L g17579 ( 
.A(n_17460),
.B(n_3591),
.Y(n_17579)
);

NAND3xp33_ASAP7_75t_SL g17580 ( 
.A(n_17509),
.B(n_17452),
.C(n_17549),
.Y(n_17580)
);

NAND3xp33_ASAP7_75t_L g17581 ( 
.A(n_17518),
.B(n_3591),
.C(n_3592),
.Y(n_17581)
);

NOR3xp33_ASAP7_75t_SL g17582 ( 
.A(n_17483),
.B(n_3592),
.C(n_3593),
.Y(n_17582)
);

AND4x1_ASAP7_75t_L g17583 ( 
.A(n_17535),
.B(n_3595),
.C(n_3593),
.D(n_3594),
.Y(n_17583)
);

NAND3xp33_ASAP7_75t_L g17584 ( 
.A(n_17510),
.B(n_3594),
.C(n_3596),
.Y(n_17584)
);

INVx1_ASAP7_75t_L g17585 ( 
.A(n_17449),
.Y(n_17585)
);

NOR2x1_ASAP7_75t_L g17586 ( 
.A(n_17470),
.B(n_17550),
.Y(n_17586)
);

NOR2xp33_ASAP7_75t_SL g17587 ( 
.A(n_17527),
.B(n_3597),
.Y(n_17587)
);

NOR2xp33_ASAP7_75t_L g17588 ( 
.A(n_17552),
.B(n_3597),
.Y(n_17588)
);

NOR2xp33_ASAP7_75t_SL g17589 ( 
.A(n_17534),
.B(n_3598),
.Y(n_17589)
);

NOR3x1_ASAP7_75t_L g17590 ( 
.A(n_17521),
.B(n_3598),
.C(n_3599),
.Y(n_17590)
);

NAND4xp75_ASAP7_75t_L g17591 ( 
.A(n_17450),
.B(n_3601),
.C(n_3599),
.D(n_3600),
.Y(n_17591)
);

OAI221xp5_ASAP7_75t_L g17592 ( 
.A1(n_17486),
.A2(n_3602),
.B1(n_3600),
.B2(n_3601),
.C(n_3603),
.Y(n_17592)
);

INVx1_ASAP7_75t_L g17593 ( 
.A(n_17545),
.Y(n_17593)
);

NOR4xp75_ASAP7_75t_L g17594 ( 
.A(n_17540),
.B(n_3606),
.C(n_3604),
.D(n_3605),
.Y(n_17594)
);

INVxp33_ASAP7_75t_L g17595 ( 
.A(n_17457),
.Y(n_17595)
);

INVx1_ASAP7_75t_L g17596 ( 
.A(n_17551),
.Y(n_17596)
);

AOI22x1_ASAP7_75t_L g17597 ( 
.A1(n_17553),
.A2(n_3607),
.B1(n_3604),
.B2(n_3606),
.Y(n_17597)
);

NAND2xp5_ASAP7_75t_SL g17598 ( 
.A(n_17446),
.B(n_3608),
.Y(n_17598)
);

NOR2xp33_ASAP7_75t_L g17599 ( 
.A(n_17525),
.B(n_3608),
.Y(n_17599)
);

AOI211xp5_ASAP7_75t_L g17600 ( 
.A1(n_17533),
.A2(n_17463),
.B(n_17520),
.C(n_17469),
.Y(n_17600)
);

NAND2xp5_ASAP7_75t_SL g17601 ( 
.A(n_17441),
.B(n_17490),
.Y(n_17601)
);

INVx1_ASAP7_75t_SL g17602 ( 
.A(n_17491),
.Y(n_17602)
);

INVx2_ASAP7_75t_SL g17603 ( 
.A(n_17480),
.Y(n_17603)
);

NOR2x1_ASAP7_75t_L g17604 ( 
.A(n_17554),
.B(n_17555),
.Y(n_17604)
);

NAND3xp33_ASAP7_75t_L g17605 ( 
.A(n_17557),
.B(n_3609),
.C(n_3610),
.Y(n_17605)
);

INVx1_ASAP7_75t_L g17606 ( 
.A(n_17492),
.Y(n_17606)
);

NOR3xp33_ASAP7_75t_L g17607 ( 
.A(n_17544),
.B(n_17490),
.C(n_17531),
.Y(n_17607)
);

AND2x2_ASAP7_75t_L g17608 ( 
.A(n_17473),
.B(n_3609),
.Y(n_17608)
);

NAND3xp33_ASAP7_75t_L g17609 ( 
.A(n_17539),
.B(n_3610),
.C(n_3611),
.Y(n_17609)
);

NOR3xp33_ASAP7_75t_L g17610 ( 
.A(n_17500),
.B(n_3611),
.C(n_3612),
.Y(n_17610)
);

INVx2_ASAP7_75t_L g17611 ( 
.A(n_17438),
.Y(n_17611)
);

NAND2xp5_ASAP7_75t_SL g17612 ( 
.A(n_17523),
.B(n_3612),
.Y(n_17612)
);

OR2x2_ASAP7_75t_L g17613 ( 
.A(n_17502),
.B(n_3613),
.Y(n_17613)
);

NAND2x1_ASAP7_75t_SL g17614 ( 
.A(n_17538),
.B(n_3613),
.Y(n_17614)
);

NAND2xp5_ASAP7_75t_L g17615 ( 
.A(n_17443),
.B(n_3614),
.Y(n_17615)
);

O2A1O1Ixp33_ASAP7_75t_L g17616 ( 
.A1(n_17445),
.A2(n_3616),
.B(n_3614),
.C(n_3615),
.Y(n_17616)
);

AOI21xp5_ASAP7_75t_L g17617 ( 
.A1(n_17439),
.A2(n_3616),
.B(n_3617),
.Y(n_17617)
);

NAND5xp2_ASAP7_75t_L g17618 ( 
.A(n_17498),
.B(n_3619),
.C(n_3617),
.D(n_3618),
.E(n_3620),
.Y(n_17618)
);

INVx1_ASAP7_75t_L g17619 ( 
.A(n_17504),
.Y(n_17619)
);

NOR3xp33_ASAP7_75t_L g17620 ( 
.A(n_17522),
.B(n_3618),
.C(n_3619),
.Y(n_17620)
);

NOR3xp33_ASAP7_75t_L g17621 ( 
.A(n_17503),
.B(n_3621),
.C(n_3622),
.Y(n_17621)
);

NOR2x1_ASAP7_75t_L g17622 ( 
.A(n_17493),
.B(n_17482),
.Y(n_17622)
);

NOR2x1_ASAP7_75t_L g17623 ( 
.A(n_17481),
.B(n_3622),
.Y(n_17623)
);

AND2x2_ASAP7_75t_L g17624 ( 
.A(n_17478),
.B(n_3623),
.Y(n_17624)
);

INVx1_ASAP7_75t_L g17625 ( 
.A(n_17474),
.Y(n_17625)
);

NAND4xp25_ASAP7_75t_L g17626 ( 
.A(n_17475),
.B(n_3625),
.C(n_3623),
.D(n_3624),
.Y(n_17626)
);

OAI22xp5_ASAP7_75t_L g17627 ( 
.A1(n_17494),
.A2(n_3626),
.B1(n_3624),
.B2(n_3625),
.Y(n_17627)
);

NAND4xp25_ASAP7_75t_L g17628 ( 
.A(n_17530),
.B(n_3628),
.C(n_3626),
.D(n_3627),
.Y(n_17628)
);

NAND3xp33_ASAP7_75t_L g17629 ( 
.A(n_17487),
.B(n_17468),
.C(n_17462),
.Y(n_17629)
);

INVx1_ASAP7_75t_L g17630 ( 
.A(n_17497),
.Y(n_17630)
);

INVx1_ASAP7_75t_L g17631 ( 
.A(n_17484),
.Y(n_17631)
);

NOR2xp67_ASAP7_75t_L g17632 ( 
.A(n_17548),
.B(n_3627),
.Y(n_17632)
);

NAND2xp5_ASAP7_75t_L g17633 ( 
.A(n_17513),
.B(n_3628),
.Y(n_17633)
);

NOR2xp33_ASAP7_75t_L g17634 ( 
.A(n_17546),
.B(n_3629),
.Y(n_17634)
);

NAND3xp33_ASAP7_75t_L g17635 ( 
.A(n_17485),
.B(n_3629),
.C(n_3630),
.Y(n_17635)
);

AOI22xp5_ASAP7_75t_SL g17636 ( 
.A1(n_17508),
.A2(n_17511),
.B1(n_17454),
.B2(n_17507),
.Y(n_17636)
);

NOR3xp33_ASAP7_75t_SL g17637 ( 
.A(n_17514),
.B(n_3630),
.C(n_3631),
.Y(n_17637)
);

NAND3xp33_ASAP7_75t_L g17638 ( 
.A(n_17537),
.B(n_3631),
.C(n_3632),
.Y(n_17638)
);

NAND2x1_ASAP7_75t_SL g17639 ( 
.A(n_17512),
.B(n_3633),
.Y(n_17639)
);

NOR4xp25_ASAP7_75t_L g17640 ( 
.A(n_17526),
.B(n_3635),
.C(n_3633),
.D(n_3634),
.Y(n_17640)
);

NAND2xp5_ASAP7_75t_L g17641 ( 
.A(n_17465),
.B(n_3634),
.Y(n_17641)
);

NAND4xp25_ASAP7_75t_SL g17642 ( 
.A(n_17558),
.B(n_3637),
.C(n_3635),
.D(n_3636),
.Y(n_17642)
);

AOI21xp5_ASAP7_75t_L g17643 ( 
.A1(n_17524),
.A2(n_3636),
.B(n_3638),
.Y(n_17643)
);

NAND2xp5_ASAP7_75t_L g17644 ( 
.A(n_17442),
.B(n_3638),
.Y(n_17644)
);

AND2x2_ASAP7_75t_SL g17645 ( 
.A(n_17547),
.B(n_3639),
.Y(n_17645)
);

AOI22xp5_ASAP7_75t_L g17646 ( 
.A1(n_17532),
.A2(n_3642),
.B1(n_3640),
.B2(n_3641),
.Y(n_17646)
);

INVx1_ASAP7_75t_L g17647 ( 
.A(n_17501),
.Y(n_17647)
);

NOR2x1_ASAP7_75t_SL g17648 ( 
.A(n_17516),
.B(n_3640),
.Y(n_17648)
);

NAND3xp33_ASAP7_75t_L g17649 ( 
.A(n_17471),
.B(n_3642),
.C(n_3643),
.Y(n_17649)
);

NOR3xp33_ASAP7_75t_L g17650 ( 
.A(n_17461),
.B(n_3643),
.C(n_3644),
.Y(n_17650)
);

NAND2xp5_ASAP7_75t_L g17651 ( 
.A(n_17472),
.B(n_3644),
.Y(n_17651)
);

AOI211x1_ASAP7_75t_L g17652 ( 
.A1(n_17464),
.A2(n_3647),
.B(n_3645),
.C(n_3646),
.Y(n_17652)
);

INVx1_ASAP7_75t_L g17653 ( 
.A(n_17459),
.Y(n_17653)
);

NOR2xp33_ASAP7_75t_L g17654 ( 
.A(n_17455),
.B(n_17456),
.Y(n_17654)
);

NOR3xp33_ASAP7_75t_L g17655 ( 
.A(n_17488),
.B(n_3645),
.C(n_3646),
.Y(n_17655)
);

NOR2xp67_ASAP7_75t_L g17656 ( 
.A(n_17496),
.B(n_3647),
.Y(n_17656)
);

INVx1_ASAP7_75t_SL g17657 ( 
.A(n_17466),
.Y(n_17657)
);

NOR3xp33_ASAP7_75t_SL g17658 ( 
.A(n_17542),
.B(n_17543),
.C(n_17515),
.Y(n_17658)
);

AND5x1_ASAP7_75t_L g17659 ( 
.A(n_17505),
.B(n_3651),
.C(n_3648),
.D(n_3650),
.E(n_3652),
.Y(n_17659)
);

HB1xp67_ASAP7_75t_L g17660 ( 
.A(n_17541),
.Y(n_17660)
);

AND2x2_ASAP7_75t_L g17661 ( 
.A(n_17457),
.B(n_3648),
.Y(n_17661)
);

NOR2xp67_ASAP7_75t_L g17662 ( 
.A(n_17495),
.B(n_3652),
.Y(n_17662)
);

NAND3xp33_ASAP7_75t_L g17663 ( 
.A(n_17556),
.B(n_3653),
.C(n_3654),
.Y(n_17663)
);

NAND2xp5_ASAP7_75t_L g17664 ( 
.A(n_17458),
.B(n_3653),
.Y(n_17664)
);

NAND3xp33_ASAP7_75t_L g17665 ( 
.A(n_17556),
.B(n_3655),
.C(n_3656),
.Y(n_17665)
);

AND2x2_ASAP7_75t_L g17666 ( 
.A(n_17457),
.B(n_3655),
.Y(n_17666)
);

INVx1_ASAP7_75t_L g17667 ( 
.A(n_17444),
.Y(n_17667)
);

NOR2x1_ASAP7_75t_L g17668 ( 
.A(n_17444),
.B(n_3656),
.Y(n_17668)
);

NOR2xp33_ASAP7_75t_L g17669 ( 
.A(n_17467),
.B(n_3657),
.Y(n_17669)
);

INVx1_ASAP7_75t_L g17670 ( 
.A(n_17444),
.Y(n_17670)
);

NAND2xp5_ASAP7_75t_L g17671 ( 
.A(n_17458),
.B(n_3657),
.Y(n_17671)
);

AOI211x1_ASAP7_75t_L g17672 ( 
.A1(n_17544),
.A2(n_3660),
.B(n_3658),
.C(n_3659),
.Y(n_17672)
);

AND2x2_ASAP7_75t_L g17673 ( 
.A(n_17457),
.B(n_3658),
.Y(n_17673)
);

NOR2xp33_ASAP7_75t_L g17674 ( 
.A(n_17467),
.B(n_3659),
.Y(n_17674)
);

NAND2xp5_ASAP7_75t_L g17675 ( 
.A(n_17458),
.B(n_3660),
.Y(n_17675)
);

NAND4xp75_ASAP7_75t_L g17676 ( 
.A(n_17477),
.B(n_3664),
.C(n_3661),
.D(n_3662),
.Y(n_17676)
);

HB1xp67_ASAP7_75t_L g17677 ( 
.A(n_17444),
.Y(n_17677)
);

NAND2xp5_ASAP7_75t_L g17678 ( 
.A(n_17458),
.B(n_3661),
.Y(n_17678)
);

NOR3x1_ASAP7_75t_L g17679 ( 
.A(n_17453),
.B(n_3662),
.C(n_3664),
.Y(n_17679)
);

NAND3xp33_ASAP7_75t_L g17680 ( 
.A(n_17556),
.B(n_3665),
.C(n_3666),
.Y(n_17680)
);

NOR3xp33_ASAP7_75t_L g17681 ( 
.A(n_17489),
.B(n_3665),
.C(n_3666),
.Y(n_17681)
);

OR2x2_ASAP7_75t_L g17682 ( 
.A(n_17618),
.B(n_3667),
.Y(n_17682)
);

NAND2xp5_ASAP7_75t_SL g17683 ( 
.A(n_17645),
.B(n_3668),
.Y(n_17683)
);

NAND2xp5_ASAP7_75t_L g17684 ( 
.A(n_17656),
.B(n_17661),
.Y(n_17684)
);

INVxp33_ASAP7_75t_SL g17685 ( 
.A(n_17634),
.Y(n_17685)
);

INVx3_ASAP7_75t_L g17686 ( 
.A(n_17562),
.Y(n_17686)
);

NOR2x1_ASAP7_75t_L g17687 ( 
.A(n_17559),
.B(n_3668),
.Y(n_17687)
);

NOR4xp75_ASAP7_75t_L g17688 ( 
.A(n_17639),
.B(n_3671),
.C(n_3669),
.D(n_3670),
.Y(n_17688)
);

INVx1_ASAP7_75t_L g17689 ( 
.A(n_17614),
.Y(n_17689)
);

NAND2xp5_ASAP7_75t_L g17690 ( 
.A(n_17666),
.B(n_3669),
.Y(n_17690)
);

NAND2xp5_ASAP7_75t_L g17691 ( 
.A(n_17673),
.B(n_3670),
.Y(n_17691)
);

NOR3xp33_ASAP7_75t_L g17692 ( 
.A(n_17580),
.B(n_3671),
.C(n_3672),
.Y(n_17692)
);

NOR2xp33_ASAP7_75t_L g17693 ( 
.A(n_17626),
.B(n_3672),
.Y(n_17693)
);

NAND2xp5_ASAP7_75t_SL g17694 ( 
.A(n_17572),
.B(n_3673),
.Y(n_17694)
);

NAND3xp33_ASAP7_75t_L g17695 ( 
.A(n_17604),
.B(n_3673),
.C(n_3674),
.Y(n_17695)
);

NOR3x1_ASAP7_75t_L g17696 ( 
.A(n_17560),
.B(n_3674),
.C(n_3675),
.Y(n_17696)
);

NAND2xp5_ASAP7_75t_L g17697 ( 
.A(n_17608),
.B(n_3675),
.Y(n_17697)
);

NOR3xp33_ASAP7_75t_SL g17698 ( 
.A(n_17612),
.B(n_3676),
.C(n_3677),
.Y(n_17698)
);

CKINVDCx20_ASAP7_75t_R g17699 ( 
.A(n_17660),
.Y(n_17699)
);

NAND2xp5_ASAP7_75t_L g17700 ( 
.A(n_17565),
.B(n_17681),
.Y(n_17700)
);

NAND4xp75_ASAP7_75t_L g17701 ( 
.A(n_17586),
.B(n_3679),
.C(n_3676),
.D(n_3678),
.Y(n_17701)
);

NOR2xp33_ASAP7_75t_L g17702 ( 
.A(n_17592),
.B(n_3679),
.Y(n_17702)
);

NAND2xp5_ASAP7_75t_L g17703 ( 
.A(n_17655),
.B(n_3680),
.Y(n_17703)
);

NOR3xp33_ASAP7_75t_L g17704 ( 
.A(n_17601),
.B(n_3680),
.C(n_3681),
.Y(n_17704)
);

O2A1O1Ixp33_ASAP7_75t_SL g17705 ( 
.A1(n_17598),
.A2(n_3683),
.B(n_3681),
.C(n_3682),
.Y(n_17705)
);

NOR3xp33_ASAP7_75t_L g17706 ( 
.A(n_17607),
.B(n_3682),
.C(n_3683),
.Y(n_17706)
);

OAI21xp33_ASAP7_75t_L g17707 ( 
.A1(n_17595),
.A2(n_3684),
.B(n_3685),
.Y(n_17707)
);

NOR2x1_ASAP7_75t_L g17708 ( 
.A(n_17668),
.B(n_3684),
.Y(n_17708)
);

AND4x1_ASAP7_75t_L g17709 ( 
.A(n_17622),
.B(n_3688),
.C(n_3686),
.D(n_3687),
.Y(n_17709)
);

NAND4xp25_ASAP7_75t_L g17710 ( 
.A(n_17672),
.B(n_17600),
.C(n_17662),
.D(n_17590),
.Y(n_17710)
);

INVx2_ASAP7_75t_L g17711 ( 
.A(n_17597),
.Y(n_17711)
);

AOI211x1_ASAP7_75t_L g17712 ( 
.A1(n_17617),
.A2(n_3688),
.B(n_3686),
.C(n_3687),
.Y(n_17712)
);

OAI21xp33_ASAP7_75t_L g17713 ( 
.A1(n_17589),
.A2(n_3689),
.B(n_3690),
.Y(n_17713)
);

AND2x2_ASAP7_75t_L g17714 ( 
.A(n_17582),
.B(n_3689),
.Y(n_17714)
);

OAI211xp5_ASAP7_75t_SL g17715 ( 
.A1(n_17658),
.A2(n_3693),
.B(n_3691),
.C(n_3692),
.Y(n_17715)
);

NOR3xp33_ASAP7_75t_SL g17716 ( 
.A(n_17642),
.B(n_3691),
.C(n_3692),
.Y(n_17716)
);

AND2x2_ASAP7_75t_L g17717 ( 
.A(n_17637),
.B(n_3693),
.Y(n_17717)
);

NAND3xp33_ASAP7_75t_L g17718 ( 
.A(n_17587),
.B(n_3694),
.C(n_3695),
.Y(n_17718)
);

NAND2xp5_ASAP7_75t_L g17719 ( 
.A(n_17623),
.B(n_3694),
.Y(n_17719)
);

NAND2xp5_ASAP7_75t_L g17720 ( 
.A(n_17620),
.B(n_3695),
.Y(n_17720)
);

NAND4xp25_ASAP7_75t_SL g17721 ( 
.A(n_17616),
.B(n_3698),
.C(n_3696),
.D(n_3697),
.Y(n_17721)
);

OR2x2_ASAP7_75t_L g17722 ( 
.A(n_17628),
.B(n_3696),
.Y(n_17722)
);

NAND2xp5_ASAP7_75t_SL g17723 ( 
.A(n_17640),
.B(n_3698),
.Y(n_17723)
);

AOI21xp5_ASAP7_75t_L g17724 ( 
.A1(n_17677),
.A2(n_3699),
.B(n_3700),
.Y(n_17724)
);

AND4x1_ASAP7_75t_L g17725 ( 
.A(n_17577),
.B(n_3701),
.C(n_3699),
.D(n_3700),
.Y(n_17725)
);

NOR2xp67_ASAP7_75t_SL g17726 ( 
.A(n_17568),
.B(n_17667),
.Y(n_17726)
);

NOR2xp67_ASAP7_75t_L g17727 ( 
.A(n_17569),
.B(n_3702),
.Y(n_17727)
);

NAND4xp25_ASAP7_75t_L g17728 ( 
.A(n_17564),
.B(n_3705),
.C(n_3703),
.D(n_3704),
.Y(n_17728)
);

OAI211xp5_ASAP7_75t_SL g17729 ( 
.A1(n_17602),
.A2(n_3706),
.B(n_3704),
.C(n_3705),
.Y(n_17729)
);

NOR2xp67_ASAP7_75t_L g17730 ( 
.A(n_17605),
.B(n_3706),
.Y(n_17730)
);

NOR2x1_ASAP7_75t_L g17731 ( 
.A(n_17676),
.B(n_3707),
.Y(n_17731)
);

INVxp33_ASAP7_75t_SL g17732 ( 
.A(n_17636),
.Y(n_17732)
);

NOR2x1_ASAP7_75t_L g17733 ( 
.A(n_17670),
.B(n_3707),
.Y(n_17733)
);

NAND3xp33_ASAP7_75t_L g17734 ( 
.A(n_17609),
.B(n_3708),
.C(n_3709),
.Y(n_17734)
);

AND5x1_ASAP7_75t_L g17735 ( 
.A(n_17567),
.B(n_3710),
.C(n_3708),
.D(n_3709),
.E(n_3711),
.Y(n_17735)
);

AND4x1_ASAP7_75t_L g17736 ( 
.A(n_17679),
.B(n_3712),
.C(n_3710),
.D(n_3711),
.Y(n_17736)
);

NAND3x1_ASAP7_75t_L g17737 ( 
.A(n_17563),
.B(n_3712),
.C(n_3713),
.Y(n_17737)
);

AND2x2_ASAP7_75t_L g17738 ( 
.A(n_17624),
.B(n_3713),
.Y(n_17738)
);

OAI21xp5_ASAP7_75t_L g17739 ( 
.A1(n_17669),
.A2(n_3714),
.B(n_3715),
.Y(n_17739)
);

NOR2xp33_ASAP7_75t_L g17740 ( 
.A(n_17573),
.B(n_17664),
.Y(n_17740)
);

OAI211xp5_ASAP7_75t_L g17741 ( 
.A1(n_17574),
.A2(n_17652),
.B(n_17615),
.C(n_17643),
.Y(n_17741)
);

NAND2xp5_ASAP7_75t_L g17742 ( 
.A(n_17621),
.B(n_3714),
.Y(n_17742)
);

OAI21xp5_ASAP7_75t_SL g17743 ( 
.A1(n_17561),
.A2(n_3715),
.B(n_3716),
.Y(n_17743)
);

NOR3xp33_ASAP7_75t_L g17744 ( 
.A(n_17653),
.B(n_3716),
.C(n_3717),
.Y(n_17744)
);

NOR2x1_ASAP7_75t_L g17745 ( 
.A(n_17591),
.B(n_3717),
.Y(n_17745)
);

NAND3xp33_ASAP7_75t_L g17746 ( 
.A(n_17649),
.B(n_3718),
.C(n_3719),
.Y(n_17746)
);

NOR2x1_ASAP7_75t_L g17747 ( 
.A(n_17576),
.B(n_3718),
.Y(n_17747)
);

NAND4xp25_ASAP7_75t_L g17748 ( 
.A(n_17674),
.B(n_17599),
.C(n_17581),
.D(n_17571),
.Y(n_17748)
);

INVx1_ASAP7_75t_L g17749 ( 
.A(n_17671),
.Y(n_17749)
);

NAND2xp5_ASAP7_75t_L g17750 ( 
.A(n_17650),
.B(n_3719),
.Y(n_17750)
);

AND5x1_ASAP7_75t_L g17751 ( 
.A(n_17588),
.B(n_3722),
.C(n_3720),
.D(n_3721),
.E(n_3723),
.Y(n_17751)
);

INVx2_ASAP7_75t_SL g17752 ( 
.A(n_17583),
.Y(n_17752)
);

NOR2x1_ASAP7_75t_L g17753 ( 
.A(n_17675),
.B(n_3720),
.Y(n_17753)
);

NAND2xp33_ASAP7_75t_L g17754 ( 
.A(n_17578),
.B(n_3722),
.Y(n_17754)
);

INVx1_ASAP7_75t_L g17755 ( 
.A(n_17678),
.Y(n_17755)
);

NAND3xp33_ASAP7_75t_SL g17756 ( 
.A(n_17657),
.B(n_3724),
.C(n_3725),
.Y(n_17756)
);

NAND2xp5_ASAP7_75t_SL g17757 ( 
.A(n_17632),
.B(n_3724),
.Y(n_17757)
);

NOR2x1_ASAP7_75t_L g17758 ( 
.A(n_17566),
.B(n_3726),
.Y(n_17758)
);

NAND3xp33_ASAP7_75t_L g17759 ( 
.A(n_17613),
.B(n_17629),
.C(n_17663),
.Y(n_17759)
);

NAND2xp5_ASAP7_75t_L g17760 ( 
.A(n_17610),
.B(n_3727),
.Y(n_17760)
);

NOR3xp33_ASAP7_75t_L g17761 ( 
.A(n_17654),
.B(n_3727),
.C(n_3728),
.Y(n_17761)
);

NOR3xp33_ASAP7_75t_L g17762 ( 
.A(n_17603),
.B(n_3728),
.C(n_3729),
.Y(n_17762)
);

INVx2_ASAP7_75t_SL g17763 ( 
.A(n_17644),
.Y(n_17763)
);

INVx3_ASAP7_75t_L g17764 ( 
.A(n_17619),
.Y(n_17764)
);

NAND4xp25_ASAP7_75t_L g17765 ( 
.A(n_17665),
.B(n_3731),
.C(n_3729),
.D(n_3730),
.Y(n_17765)
);

NAND5xp2_ASAP7_75t_L g17766 ( 
.A(n_17606),
.B(n_3733),
.C(n_3730),
.D(n_3732),
.E(n_3734),
.Y(n_17766)
);

INVx1_ASAP7_75t_L g17767 ( 
.A(n_17579),
.Y(n_17767)
);

INVx1_ASAP7_75t_L g17768 ( 
.A(n_17594),
.Y(n_17768)
);

AOI211x1_ASAP7_75t_L g17769 ( 
.A1(n_17680),
.A2(n_3735),
.B(n_3732),
.C(n_3733),
.Y(n_17769)
);

NOR3x1_ASAP7_75t_L g17770 ( 
.A(n_17584),
.B(n_3736),
.C(n_3737),
.Y(n_17770)
);

NOR2x1_ASAP7_75t_L g17771 ( 
.A(n_17635),
.B(n_3736),
.Y(n_17771)
);

AND2x2_ASAP7_75t_L g17772 ( 
.A(n_17570),
.B(n_3737),
.Y(n_17772)
);

NAND2xp5_ASAP7_75t_L g17773 ( 
.A(n_17648),
.B(n_3738),
.Y(n_17773)
);

NAND3xp33_ASAP7_75t_L g17774 ( 
.A(n_17638),
.B(n_3739),
.C(n_3740),
.Y(n_17774)
);

NAND3xp33_ASAP7_75t_L g17775 ( 
.A(n_17575),
.B(n_3739),
.C(n_3740),
.Y(n_17775)
);

OR3x1_ASAP7_75t_L g17776 ( 
.A(n_17585),
.B(n_3741),
.C(n_3742),
.Y(n_17776)
);

INVx2_ASAP7_75t_SL g17777 ( 
.A(n_17651),
.Y(n_17777)
);

NAND4xp25_ASAP7_75t_SL g17778 ( 
.A(n_17633),
.B(n_3743),
.C(n_3741),
.D(n_3742),
.Y(n_17778)
);

NOR2x1_ASAP7_75t_L g17779 ( 
.A(n_17641),
.B(n_3743),
.Y(n_17779)
);

NAND3xp33_ASAP7_75t_L g17780 ( 
.A(n_17647),
.B(n_3744),
.C(n_3745),
.Y(n_17780)
);

NOR3xp33_ASAP7_75t_L g17781 ( 
.A(n_17611),
.B(n_17596),
.C(n_17593),
.Y(n_17781)
);

AND2x4_ASAP7_75t_L g17782 ( 
.A(n_17659),
.B(n_3744),
.Y(n_17782)
);

NAND3xp33_ASAP7_75t_SL g17783 ( 
.A(n_17625),
.B(n_3745),
.C(n_3746),
.Y(n_17783)
);

NAND4xp25_ASAP7_75t_L g17784 ( 
.A(n_17630),
.B(n_3748),
.C(n_3746),
.D(n_3747),
.Y(n_17784)
);

NOR2x1_ASAP7_75t_L g17785 ( 
.A(n_17627),
.B(n_3747),
.Y(n_17785)
);

AOI211x1_ASAP7_75t_L g17786 ( 
.A1(n_17631),
.A2(n_3750),
.B(n_3748),
.C(n_3749),
.Y(n_17786)
);

INVx1_ASAP7_75t_L g17787 ( 
.A(n_17646),
.Y(n_17787)
);

NOR4xp75_ASAP7_75t_L g17788 ( 
.A(n_17639),
.B(n_3751),
.C(n_3749),
.D(n_3750),
.Y(n_17788)
);

AND2x2_ASAP7_75t_L g17789 ( 
.A(n_17661),
.B(n_3751),
.Y(n_17789)
);

NOR3x1_ASAP7_75t_L g17790 ( 
.A(n_17560),
.B(n_3752),
.C(n_3753),
.Y(n_17790)
);

NOR2x1p5_ASAP7_75t_L g17791 ( 
.A(n_17591),
.B(n_3753),
.Y(n_17791)
);

NOR3xp33_ASAP7_75t_L g17792 ( 
.A(n_17580),
.B(n_3754),
.C(n_3755),
.Y(n_17792)
);

INVx2_ASAP7_75t_SL g17793 ( 
.A(n_17614),
.Y(n_17793)
);

NOR3xp33_ASAP7_75t_L g17794 ( 
.A(n_17580),
.B(n_3754),
.C(n_3755),
.Y(n_17794)
);

AOI221x1_ASAP7_75t_L g17795 ( 
.A1(n_17607),
.A2(n_3758),
.B1(n_3756),
.B2(n_3757),
.C(n_3759),
.Y(n_17795)
);

NOR3xp33_ASAP7_75t_L g17796 ( 
.A(n_17580),
.B(n_3756),
.C(n_3757),
.Y(n_17796)
);

NAND4xp75_ASAP7_75t_L g17797 ( 
.A(n_17604),
.B(n_3761),
.C(n_3758),
.D(n_3760),
.Y(n_17797)
);

INVx1_ASAP7_75t_L g17798 ( 
.A(n_17614),
.Y(n_17798)
);

AND2x2_ASAP7_75t_L g17799 ( 
.A(n_17661),
.B(n_3760),
.Y(n_17799)
);

NOR2xp33_ASAP7_75t_L g17800 ( 
.A(n_17626),
.B(n_3761),
.Y(n_17800)
);

OAI21xp5_ASAP7_75t_L g17801 ( 
.A1(n_17604),
.A2(n_3762),
.B(n_3763),
.Y(n_17801)
);

NOR3xp33_ASAP7_75t_L g17802 ( 
.A(n_17580),
.B(n_3762),
.C(n_3763),
.Y(n_17802)
);

NAND4xp75_ASAP7_75t_L g17803 ( 
.A(n_17604),
.B(n_3766),
.C(n_3764),
.D(n_3765),
.Y(n_17803)
);

NAND4xp25_ASAP7_75t_L g17804 ( 
.A(n_17634),
.B(n_3766),
.C(n_3764),
.D(n_3765),
.Y(n_17804)
);

AND4x1_ASAP7_75t_L g17805 ( 
.A(n_17634),
.B(n_3769),
.C(n_3767),
.D(n_3768),
.Y(n_17805)
);

NAND2xp5_ASAP7_75t_L g17806 ( 
.A(n_17645),
.B(n_3767),
.Y(n_17806)
);

NAND3xp33_ASAP7_75t_L g17807 ( 
.A(n_17634),
.B(n_3768),
.C(n_3769),
.Y(n_17807)
);

NAND4xp75_ASAP7_75t_L g17808 ( 
.A(n_17604),
.B(n_3772),
.C(n_3770),
.D(n_3771),
.Y(n_17808)
);

NOR2x1_ASAP7_75t_L g17809 ( 
.A(n_17559),
.B(n_3772),
.Y(n_17809)
);

NAND2x1p5_ASAP7_75t_L g17810 ( 
.A(n_17559),
.B(n_3770),
.Y(n_17810)
);

AND2x2_ASAP7_75t_SL g17811 ( 
.A(n_17634),
.B(n_3773),
.Y(n_17811)
);

NOR2xp67_ASAP7_75t_L g17812 ( 
.A(n_17569),
.B(n_3774),
.Y(n_17812)
);

NAND5xp2_ASAP7_75t_L g17813 ( 
.A(n_17600),
.B(n_3775),
.C(n_3773),
.D(n_3774),
.E(n_3776),
.Y(n_17813)
);

INVx1_ASAP7_75t_SL g17814 ( 
.A(n_17614),
.Y(n_17814)
);

O2A1O1Ixp33_ASAP7_75t_L g17815 ( 
.A1(n_17660),
.A2(n_3778),
.B(n_3776),
.C(n_3777),
.Y(n_17815)
);

OAI211xp5_ASAP7_75t_L g17816 ( 
.A1(n_17614),
.A2(n_3779),
.B(n_3780),
.C(n_3778),
.Y(n_17816)
);

NAND4xp25_ASAP7_75t_L g17817 ( 
.A(n_17634),
.B(n_3781),
.C(n_3777),
.D(n_3780),
.Y(n_17817)
);

NAND4xp75_ASAP7_75t_L g17818 ( 
.A(n_17604),
.B(n_3783),
.C(n_3781),
.D(n_3782),
.Y(n_17818)
);

AOI21xp33_ASAP7_75t_SL g17819 ( 
.A1(n_17562),
.A2(n_3782),
.B(n_3784),
.Y(n_17819)
);

AND2x2_ASAP7_75t_L g17820 ( 
.A(n_17661),
.B(n_3784),
.Y(n_17820)
);

NOR3xp33_ASAP7_75t_L g17821 ( 
.A(n_17580),
.B(n_3785),
.C(n_3786),
.Y(n_17821)
);

AOI21xp5_ASAP7_75t_L g17822 ( 
.A1(n_17612),
.A2(n_3785),
.B(n_3786),
.Y(n_17822)
);

NOR2x1_ASAP7_75t_L g17823 ( 
.A(n_17559),
.B(n_3788),
.Y(n_17823)
);

NAND4xp25_ASAP7_75t_L g17824 ( 
.A(n_17634),
.B(n_3791),
.C(n_3787),
.D(n_3789),
.Y(n_17824)
);

NAND2xp5_ASAP7_75t_L g17825 ( 
.A(n_17645),
.B(n_3791),
.Y(n_17825)
);

NOR2x1_ASAP7_75t_L g17826 ( 
.A(n_17559),
.B(n_3792),
.Y(n_17826)
);

INVx1_ASAP7_75t_L g17827 ( 
.A(n_17614),
.Y(n_17827)
);

NOR2x1_ASAP7_75t_L g17828 ( 
.A(n_17559),
.B(n_3792),
.Y(n_17828)
);

AND2x2_ASAP7_75t_L g17829 ( 
.A(n_17661),
.B(n_3789),
.Y(n_17829)
);

NOR3xp33_ASAP7_75t_L g17830 ( 
.A(n_17580),
.B(n_3793),
.C(n_3794),
.Y(n_17830)
);

NOR3xp33_ASAP7_75t_L g17831 ( 
.A(n_17580),
.B(n_3793),
.C(n_3794),
.Y(n_17831)
);

AOI211xp5_ASAP7_75t_L g17832 ( 
.A1(n_17592),
.A2(n_3797),
.B(n_3795),
.C(n_3796),
.Y(n_17832)
);

NOR2xp33_ASAP7_75t_L g17833 ( 
.A(n_17626),
.B(n_4575),
.Y(n_17833)
);

NOR2x1_ASAP7_75t_L g17834 ( 
.A(n_17559),
.B(n_3798),
.Y(n_17834)
);

NOR2x1_ASAP7_75t_L g17835 ( 
.A(n_17559),
.B(n_3798),
.Y(n_17835)
);

NAND4xp25_ASAP7_75t_L g17836 ( 
.A(n_17634),
.B(n_3800),
.C(n_3795),
.D(n_3799),
.Y(n_17836)
);

NOR3xp33_ASAP7_75t_L g17837 ( 
.A(n_17580),
.B(n_3799),
.C(n_3800),
.Y(n_17837)
);

NOR3xp33_ASAP7_75t_L g17838 ( 
.A(n_17580),
.B(n_3801),
.C(n_3802),
.Y(n_17838)
);

NOR2xp67_ASAP7_75t_L g17839 ( 
.A(n_17569),
.B(n_3802),
.Y(n_17839)
);

NAND3xp33_ASAP7_75t_L g17840 ( 
.A(n_17634),
.B(n_3801),
.C(n_3803),
.Y(n_17840)
);

NOR2x1_ASAP7_75t_SL g17841 ( 
.A(n_17560),
.B(n_3805),
.Y(n_17841)
);

NOR3xp33_ASAP7_75t_SL g17842 ( 
.A(n_17580),
.B(n_3804),
.C(n_3806),
.Y(n_17842)
);

NOR3xp33_ASAP7_75t_SL g17843 ( 
.A(n_17580),
.B(n_3804),
.C(n_3806),
.Y(n_17843)
);

NOR3xp33_ASAP7_75t_L g17844 ( 
.A(n_17580),
.B(n_3807),
.C(n_3808),
.Y(n_17844)
);

NAND4xp25_ASAP7_75t_L g17845 ( 
.A(n_17634),
.B(n_3809),
.C(n_3807),
.D(n_3808),
.Y(n_17845)
);

HB1xp67_ASAP7_75t_L g17846 ( 
.A(n_17688),
.Y(n_17846)
);

AOI211xp5_ASAP7_75t_L g17847 ( 
.A1(n_17819),
.A2(n_3811),
.B(n_3809),
.C(n_3810),
.Y(n_17847)
);

NOR3xp33_ASAP7_75t_L g17848 ( 
.A(n_17764),
.B(n_3810),
.C(n_3811),
.Y(n_17848)
);

OAI22xp5_ASAP7_75t_L g17849 ( 
.A1(n_17699),
.A2(n_3814),
.B1(n_3812),
.B2(n_3813),
.Y(n_17849)
);

OAI222xp33_ASAP7_75t_L g17850 ( 
.A1(n_17726),
.A2(n_3815),
.B1(n_3817),
.B2(n_3812),
.C1(n_3814),
.C2(n_3816),
.Y(n_17850)
);

O2A1O1Ixp33_ASAP7_75t_L g17851 ( 
.A1(n_17754),
.A2(n_3826),
.B(n_3834),
.C(n_3818),
.Y(n_17851)
);

OAI21xp33_ASAP7_75t_SL g17852 ( 
.A1(n_17687),
.A2(n_3819),
.B(n_3820),
.Y(n_17852)
);

AOI22xp5_ASAP7_75t_L g17853 ( 
.A1(n_17732),
.A2(n_3821),
.B1(n_3819),
.B2(n_3820),
.Y(n_17853)
);

O2A1O1Ixp33_ASAP7_75t_SL g17854 ( 
.A1(n_17683),
.A2(n_3824),
.B(n_3822),
.C(n_3823),
.Y(n_17854)
);

INVx2_ASAP7_75t_SL g17855 ( 
.A(n_17708),
.Y(n_17855)
);

AOI222xp33_ASAP7_75t_L g17856 ( 
.A1(n_17694),
.A2(n_3825),
.B1(n_3828),
.B2(n_3823),
.C1(n_3824),
.C2(n_3827),
.Y(n_17856)
);

NOR2xp67_ASAP7_75t_SL g17857 ( 
.A(n_17686),
.B(n_3825),
.Y(n_17857)
);

XOR2x2_ASAP7_75t_L g17858 ( 
.A(n_17788),
.B(n_3827),
.Y(n_17858)
);

XOR2xp5_ASAP7_75t_L g17859 ( 
.A(n_17776),
.B(n_3828),
.Y(n_17859)
);

AOI221xp5_ASAP7_75t_SL g17860 ( 
.A1(n_17757),
.A2(n_3831),
.B1(n_3829),
.B2(n_3830),
.C(n_3832),
.Y(n_17860)
);

NOR2xp33_ASAP7_75t_L g17861 ( 
.A(n_17728),
.B(n_3830),
.Y(n_17861)
);

AOI211xp5_ASAP7_75t_L g17862 ( 
.A1(n_17816),
.A2(n_3834),
.B(n_3832),
.C(n_3833),
.Y(n_17862)
);

AOI211xp5_ASAP7_75t_SL g17863 ( 
.A1(n_17764),
.A2(n_17705),
.B(n_17741),
.C(n_17689),
.Y(n_17863)
);

AOI221xp5_ASAP7_75t_L g17864 ( 
.A1(n_17721),
.A2(n_3837),
.B1(n_3835),
.B2(n_3836),
.C(n_3838),
.Y(n_17864)
);

AOI211xp5_ASAP7_75t_L g17865 ( 
.A1(n_17715),
.A2(n_3837),
.B(n_3835),
.C(n_3836),
.Y(n_17865)
);

AOI22xp5_ASAP7_75t_L g17866 ( 
.A1(n_17727),
.A2(n_3840),
.B1(n_3838),
.B2(n_3839),
.Y(n_17866)
);

AOI221x1_ASAP7_75t_L g17867 ( 
.A1(n_17781),
.A2(n_17710),
.B1(n_17827),
.B2(n_17798),
.C(n_17692),
.Y(n_17867)
);

INVx1_ASAP7_75t_L g17868 ( 
.A(n_17733),
.Y(n_17868)
);

AOI21xp5_ASAP7_75t_L g17869 ( 
.A1(n_17773),
.A2(n_3839),
.B(n_3841),
.Y(n_17869)
);

OAI31xp33_ASAP7_75t_SL g17870 ( 
.A1(n_17809),
.A2(n_4572),
.A3(n_4573),
.B(n_4571),
.Y(n_17870)
);

AOI211xp5_ASAP7_75t_L g17871 ( 
.A1(n_17713),
.A2(n_17792),
.B(n_17796),
.C(n_17794),
.Y(n_17871)
);

OAI21xp5_ASAP7_75t_SL g17872 ( 
.A1(n_17743),
.A2(n_3842),
.B(n_3843),
.Y(n_17872)
);

INVx1_ASAP7_75t_SL g17873 ( 
.A(n_17789),
.Y(n_17873)
);

AOI222xp33_ASAP7_75t_L g17874 ( 
.A1(n_17812),
.A2(n_3844),
.B1(n_3846),
.B2(n_3842),
.C1(n_3843),
.C2(n_3845),
.Y(n_17874)
);

OAI211xp5_ASAP7_75t_SL g17875 ( 
.A1(n_17747),
.A2(n_3847),
.B(n_3844),
.C(n_3846),
.Y(n_17875)
);

O2A1O1Ixp5_ASAP7_75t_L g17876 ( 
.A1(n_17723),
.A2(n_3849),
.B(n_3847),
.C(n_3848),
.Y(n_17876)
);

AOI21xp5_ASAP7_75t_L g17877 ( 
.A1(n_17793),
.A2(n_3848),
.B(n_3849),
.Y(n_17877)
);

NAND2xp5_ASAP7_75t_L g17878 ( 
.A(n_17799),
.B(n_3850),
.Y(n_17878)
);

OAI211xp5_ASAP7_75t_L g17879 ( 
.A1(n_17739),
.A2(n_3852),
.B(n_3853),
.C(n_3851),
.Y(n_17879)
);

AOI221xp5_ASAP7_75t_L g17880 ( 
.A1(n_17769),
.A2(n_3852),
.B1(n_3850),
.B2(n_3851),
.C(n_3853),
.Y(n_17880)
);

INVx2_ASAP7_75t_L g17881 ( 
.A(n_17797),
.Y(n_17881)
);

OAI211xp5_ASAP7_75t_SL g17882 ( 
.A1(n_17814),
.A2(n_3856),
.B(n_3854),
.C(n_3855),
.Y(n_17882)
);

NAND2xp5_ASAP7_75t_L g17883 ( 
.A(n_17820),
.B(n_3855),
.Y(n_17883)
);

AOI221x1_ASAP7_75t_L g17884 ( 
.A1(n_17802),
.A2(n_3858),
.B1(n_3856),
.B2(n_3857),
.C(n_3859),
.Y(n_17884)
);

A2O1A1Ixp33_ASAP7_75t_L g17885 ( 
.A1(n_17815),
.A2(n_4579),
.B(n_4570),
.C(n_3859),
.Y(n_17885)
);

OAI21xp5_ASAP7_75t_L g17886 ( 
.A1(n_17737),
.A2(n_3857),
.B(n_3858),
.Y(n_17886)
);

AOI221xp5_ASAP7_75t_L g17887 ( 
.A1(n_17712),
.A2(n_17831),
.B1(n_17837),
.B2(n_17830),
.C(n_17821),
.Y(n_17887)
);

OAI211xp5_ASAP7_75t_SL g17888 ( 
.A1(n_17823),
.A2(n_3862),
.B(n_3860),
.C(n_3861),
.Y(n_17888)
);

AOI21xp33_ASAP7_75t_L g17889 ( 
.A1(n_17702),
.A2(n_3860),
.B(n_3861),
.Y(n_17889)
);

INVx2_ASAP7_75t_L g17890 ( 
.A(n_17803),
.Y(n_17890)
);

OAI211xp5_ASAP7_75t_SL g17891 ( 
.A1(n_17826),
.A2(n_3864),
.B(n_3862),
.C(n_3863),
.Y(n_17891)
);

HB1xp67_ASAP7_75t_L g17892 ( 
.A(n_17709),
.Y(n_17892)
);

AOI21xp5_ASAP7_75t_L g17893 ( 
.A1(n_17684),
.A2(n_3864),
.B(n_3865),
.Y(n_17893)
);

AOI211x1_ASAP7_75t_SL g17894 ( 
.A1(n_17839),
.A2(n_3867),
.B(n_3865),
.C(n_3866),
.Y(n_17894)
);

OAI211xp5_ASAP7_75t_L g17895 ( 
.A1(n_17838),
.A2(n_3868),
.B(n_3869),
.C(n_3867),
.Y(n_17895)
);

OAI21xp33_ASAP7_75t_L g17896 ( 
.A1(n_17842),
.A2(n_3866),
.B(n_3868),
.Y(n_17896)
);

AOI221xp5_ASAP7_75t_SL g17897 ( 
.A1(n_17748),
.A2(n_3872),
.B1(n_3869),
.B2(n_3870),
.C(n_3873),
.Y(n_17897)
);

NAND4xp25_ASAP7_75t_SL g17898 ( 
.A(n_17832),
.B(n_3873),
.C(n_3870),
.D(n_3872),
.Y(n_17898)
);

INVx1_ASAP7_75t_L g17899 ( 
.A(n_17738),
.Y(n_17899)
);

OAI21xp33_ASAP7_75t_SL g17900 ( 
.A1(n_17828),
.A2(n_3874),
.B(n_3875),
.Y(n_17900)
);

A2O1A1Ixp33_ASAP7_75t_L g17901 ( 
.A1(n_17693),
.A2(n_4579),
.B(n_4570),
.C(n_3876),
.Y(n_17901)
);

AOI222xp33_ASAP7_75t_L g17902 ( 
.A1(n_17730),
.A2(n_3876),
.B1(n_3878),
.B2(n_3874),
.C1(n_3875),
.C2(n_3877),
.Y(n_17902)
);

NOR2xp33_ASAP7_75t_R g17903 ( 
.A(n_17686),
.B(n_3879),
.Y(n_17903)
);

NAND3xp33_ASAP7_75t_SL g17904 ( 
.A(n_17844),
.B(n_3878),
.C(n_3879),
.Y(n_17904)
);

AOI22xp33_ASAP7_75t_L g17905 ( 
.A1(n_17782),
.A2(n_3882),
.B1(n_3880),
.B2(n_3881),
.Y(n_17905)
);

O2A1O1Ixp33_ASAP7_75t_L g17906 ( 
.A1(n_17719),
.A2(n_3890),
.B(n_3900),
.C(n_3880),
.Y(n_17906)
);

INVx1_ASAP7_75t_L g17907 ( 
.A(n_17682),
.Y(n_17907)
);

OAI21xp33_ASAP7_75t_L g17908 ( 
.A1(n_17843),
.A2(n_3883),
.B(n_3884),
.Y(n_17908)
);

AOI222xp33_ASAP7_75t_L g17909 ( 
.A1(n_17841),
.A2(n_3886),
.B1(n_3888),
.B2(n_3884),
.C1(n_3885),
.C2(n_3887),
.Y(n_17909)
);

INVxp67_ASAP7_75t_L g17910 ( 
.A(n_17829),
.Y(n_17910)
);

AOI21xp5_ASAP7_75t_L g17911 ( 
.A1(n_17772),
.A2(n_3885),
.B(n_3886),
.Y(n_17911)
);

INVx1_ASAP7_75t_L g17912 ( 
.A(n_17811),
.Y(n_17912)
);

AOI322xp5_ASAP7_75t_L g17913 ( 
.A1(n_17800),
.A2(n_3893),
.A3(n_3892),
.B1(n_3889),
.B2(n_3887),
.C1(n_3888),
.C2(n_3891),
.Y(n_17913)
);

AOI21xp5_ASAP7_75t_L g17914 ( 
.A1(n_17752),
.A2(n_3891),
.B(n_3892),
.Y(n_17914)
);

NOR2xp33_ASAP7_75t_L g17915 ( 
.A(n_17765),
.B(n_3895),
.Y(n_17915)
);

NAND2xp5_ASAP7_75t_L g17916 ( 
.A(n_17706),
.B(n_3895),
.Y(n_17916)
);

INVx1_ASAP7_75t_SL g17917 ( 
.A(n_17690),
.Y(n_17917)
);

INVx1_ASAP7_75t_L g17918 ( 
.A(n_17810),
.Y(n_17918)
);

NOR3xp33_ASAP7_75t_L g17919 ( 
.A(n_17759),
.B(n_3897),
.C(n_3898),
.Y(n_17919)
);

HB1xp67_ASAP7_75t_L g17920 ( 
.A(n_17808),
.Y(n_17920)
);

OAI221xp5_ASAP7_75t_L g17921 ( 
.A1(n_17725),
.A2(n_3899),
.B1(n_3897),
.B2(n_3898),
.C(n_3900),
.Y(n_17921)
);

OAI211xp5_ASAP7_75t_L g17922 ( 
.A1(n_17753),
.A2(n_3902),
.B(n_3903),
.C(n_3901),
.Y(n_17922)
);

OAI221xp5_ASAP7_75t_L g17923 ( 
.A1(n_17736),
.A2(n_3902),
.B1(n_3899),
.B2(n_3901),
.C(n_3903),
.Y(n_17923)
);

OAI211xp5_ASAP7_75t_SL g17924 ( 
.A1(n_17834),
.A2(n_3906),
.B(n_3904),
.C(n_3905),
.Y(n_17924)
);

AOI21xp5_ASAP7_75t_L g17925 ( 
.A1(n_17806),
.A2(n_3904),
.B(n_3905),
.Y(n_17925)
);

AOI222xp33_ASAP7_75t_L g17926 ( 
.A1(n_17782),
.A2(n_3908),
.B1(n_3910),
.B2(n_3906),
.C1(n_3907),
.C2(n_3909),
.Y(n_17926)
);

OAI221xp5_ASAP7_75t_SL g17927 ( 
.A1(n_17722),
.A2(n_3910),
.B1(n_3907),
.B2(n_3908),
.C(n_3911),
.Y(n_17927)
);

BUFx2_ASAP7_75t_L g17928 ( 
.A(n_17835),
.Y(n_17928)
);

INVx1_ASAP7_75t_L g17929 ( 
.A(n_17825),
.Y(n_17929)
);

OA22x2_ASAP7_75t_SL g17930 ( 
.A1(n_17768),
.A2(n_3913),
.B1(n_3911),
.B2(n_3912),
.Y(n_17930)
);

OA211x2_ASAP7_75t_L g17931 ( 
.A1(n_17801),
.A2(n_17778),
.B(n_17756),
.C(n_17783),
.Y(n_17931)
);

OAI211xp5_ASAP7_75t_L g17932 ( 
.A1(n_17779),
.A2(n_3915),
.B(n_3916),
.C(n_3914),
.Y(n_17932)
);

AOI211x1_ASAP7_75t_L g17933 ( 
.A1(n_17822),
.A2(n_3915),
.B(n_3912),
.C(n_3914),
.Y(n_17933)
);

AOI211xp5_ASAP7_75t_L g17934 ( 
.A1(n_17746),
.A2(n_3920),
.B(n_3917),
.C(n_3919),
.Y(n_17934)
);

AOI22xp5_ASAP7_75t_L g17935 ( 
.A1(n_17833),
.A2(n_3922),
.B1(n_3920),
.B2(n_3921),
.Y(n_17935)
);

AOI221xp5_ASAP7_75t_L g17936 ( 
.A1(n_17774),
.A2(n_3923),
.B1(n_3921),
.B2(n_3922),
.C(n_3924),
.Y(n_17936)
);

AOI22xp5_ASAP7_75t_L g17937 ( 
.A1(n_17714),
.A2(n_3925),
.B1(n_3923),
.B2(n_3924),
.Y(n_17937)
);

NOR2xp67_ASAP7_75t_L g17938 ( 
.A(n_17766),
.B(n_4572),
.Y(n_17938)
);

INVxp67_ASAP7_75t_L g17939 ( 
.A(n_17691),
.Y(n_17939)
);

NOR3xp33_ASAP7_75t_SL g17940 ( 
.A(n_17740),
.B(n_3925),
.C(n_3926),
.Y(n_17940)
);

NOR3x2_ASAP7_75t_L g17941 ( 
.A(n_17818),
.B(n_3926),
.C(n_3927),
.Y(n_17941)
);

OAI211xp5_ASAP7_75t_L g17942 ( 
.A1(n_17745),
.A2(n_3929),
.B(n_3930),
.C(n_3928),
.Y(n_17942)
);

AOI22xp5_ASAP7_75t_L g17943 ( 
.A1(n_17704),
.A2(n_3929),
.B1(n_3927),
.B2(n_3928),
.Y(n_17943)
);

AOI21xp5_ASAP7_75t_L g17944 ( 
.A1(n_17717),
.A2(n_3930),
.B(n_3931),
.Y(n_17944)
);

AOI22xp5_ASAP7_75t_L g17945 ( 
.A1(n_17685),
.A2(n_3934),
.B1(n_3932),
.B2(n_3933),
.Y(n_17945)
);

NAND5xp2_ASAP7_75t_SL g17946 ( 
.A(n_17762),
.B(n_3934),
.C(n_3936),
.D(n_3933),
.E(n_3935),
.Y(n_17946)
);

INVx1_ASAP7_75t_L g17947 ( 
.A(n_17697),
.Y(n_17947)
);

CKINVDCx20_ASAP7_75t_R g17948 ( 
.A(n_17767),
.Y(n_17948)
);

OAI221xp5_ASAP7_75t_SL g17949 ( 
.A1(n_17720),
.A2(n_3936),
.B1(n_3932),
.B2(n_3935),
.C(n_3937),
.Y(n_17949)
);

HB1xp67_ASAP7_75t_L g17950 ( 
.A(n_17701),
.Y(n_17950)
);

AND2x2_ASAP7_75t_L g17951 ( 
.A(n_17698),
.B(n_3937),
.Y(n_17951)
);

OA211x2_ASAP7_75t_L g17952 ( 
.A1(n_17707),
.A2(n_3940),
.B(n_3938),
.C(n_3939),
.Y(n_17952)
);

NAND4xp25_ASAP7_75t_L g17953 ( 
.A(n_17696),
.B(n_4583),
.C(n_4569),
.D(n_3942),
.Y(n_17953)
);

OA22x2_ASAP7_75t_L g17954 ( 
.A1(n_17795),
.A2(n_3942),
.B1(n_3939),
.B2(n_3941),
.Y(n_17954)
);

AOI221xp5_ASAP7_75t_L g17955 ( 
.A1(n_17734),
.A2(n_3944),
.B1(n_3941),
.B2(n_3943),
.C(n_3945),
.Y(n_17955)
);

AOI21xp5_ASAP7_75t_L g17956 ( 
.A1(n_17700),
.A2(n_17742),
.B(n_17750),
.Y(n_17956)
);

NAND3xp33_ASAP7_75t_L g17957 ( 
.A(n_17718),
.B(n_3944),
.C(n_3945),
.Y(n_17957)
);

OAI211xp5_ASAP7_75t_L g17958 ( 
.A1(n_17731),
.A2(n_3948),
.B(n_3949),
.C(n_3947),
.Y(n_17958)
);

AOI211xp5_ASAP7_75t_SL g17959 ( 
.A1(n_17787),
.A2(n_17755),
.B(n_17749),
.C(n_17703),
.Y(n_17959)
);

OAI211xp5_ASAP7_75t_L g17960 ( 
.A1(n_17771),
.A2(n_3948),
.B(n_3949),
.C(n_3947),
.Y(n_17960)
);

AOI222xp33_ASAP7_75t_L g17961 ( 
.A1(n_17791),
.A2(n_3951),
.B1(n_3953),
.B2(n_3946),
.C1(n_3950),
.C2(n_3952),
.Y(n_17961)
);

AOI22xp5_ASAP7_75t_L g17962 ( 
.A1(n_17729),
.A2(n_3951),
.B1(n_3946),
.B2(n_3950),
.Y(n_17962)
);

O2A1O1Ixp33_ASAP7_75t_L g17963 ( 
.A1(n_17711),
.A2(n_3960),
.B(n_3969),
.C(n_3952),
.Y(n_17963)
);

INVx2_ASAP7_75t_SL g17964 ( 
.A(n_17805),
.Y(n_17964)
);

AOI221xp5_ASAP7_75t_L g17965 ( 
.A1(n_17760),
.A2(n_17716),
.B1(n_17763),
.B2(n_17777),
.C(n_17786),
.Y(n_17965)
);

INVx1_ASAP7_75t_SL g17966 ( 
.A(n_17785),
.Y(n_17966)
);

NAND3xp33_ASAP7_75t_L g17967 ( 
.A(n_17775),
.B(n_3953),
.C(n_3954),
.Y(n_17967)
);

AOI211xp5_ASAP7_75t_L g17968 ( 
.A1(n_17695),
.A2(n_3956),
.B(n_3954),
.C(n_3955),
.Y(n_17968)
);

NOR2x1_ASAP7_75t_L g17969 ( 
.A(n_17780),
.B(n_4569),
.Y(n_17969)
);

OAI211xp5_ASAP7_75t_L g17970 ( 
.A1(n_17724),
.A2(n_3957),
.B(n_3958),
.C(n_3956),
.Y(n_17970)
);

INVx2_ASAP7_75t_L g17971 ( 
.A(n_17790),
.Y(n_17971)
);

AOI221xp5_ASAP7_75t_L g17972 ( 
.A1(n_17813),
.A2(n_3958),
.B1(n_3955),
.B2(n_3957),
.C(n_3959),
.Y(n_17972)
);

AOI221x1_ASAP7_75t_L g17973 ( 
.A1(n_17761),
.A2(n_3961),
.B1(n_3959),
.B2(n_3960),
.C(n_3962),
.Y(n_17973)
);

OAI211xp5_ASAP7_75t_SL g17974 ( 
.A1(n_17758),
.A2(n_3964),
.B(n_3961),
.C(n_3963),
.Y(n_17974)
);

AOI211xp5_ASAP7_75t_L g17975 ( 
.A1(n_17807),
.A2(n_3965),
.B(n_3963),
.C(n_3964),
.Y(n_17975)
);

NAND2xp5_ASAP7_75t_L g17976 ( 
.A(n_17857),
.B(n_17744),
.Y(n_17976)
);

NOR2x1_ASAP7_75t_L g17977 ( 
.A(n_17868),
.B(n_17928),
.Y(n_17977)
);

INVx1_ASAP7_75t_L g17978 ( 
.A(n_17954),
.Y(n_17978)
);

NAND4xp75_ASAP7_75t_L g17979 ( 
.A(n_17867),
.B(n_17770),
.C(n_17751),
.D(n_17735),
.Y(n_17979)
);

OR2x2_ASAP7_75t_L g17980 ( 
.A(n_17953),
.B(n_17840),
.Y(n_17980)
);

NAND2xp5_ASAP7_75t_L g17981 ( 
.A(n_17905),
.B(n_17804),
.Y(n_17981)
);

NOR2xp67_ASAP7_75t_L g17982 ( 
.A(n_17852),
.B(n_17817),
.Y(n_17982)
);

AO21x1_ASAP7_75t_L g17983 ( 
.A1(n_17944),
.A2(n_17824),
.B(n_17836),
.Y(n_17983)
);

NOR2x1_ASAP7_75t_L g17984 ( 
.A(n_17918),
.B(n_17845),
.Y(n_17984)
);

OR2x2_ASAP7_75t_L g17985 ( 
.A(n_17898),
.B(n_17784),
.Y(n_17985)
);

OAI21xp33_ASAP7_75t_L g17986 ( 
.A1(n_17870),
.A2(n_17908),
.B(n_17896),
.Y(n_17986)
);

OAI22xp33_ASAP7_75t_SL g17987 ( 
.A1(n_17921),
.A2(n_4566),
.B1(n_4567),
.B2(n_4565),
.Y(n_17987)
);

NAND4xp75_ASAP7_75t_L g17988 ( 
.A(n_17965),
.B(n_3968),
.C(n_3965),
.D(n_3967),
.Y(n_17988)
);

NAND2x1_ASAP7_75t_SL g17989 ( 
.A(n_17846),
.B(n_3967),
.Y(n_17989)
);

NOR3x1_ASAP7_75t_L g17990 ( 
.A(n_17942),
.B(n_4567),
.C(n_4566),
.Y(n_17990)
);

NAND2xp5_ASAP7_75t_L g17991 ( 
.A(n_17909),
.B(n_3968),
.Y(n_17991)
);

NAND2xp5_ASAP7_75t_L g17992 ( 
.A(n_17894),
.B(n_3969),
.Y(n_17992)
);

AND2x2_ASAP7_75t_L g17993 ( 
.A(n_17951),
.B(n_3970),
.Y(n_17993)
);

NAND2xp5_ASAP7_75t_L g17994 ( 
.A(n_17874),
.B(n_3971),
.Y(n_17994)
);

NAND4xp25_ASAP7_75t_L g17995 ( 
.A(n_17863),
.B(n_3973),
.C(n_3971),
.D(n_3972),
.Y(n_17995)
);

NOR3x1_ASAP7_75t_L g17996 ( 
.A(n_17958),
.B(n_4577),
.C(n_4576),
.Y(n_17996)
);

NOR2x1_ASAP7_75t_L g17997 ( 
.A(n_17912),
.B(n_17932),
.Y(n_17997)
);

NOR2x1_ASAP7_75t_L g17998 ( 
.A(n_17922),
.B(n_3974),
.Y(n_17998)
);

INVx2_ASAP7_75t_L g17999 ( 
.A(n_17930),
.Y(n_17999)
);

NAND2xp5_ASAP7_75t_L g18000 ( 
.A(n_17911),
.B(n_3974),
.Y(n_18000)
);

NOR2x1_ASAP7_75t_L g18001 ( 
.A(n_17888),
.B(n_3975),
.Y(n_18001)
);

NOR2x1_ASAP7_75t_L g18002 ( 
.A(n_17891),
.B(n_3976),
.Y(n_18002)
);

NOR2x1_ASAP7_75t_L g18003 ( 
.A(n_17924),
.B(n_3976),
.Y(n_18003)
);

AND2x2_ASAP7_75t_L g18004 ( 
.A(n_17938),
.B(n_3977),
.Y(n_18004)
);

OR2x6_ASAP7_75t_L g18005 ( 
.A(n_17855),
.B(n_3977),
.Y(n_18005)
);

INVxp33_ASAP7_75t_L g18006 ( 
.A(n_17859),
.Y(n_18006)
);

HB1xp67_ASAP7_75t_L g18007 ( 
.A(n_17903),
.Y(n_18007)
);

AND2x2_ASAP7_75t_L g18008 ( 
.A(n_17940),
.B(n_3978),
.Y(n_18008)
);

INVx2_ASAP7_75t_L g18009 ( 
.A(n_17858),
.Y(n_18009)
);

INVx2_ASAP7_75t_L g18010 ( 
.A(n_17941),
.Y(n_18010)
);

NAND2x1p5_ASAP7_75t_L g18011 ( 
.A(n_17964),
.B(n_3978),
.Y(n_18011)
);

NOR2x1_ASAP7_75t_SL g18012 ( 
.A(n_17960),
.B(n_3979),
.Y(n_18012)
);

NAND3xp33_ASAP7_75t_SL g18013 ( 
.A(n_17948),
.B(n_3980),
.C(n_3981),
.Y(n_18013)
);

NOR2xp67_ASAP7_75t_L g18014 ( 
.A(n_17900),
.B(n_3981),
.Y(n_18014)
);

NAND3xp33_ASAP7_75t_SL g18015 ( 
.A(n_17873),
.B(n_3982),
.C(n_3983),
.Y(n_18015)
);

NAND3xp33_ASAP7_75t_L g18016 ( 
.A(n_17959),
.B(n_3992),
.C(n_3982),
.Y(n_18016)
);

HB1xp67_ASAP7_75t_L g18017 ( 
.A(n_17886),
.Y(n_18017)
);

AOI22xp5_ASAP7_75t_L g18018 ( 
.A1(n_17861),
.A2(n_3987),
.B1(n_3985),
.B2(n_3986),
.Y(n_18018)
);

OR2x2_ASAP7_75t_L g18019 ( 
.A(n_17904),
.B(n_3985),
.Y(n_18019)
);

INVx1_ASAP7_75t_L g18020 ( 
.A(n_17866),
.Y(n_18020)
);

NOR3xp33_ASAP7_75t_SL g18021 ( 
.A(n_17974),
.B(n_3986),
.C(n_3987),
.Y(n_18021)
);

OAI22xp5_ASAP7_75t_L g18022 ( 
.A1(n_17943),
.A2(n_3990),
.B1(n_3988),
.B2(n_3989),
.Y(n_18022)
);

NOR2x1_ASAP7_75t_L g18023 ( 
.A(n_17875),
.B(n_3988),
.Y(n_18023)
);

INVx2_ASAP7_75t_L g18024 ( 
.A(n_17878),
.Y(n_18024)
);

NOR2xp33_ASAP7_75t_R g18025 ( 
.A(n_17946),
.B(n_3989),
.Y(n_18025)
);

NAND3xp33_ASAP7_75t_L g18026 ( 
.A(n_17902),
.B(n_4000),
.C(n_3990),
.Y(n_18026)
);

NOR3x1_ASAP7_75t_L g18027 ( 
.A(n_17923),
.B(n_4582),
.C(n_4578),
.Y(n_18027)
);

NOR2x1_ASAP7_75t_L g18028 ( 
.A(n_17967),
.B(n_17899),
.Y(n_18028)
);

AND2x2_ASAP7_75t_L g18029 ( 
.A(n_17972),
.B(n_3991),
.Y(n_18029)
);

NAND4xp75_ASAP7_75t_L g18030 ( 
.A(n_17931),
.B(n_3994),
.C(n_3991),
.D(n_3993),
.Y(n_18030)
);

OAI22xp5_ASAP7_75t_L g18031 ( 
.A1(n_17962),
.A2(n_3995),
.B1(n_3993),
.B2(n_3994),
.Y(n_18031)
);

NOR2xp67_ASAP7_75t_L g18032 ( 
.A(n_17970),
.B(n_3995),
.Y(n_18032)
);

OAI21x1_ASAP7_75t_SL g18033 ( 
.A1(n_17851),
.A2(n_4006),
.B(n_3996),
.Y(n_18033)
);

NOR3xp33_ASAP7_75t_L g18034 ( 
.A(n_17910),
.B(n_3996),
.C(n_3997),
.Y(n_18034)
);

NAND2xp5_ASAP7_75t_L g18035 ( 
.A(n_17847),
.B(n_3997),
.Y(n_18035)
);

NOR3xp33_ASAP7_75t_L g18036 ( 
.A(n_17907),
.B(n_3998),
.C(n_4001),
.Y(n_18036)
);

NOR2x1_ASAP7_75t_L g18037 ( 
.A(n_17957),
.B(n_4001),
.Y(n_18037)
);

INVx1_ASAP7_75t_SL g18038 ( 
.A(n_17883),
.Y(n_18038)
);

OAI21xp5_ASAP7_75t_L g18039 ( 
.A1(n_17876),
.A2(n_4002),
.B(n_4003),
.Y(n_18039)
);

NOR2x1_ASAP7_75t_L g18040 ( 
.A(n_17971),
.B(n_4002),
.Y(n_18040)
);

NOR2xp33_ASAP7_75t_L g18041 ( 
.A(n_17872),
.B(n_4004),
.Y(n_18041)
);

INVx1_ASAP7_75t_L g18042 ( 
.A(n_17952),
.Y(n_18042)
);

NAND4xp25_ASAP7_75t_L g18043 ( 
.A(n_17915),
.B(n_4007),
.C(n_4005),
.D(n_4006),
.Y(n_18043)
);

NAND2xp5_ASAP7_75t_SL g18044 ( 
.A(n_17864),
.B(n_4005),
.Y(n_18044)
);

OR2x2_ASAP7_75t_L g18045 ( 
.A(n_17916),
.B(n_4007),
.Y(n_18045)
);

NOR3xp33_ASAP7_75t_L g18046 ( 
.A(n_17966),
.B(n_4008),
.C(n_4009),
.Y(n_18046)
);

NOR3xp33_ASAP7_75t_L g18047 ( 
.A(n_17939),
.B(n_4009),
.C(n_4010),
.Y(n_18047)
);

INVx1_ASAP7_75t_L g18048 ( 
.A(n_17854),
.Y(n_18048)
);

NOR3xp33_ASAP7_75t_L g18049 ( 
.A(n_17947),
.B(n_17929),
.C(n_17917),
.Y(n_18049)
);

CKINVDCx5p33_ASAP7_75t_R g18050 ( 
.A(n_17920),
.Y(n_18050)
);

INVxp33_ASAP7_75t_SL g18051 ( 
.A(n_17950),
.Y(n_18051)
);

OAI22xp5_ASAP7_75t_L g18052 ( 
.A1(n_17865),
.A2(n_4012),
.B1(n_4010),
.B2(n_4011),
.Y(n_18052)
);

NAND2xp5_ASAP7_75t_L g18053 ( 
.A(n_17961),
.B(n_4011),
.Y(n_18053)
);

NOR2xp67_ASAP7_75t_L g18054 ( 
.A(n_17879),
.B(n_4012),
.Y(n_18054)
);

NAND4xp75_ASAP7_75t_L g18055 ( 
.A(n_17933),
.B(n_4015),
.C(n_4013),
.D(n_4014),
.Y(n_18055)
);

NOR2x1_ASAP7_75t_L g18056 ( 
.A(n_17881),
.B(n_4014),
.Y(n_18056)
);

AND3x4_ASAP7_75t_L g18057 ( 
.A(n_17969),
.B(n_4023),
.C(n_4015),
.Y(n_18057)
);

NOR2xp67_ASAP7_75t_L g18058 ( 
.A(n_17895),
.B(n_4016),
.Y(n_18058)
);

INVx1_ASAP7_75t_L g18059 ( 
.A(n_17892),
.Y(n_18059)
);

AND2x2_ASAP7_75t_L g18060 ( 
.A(n_17890),
.B(n_4016),
.Y(n_18060)
);

AND2x2_ASAP7_75t_L g18061 ( 
.A(n_17860),
.B(n_4017),
.Y(n_18061)
);

AND2x4_ASAP7_75t_L g18062 ( 
.A(n_17869),
.B(n_4018),
.Y(n_18062)
);

OA22x2_ASAP7_75t_L g18063 ( 
.A1(n_17884),
.A2(n_4020),
.B1(n_4018),
.B2(n_4019),
.Y(n_18063)
);

INVxp33_ASAP7_75t_SL g18064 ( 
.A(n_17956),
.Y(n_18064)
);

NOR2x1_ASAP7_75t_L g18065 ( 
.A(n_17882),
.B(n_4019),
.Y(n_18065)
);

INVx2_ASAP7_75t_L g18066 ( 
.A(n_17853),
.Y(n_18066)
);

NOR2x1_ASAP7_75t_L g18067 ( 
.A(n_17901),
.B(n_4020),
.Y(n_18067)
);

NOR2x1_ASAP7_75t_L g18068 ( 
.A(n_17906),
.B(n_4021),
.Y(n_18068)
);

NOR2x1p5_ASAP7_75t_L g18069 ( 
.A(n_17871),
.B(n_4021),
.Y(n_18069)
);

XOR2x2_ASAP7_75t_L g18070 ( 
.A(n_17979),
.B(n_17862),
.Y(n_18070)
);

NOR2x1_ASAP7_75t_L g18071 ( 
.A(n_18040),
.B(n_17877),
.Y(n_18071)
);

INVx2_ASAP7_75t_SL g18072 ( 
.A(n_17989),
.Y(n_18072)
);

INVx1_ASAP7_75t_L g18073 ( 
.A(n_18063),
.Y(n_18073)
);

OAI21xp5_ASAP7_75t_L g18074 ( 
.A1(n_17977),
.A2(n_17885),
.B(n_17887),
.Y(n_18074)
);

NOR2xp67_ASAP7_75t_L g18075 ( 
.A(n_17992),
.B(n_17925),
.Y(n_18075)
);

INVx1_ASAP7_75t_L g18076 ( 
.A(n_18056),
.Y(n_18076)
);

INVx1_ASAP7_75t_L g18077 ( 
.A(n_17993),
.Y(n_18077)
);

INVx1_ASAP7_75t_L g18078 ( 
.A(n_18060),
.Y(n_18078)
);

NOR2x1_ASAP7_75t_L g18079 ( 
.A(n_17995),
.B(n_17914),
.Y(n_18079)
);

NOR2x1_ASAP7_75t_L g18080 ( 
.A(n_18016),
.B(n_17893),
.Y(n_18080)
);

NOR2x1_ASAP7_75t_L g18081 ( 
.A(n_18030),
.B(n_17963),
.Y(n_18081)
);

INVx2_ASAP7_75t_L g18082 ( 
.A(n_18005),
.Y(n_18082)
);

NOR2x1_ASAP7_75t_L g18083 ( 
.A(n_17988),
.B(n_17850),
.Y(n_18083)
);

AND2x4_ASAP7_75t_L g18084 ( 
.A(n_18014),
.B(n_17919),
.Y(n_18084)
);

NAND2xp5_ASAP7_75t_L g18085 ( 
.A(n_18004),
.B(n_17968),
.Y(n_18085)
);

AOI22xp5_ASAP7_75t_L g18086 ( 
.A1(n_18051),
.A2(n_17880),
.B1(n_17936),
.B2(n_17955),
.Y(n_18086)
);

XNOR2xp5_ASAP7_75t_L g18087 ( 
.A(n_18057),
.B(n_17934),
.Y(n_18087)
);

NAND2x1p5_ASAP7_75t_L g18088 ( 
.A(n_18042),
.B(n_17937),
.Y(n_18088)
);

OR2x2_ASAP7_75t_L g18089 ( 
.A(n_18013),
.B(n_18015),
.Y(n_18089)
);

NAND4xp75_ASAP7_75t_L g18090 ( 
.A(n_17997),
.B(n_17973),
.C(n_17889),
.D(n_17897),
.Y(n_18090)
);

OR2x2_ASAP7_75t_L g18091 ( 
.A(n_18043),
.B(n_17927),
.Y(n_18091)
);

INVx1_ASAP7_75t_L g18092 ( 
.A(n_18069),
.Y(n_18092)
);

INVx2_ASAP7_75t_L g18093 ( 
.A(n_18005),
.Y(n_18093)
);

XOR2x2_ASAP7_75t_L g18094 ( 
.A(n_18055),
.B(n_17975),
.Y(n_18094)
);

AND2x4_ASAP7_75t_L g18095 ( 
.A(n_17982),
.B(n_17848),
.Y(n_18095)
);

NAND2x1p5_ASAP7_75t_L g18096 ( 
.A(n_17999),
.B(n_17935),
.Y(n_18096)
);

NOR2x1p5_ASAP7_75t_L g18097 ( 
.A(n_17991),
.B(n_17926),
.Y(n_18097)
);

NOR2xp33_ASAP7_75t_L g18098 ( 
.A(n_17987),
.B(n_17949),
.Y(n_18098)
);

INVx1_ASAP7_75t_L g18099 ( 
.A(n_18045),
.Y(n_18099)
);

OR2x2_ASAP7_75t_L g18100 ( 
.A(n_17994),
.B(n_17849),
.Y(n_18100)
);

NAND4xp25_ASAP7_75t_L g18101 ( 
.A(n_18049),
.B(n_17856),
.C(n_17913),
.D(n_17945),
.Y(n_18101)
);

NAND2xp5_ASAP7_75t_L g18102 ( 
.A(n_18008),
.B(n_4022),
.Y(n_18102)
);

NAND4xp75_ASAP7_75t_L g18103 ( 
.A(n_17984),
.B(n_4025),
.C(n_4022),
.D(n_4024),
.Y(n_18103)
);

INVx1_ASAP7_75t_L g18104 ( 
.A(n_18000),
.Y(n_18104)
);

NAND2xp5_ASAP7_75t_L g18105 ( 
.A(n_18011),
.B(n_4024),
.Y(n_18105)
);

NOR2x1_ASAP7_75t_L g18106 ( 
.A(n_17978),
.B(n_18010),
.Y(n_18106)
);

AND2x4_ASAP7_75t_L g18107 ( 
.A(n_18037),
.B(n_4026),
.Y(n_18107)
);

NAND2xp5_ASAP7_75t_L g18108 ( 
.A(n_18046),
.B(n_4026),
.Y(n_18108)
);

HB1xp67_ASAP7_75t_L g18109 ( 
.A(n_18025),
.Y(n_18109)
);

INVx1_ASAP7_75t_L g18110 ( 
.A(n_18012),
.Y(n_18110)
);

NAND4xp75_ASAP7_75t_L g18111 ( 
.A(n_18028),
.B(n_4029),
.C(n_4027),
.D(n_4028),
.Y(n_18111)
);

NAND4xp75_ASAP7_75t_L g18112 ( 
.A(n_18059),
.B(n_4031),
.C(n_4029),
.D(n_4030),
.Y(n_18112)
);

NAND2xp5_ASAP7_75t_L g18113 ( 
.A(n_18032),
.B(n_4030),
.Y(n_18113)
);

HB1xp67_ASAP7_75t_L g18114 ( 
.A(n_18054),
.Y(n_18114)
);

NOR2x1_ASAP7_75t_L g18115 ( 
.A(n_18048),
.B(n_4031),
.Y(n_18115)
);

NOR2x1_ASAP7_75t_L g18116 ( 
.A(n_17998),
.B(n_4032),
.Y(n_18116)
);

INVxp67_ASAP7_75t_SL g18117 ( 
.A(n_18053),
.Y(n_18117)
);

OAI211xp5_ASAP7_75t_L g18118 ( 
.A1(n_17986),
.A2(n_18007),
.B(n_18050),
.C(n_18017),
.Y(n_18118)
);

INVx1_ASAP7_75t_L g18119 ( 
.A(n_18033),
.Y(n_18119)
);

XOR2xp5_ASAP7_75t_L g18120 ( 
.A(n_18006),
.B(n_17985),
.Y(n_18120)
);

AOI22xp5_ASAP7_75t_L g18121 ( 
.A1(n_18041),
.A2(n_4034),
.B1(n_4035),
.B2(n_4033),
.Y(n_18121)
);

INVx2_ASAP7_75t_L g18122 ( 
.A(n_17990),
.Y(n_18122)
);

HB1xp67_ASAP7_75t_L g18123 ( 
.A(n_17996),
.Y(n_18123)
);

XNOR2xp5_ASAP7_75t_L g18124 ( 
.A(n_18023),
.B(n_4032),
.Y(n_18124)
);

INVx1_ASAP7_75t_L g18125 ( 
.A(n_18019),
.Y(n_18125)
);

XNOR2xp5_ASAP7_75t_L g18126 ( 
.A(n_18001),
.B(n_4034),
.Y(n_18126)
);

AND3x2_ASAP7_75t_L g18127 ( 
.A(n_18036),
.B(n_4035),
.C(n_4036),
.Y(n_18127)
);

INVx1_ASAP7_75t_L g18128 ( 
.A(n_18002),
.Y(n_18128)
);

NOR2xp67_ASAP7_75t_L g18129 ( 
.A(n_18026),
.B(n_4038),
.Y(n_18129)
);

XNOR2xp5_ASAP7_75t_L g18130 ( 
.A(n_18003),
.B(n_4037),
.Y(n_18130)
);

NOR3xp33_ASAP7_75t_L g18131 ( 
.A(n_18009),
.B(n_4037),
.C(n_4038),
.Y(n_18131)
);

INVx1_ASAP7_75t_SL g18132 ( 
.A(n_18062),
.Y(n_18132)
);

OAI22x1_ASAP7_75t_L g18133 ( 
.A1(n_18018),
.A2(n_4041),
.B1(n_4039),
.B2(n_4040),
.Y(n_18133)
);

INVxp33_ASAP7_75t_SL g18134 ( 
.A(n_18027),
.Y(n_18134)
);

HB1xp67_ASAP7_75t_L g18135 ( 
.A(n_18058),
.Y(n_18135)
);

AOI21xp33_ASAP7_75t_L g18136 ( 
.A1(n_17980),
.A2(n_4039),
.B(n_4040),
.Y(n_18136)
);

NOR2xp67_ASAP7_75t_L g18137 ( 
.A(n_18062),
.B(n_4042),
.Y(n_18137)
);

AND2x2_ASAP7_75t_L g18138 ( 
.A(n_18021),
.B(n_4041),
.Y(n_18138)
);

NAND4xp75_ASAP7_75t_L g18139 ( 
.A(n_18068),
.B(n_4046),
.C(n_4044),
.D(n_4045),
.Y(n_18139)
);

INVx1_ASAP7_75t_L g18140 ( 
.A(n_18102),
.Y(n_18140)
);

AND2x2_ASAP7_75t_L g18141 ( 
.A(n_18138),
.B(n_18061),
.Y(n_18141)
);

INVx1_ASAP7_75t_L g18142 ( 
.A(n_18105),
.Y(n_18142)
);

INVx1_ASAP7_75t_L g18143 ( 
.A(n_18115),
.Y(n_18143)
);

NOR2x1_ASAP7_75t_L g18144 ( 
.A(n_18076),
.B(n_18024),
.Y(n_18144)
);

INVx2_ASAP7_75t_L g18145 ( 
.A(n_18112),
.Y(n_18145)
);

NOR2x1_ASAP7_75t_L g18146 ( 
.A(n_18116),
.B(n_18067),
.Y(n_18146)
);

INVx1_ASAP7_75t_L g18147 ( 
.A(n_18139),
.Y(n_18147)
);

NAND2xp5_ASAP7_75t_L g18148 ( 
.A(n_18127),
.B(n_18137),
.Y(n_18148)
);

INVxp67_ASAP7_75t_SL g18149 ( 
.A(n_18113),
.Y(n_18149)
);

INVx1_ASAP7_75t_L g18150 ( 
.A(n_18124),
.Y(n_18150)
);

INVx2_ASAP7_75t_L g18151 ( 
.A(n_18103),
.Y(n_18151)
);

NAND2xp5_ASAP7_75t_L g18152 ( 
.A(n_18107),
.B(n_18052),
.Y(n_18152)
);

NAND2x1p5_ASAP7_75t_L g18153 ( 
.A(n_18071),
.B(n_18038),
.Y(n_18153)
);

INVx1_ASAP7_75t_L g18154 ( 
.A(n_18126),
.Y(n_18154)
);

INVx2_ASAP7_75t_L g18155 ( 
.A(n_18111),
.Y(n_18155)
);

INVxp67_ASAP7_75t_L g18156 ( 
.A(n_18107),
.Y(n_18156)
);

INVx2_ASAP7_75t_L g18157 ( 
.A(n_18133),
.Y(n_18157)
);

NAND2x1p5_ASAP7_75t_L g18158 ( 
.A(n_18072),
.B(n_18020),
.Y(n_18158)
);

NAND4xp75_ASAP7_75t_L g18159 ( 
.A(n_18106),
.B(n_18075),
.C(n_18074),
.D(n_18128),
.Y(n_18159)
);

OAI21xp33_ASAP7_75t_L g18160 ( 
.A1(n_18134),
.A2(n_18064),
.B(n_17981),
.Y(n_18160)
);

NAND4xp75_ASAP7_75t_L g18161 ( 
.A(n_18110),
.B(n_18065),
.C(n_17983),
.D(n_17976),
.Y(n_18161)
);

XNOR2x1_ASAP7_75t_L g18162 ( 
.A(n_18070),
.B(n_18066),
.Y(n_18162)
);

AND2x2_ASAP7_75t_SL g18163 ( 
.A(n_18084),
.B(n_18029),
.Y(n_18163)
);

XOR2x1_ASAP7_75t_L g18164 ( 
.A(n_18088),
.B(n_18031),
.Y(n_18164)
);

INVx2_ASAP7_75t_SL g18165 ( 
.A(n_18094),
.Y(n_18165)
);

AOI21xp33_ASAP7_75t_L g18166 ( 
.A1(n_18130),
.A2(n_18118),
.B(n_18120),
.Y(n_18166)
);

NAND2xp5_ASAP7_75t_L g18167 ( 
.A(n_18131),
.B(n_18034),
.Y(n_18167)
);

XNOR2x1_ASAP7_75t_L g18168 ( 
.A(n_18090),
.B(n_18039),
.Y(n_18168)
);

INVx1_ASAP7_75t_L g18169 ( 
.A(n_18108),
.Y(n_18169)
);

INVx1_ASAP7_75t_L g18170 ( 
.A(n_18083),
.Y(n_18170)
);

XOR2xp5_ASAP7_75t_L g18171 ( 
.A(n_18087),
.B(n_18035),
.Y(n_18171)
);

NAND2x1p5_ASAP7_75t_L g18172 ( 
.A(n_18073),
.B(n_18044),
.Y(n_18172)
);

NOR2x1_ASAP7_75t_L g18173 ( 
.A(n_18082),
.B(n_18022),
.Y(n_18173)
);

OR2x2_ASAP7_75t_L g18174 ( 
.A(n_18089),
.B(n_18047),
.Y(n_18174)
);

NAND2xp5_ASAP7_75t_L g18175 ( 
.A(n_18129),
.B(n_4045),
.Y(n_18175)
);

AOI21xp5_ASAP7_75t_SL g18176 ( 
.A1(n_18084),
.A2(n_4044),
.B(n_4046),
.Y(n_18176)
);

NAND4xp75_ASAP7_75t_L g18177 ( 
.A(n_18078),
.B(n_4049),
.C(n_4047),
.D(n_4048),
.Y(n_18177)
);

BUFx12f_ASAP7_75t_L g18178 ( 
.A(n_18095),
.Y(n_18178)
);

AOI21xp5_ASAP7_75t_SL g18179 ( 
.A1(n_18093),
.A2(n_4047),
.B(n_4048),
.Y(n_18179)
);

INVx2_ASAP7_75t_L g18180 ( 
.A(n_18097),
.Y(n_18180)
);

INVx1_ASAP7_75t_L g18181 ( 
.A(n_18081),
.Y(n_18181)
);

NAND4xp75_ASAP7_75t_L g18182 ( 
.A(n_18119),
.B(n_4051),
.C(n_4049),
.D(n_4050),
.Y(n_18182)
);

AND2x4_ASAP7_75t_L g18183 ( 
.A(n_18079),
.B(n_4051),
.Y(n_18183)
);

NAND2x1p5_ASAP7_75t_L g18184 ( 
.A(n_18132),
.B(n_4052),
.Y(n_18184)
);

NAND2xp5_ASAP7_75t_L g18185 ( 
.A(n_18121),
.B(n_4054),
.Y(n_18185)
);

XNOR2x1_ASAP7_75t_L g18186 ( 
.A(n_18096),
.B(n_4053),
.Y(n_18186)
);

XOR2xp5_ASAP7_75t_L g18187 ( 
.A(n_18109),
.B(n_4053),
.Y(n_18187)
);

NOR2xp33_ASAP7_75t_L g18188 ( 
.A(n_18101),
.B(n_4054),
.Y(n_18188)
);

INVx2_ASAP7_75t_L g18189 ( 
.A(n_18091),
.Y(n_18189)
);

BUFx3_ASAP7_75t_L g18190 ( 
.A(n_18122),
.Y(n_18190)
);

INVxp67_ASAP7_75t_SL g18191 ( 
.A(n_18123),
.Y(n_18191)
);

AOI22xp5_ASAP7_75t_L g18192 ( 
.A1(n_18098),
.A2(n_4063),
.B1(n_4071),
.B2(n_4055),
.Y(n_18192)
);

NOR2xp33_ASAP7_75t_L g18193 ( 
.A(n_18077),
.B(n_4055),
.Y(n_18193)
);

NOR2x1_ASAP7_75t_L g18194 ( 
.A(n_18092),
.B(n_4056),
.Y(n_18194)
);

XNOR2xp5_ASAP7_75t_L g18195 ( 
.A(n_18086),
.B(n_4056),
.Y(n_18195)
);

INVx1_ASAP7_75t_L g18196 ( 
.A(n_18085),
.Y(n_18196)
);

INVx1_ASAP7_75t_L g18197 ( 
.A(n_18135),
.Y(n_18197)
);

XOR2xp5_ASAP7_75t_L g18198 ( 
.A(n_18114),
.B(n_4057),
.Y(n_18198)
);

OR2x2_ASAP7_75t_L g18199 ( 
.A(n_18100),
.B(n_4057),
.Y(n_18199)
);

HB1xp67_ASAP7_75t_L g18200 ( 
.A(n_18080),
.Y(n_18200)
);

INVx1_ASAP7_75t_L g18201 ( 
.A(n_18099),
.Y(n_18201)
);

NOR2x1p5_ASAP7_75t_L g18202 ( 
.A(n_18117),
.B(n_4058),
.Y(n_18202)
);

OR2x2_ASAP7_75t_L g18203 ( 
.A(n_18125),
.B(n_4058),
.Y(n_18203)
);

INVx2_ASAP7_75t_L g18204 ( 
.A(n_18095),
.Y(n_18204)
);

AND2x2_ASAP7_75t_SL g18205 ( 
.A(n_18104),
.B(n_4059),
.Y(n_18205)
);

OAI21xp5_ASAP7_75t_L g18206 ( 
.A1(n_18136),
.A2(n_4059),
.B(n_4060),
.Y(n_18206)
);

INVx1_ASAP7_75t_L g18207 ( 
.A(n_18102),
.Y(n_18207)
);

XNOR2xp5_ASAP7_75t_L g18208 ( 
.A(n_18120),
.B(n_4060),
.Y(n_18208)
);

AOI22xp5_ASAP7_75t_L g18209 ( 
.A1(n_18134),
.A2(n_4069),
.B1(n_4079),
.B2(n_4061),
.Y(n_18209)
);

NAND3xp33_ASAP7_75t_L g18210 ( 
.A(n_18106),
.B(n_4061),
.C(n_4062),
.Y(n_18210)
);

AND2x4_ASAP7_75t_L g18211 ( 
.A(n_18137),
.B(n_4062),
.Y(n_18211)
);

INVx2_ASAP7_75t_L g18212 ( 
.A(n_18112),
.Y(n_18212)
);

AOI22xp5_ASAP7_75t_L g18213 ( 
.A1(n_18134),
.A2(n_4072),
.B1(n_4082),
.B2(n_4063),
.Y(n_18213)
);

INVx1_ASAP7_75t_L g18214 ( 
.A(n_18102),
.Y(n_18214)
);

XOR2xp5_ASAP7_75t_L g18215 ( 
.A(n_18120),
.B(n_4064),
.Y(n_18215)
);

INVx1_ASAP7_75t_L g18216 ( 
.A(n_18102),
.Y(n_18216)
);

XNOR2xp5_ASAP7_75t_L g18217 ( 
.A(n_18120),
.B(n_4065),
.Y(n_18217)
);

NOR5xp2_ASAP7_75t_L g18218 ( 
.A(n_18200),
.B(n_4067),
.C(n_4069),
.D(n_4066),
.E(n_4068),
.Y(n_18218)
);

NOR3xp33_ASAP7_75t_SL g18219 ( 
.A(n_18159),
.B(n_4065),
.C(n_4067),
.Y(n_18219)
);

AOI22xp33_ASAP7_75t_L g18220 ( 
.A1(n_18178),
.A2(n_4073),
.B1(n_4068),
.B2(n_4070),
.Y(n_18220)
);

AOI22xp5_ASAP7_75t_L g18221 ( 
.A1(n_18188),
.A2(n_4074),
.B1(n_4070),
.B2(n_4073),
.Y(n_18221)
);

NAND4xp25_ASAP7_75t_L g18222 ( 
.A(n_18166),
.B(n_4076),
.C(n_4074),
.D(n_4075),
.Y(n_18222)
);

NOR4xp25_ASAP7_75t_L g18223 ( 
.A(n_18160),
.B(n_4077),
.C(n_4075),
.D(n_4076),
.Y(n_18223)
);

OAI311xp33_ASAP7_75t_L g18224 ( 
.A1(n_18148),
.A2(n_4080),
.A3(n_4077),
.B1(n_4079),
.C1(n_4083),
.Y(n_18224)
);

OAI211xp5_ASAP7_75t_SL g18225 ( 
.A1(n_18170),
.A2(n_4084),
.B(n_4080),
.C(n_4083),
.Y(n_18225)
);

NAND3xp33_ASAP7_75t_SL g18226 ( 
.A(n_18153),
.B(n_4084),
.C(n_4085),
.Y(n_18226)
);

NOR2xp33_ASAP7_75t_L g18227 ( 
.A(n_18175),
.B(n_4085),
.Y(n_18227)
);

INVx2_ASAP7_75t_L g18228 ( 
.A(n_18184),
.Y(n_18228)
);

NOR3xp33_ASAP7_75t_L g18229 ( 
.A(n_18181),
.B(n_18191),
.C(n_18144),
.Y(n_18229)
);

INVx1_ASAP7_75t_L g18230 ( 
.A(n_18211),
.Y(n_18230)
);

NAND4xp25_ASAP7_75t_L g18231 ( 
.A(n_18201),
.B(n_4088),
.C(n_4086),
.D(n_4087),
.Y(n_18231)
);

AOI22xp5_ASAP7_75t_L g18232 ( 
.A1(n_18165),
.A2(n_4088),
.B1(n_4086),
.B2(n_4087),
.Y(n_18232)
);

NOR3xp33_ASAP7_75t_SL g18233 ( 
.A(n_18161),
.B(n_4089),
.C(n_4090),
.Y(n_18233)
);

AND2x4_ASAP7_75t_L g18234 ( 
.A(n_18146),
.B(n_4573),
.Y(n_18234)
);

AOI221xp5_ASAP7_75t_L g18235 ( 
.A1(n_18197),
.A2(n_18147),
.B1(n_18185),
.B2(n_18156),
.C(n_18143),
.Y(n_18235)
);

INVx1_ASAP7_75t_L g18236 ( 
.A(n_18186),
.Y(n_18236)
);

OAI322xp33_ASAP7_75t_L g18237 ( 
.A1(n_18158),
.A2(n_4094),
.A3(n_4093),
.B1(n_4091),
.B2(n_4089),
.C1(n_4090),
.C2(n_4092),
.Y(n_18237)
);

NOR3xp33_ASAP7_75t_L g18238 ( 
.A(n_18204),
.B(n_18180),
.C(n_18189),
.Y(n_18238)
);

NAND4xp25_ASAP7_75t_L g18239 ( 
.A(n_18190),
.B(n_4093),
.C(n_4091),
.D(n_4092),
.Y(n_18239)
);

AOI21xp5_ASAP7_75t_L g18240 ( 
.A1(n_18162),
.A2(n_4094),
.B(n_4096),
.Y(n_18240)
);

NAND5xp2_ASAP7_75t_L g18241 ( 
.A(n_18172),
.B(n_4098),
.C(n_4100),
.D(n_4097),
.E(n_4099),
.Y(n_18241)
);

NOR2x1p5_ASAP7_75t_L g18242 ( 
.A(n_18164),
.B(n_4096),
.Y(n_18242)
);

AOI22xp5_ASAP7_75t_L g18243 ( 
.A1(n_18196),
.A2(n_4100),
.B1(n_4097),
.B2(n_4099),
.Y(n_18243)
);

NAND2xp5_ASAP7_75t_L g18244 ( 
.A(n_18202),
.B(n_4101),
.Y(n_18244)
);

AOI22xp5_ASAP7_75t_L g18245 ( 
.A1(n_18151),
.A2(n_18155),
.B1(n_18173),
.B2(n_18145),
.Y(n_18245)
);

AOI22xp5_ASAP7_75t_L g18246 ( 
.A1(n_18212),
.A2(n_18163),
.B1(n_18149),
.B2(n_18194),
.Y(n_18246)
);

AND4x1_ASAP7_75t_L g18247 ( 
.A(n_18141),
.B(n_4103),
.C(n_4104),
.D(n_4102),
.Y(n_18247)
);

NAND4xp25_ASAP7_75t_SL g18248 ( 
.A(n_18179),
.B(n_18176),
.C(n_18206),
.D(n_18210),
.Y(n_18248)
);

INVx1_ASAP7_75t_L g18249 ( 
.A(n_18195),
.Y(n_18249)
);

XOR2xp5_ASAP7_75t_L g18250 ( 
.A(n_18168),
.B(n_4101),
.Y(n_18250)
);

NAND4xp25_ASAP7_75t_L g18251 ( 
.A(n_18174),
.B(n_4106),
.C(n_4103),
.D(n_4105),
.Y(n_18251)
);

INVx1_ASAP7_75t_L g18252 ( 
.A(n_18208),
.Y(n_18252)
);

NAND2xp5_ASAP7_75t_L g18253 ( 
.A(n_18205),
.B(n_4106),
.Y(n_18253)
);

INVx1_ASAP7_75t_L g18254 ( 
.A(n_18217),
.Y(n_18254)
);

NAND2xp5_ASAP7_75t_SL g18255 ( 
.A(n_18183),
.B(n_4107),
.Y(n_18255)
);

AOI211xp5_ASAP7_75t_L g18256 ( 
.A1(n_18150),
.A2(n_18154),
.B(n_18157),
.C(n_18152),
.Y(n_18256)
);

NOR4xp25_ASAP7_75t_L g18257 ( 
.A(n_18142),
.B(n_4109),
.C(n_4107),
.D(n_4108),
.Y(n_18257)
);

XOR2xp5_ASAP7_75t_L g18258 ( 
.A(n_18171),
.B(n_4108),
.Y(n_18258)
);

AOI22xp5_ASAP7_75t_L g18259 ( 
.A1(n_18140),
.A2(n_4111),
.B1(n_4109),
.B2(n_4110),
.Y(n_18259)
);

OAI221xp5_ASAP7_75t_L g18260 ( 
.A1(n_18167),
.A2(n_4112),
.B1(n_4110),
.B2(n_4111),
.C(n_4113),
.Y(n_18260)
);

AOI21xp33_ASAP7_75t_SL g18261 ( 
.A1(n_18207),
.A2(n_4112),
.B(n_4113),
.Y(n_18261)
);

NAND2xp5_ASAP7_75t_L g18262 ( 
.A(n_18215),
.B(n_4114),
.Y(n_18262)
);

OAI211xp5_ASAP7_75t_L g18263 ( 
.A1(n_18214),
.A2(n_4117),
.B(n_4115),
.C(n_4116),
.Y(n_18263)
);

NAND2xp33_ASAP7_75t_L g18264 ( 
.A(n_18216),
.B(n_4115),
.Y(n_18264)
);

OA22x2_ASAP7_75t_L g18265 ( 
.A1(n_18192),
.A2(n_4118),
.B1(n_4116),
.B2(n_4117),
.Y(n_18265)
);

INVx1_ASAP7_75t_L g18266 ( 
.A(n_18187),
.Y(n_18266)
);

OR2x2_ASAP7_75t_L g18267 ( 
.A(n_18169),
.B(n_4118),
.Y(n_18267)
);

NAND2xp5_ASAP7_75t_L g18268 ( 
.A(n_18177),
.B(n_4119),
.Y(n_18268)
);

OAI222xp33_ASAP7_75t_L g18269 ( 
.A1(n_18209),
.A2(n_4122),
.B1(n_4125),
.B2(n_4120),
.C1(n_4121),
.C2(n_4124),
.Y(n_18269)
);

OAI22xp5_ASAP7_75t_L g18270 ( 
.A1(n_18198),
.A2(n_4124),
.B1(n_4121),
.B2(n_4122),
.Y(n_18270)
);

AOI22xp5_ASAP7_75t_L g18271 ( 
.A1(n_18182),
.A2(n_4128),
.B1(n_4126),
.B2(n_4127),
.Y(n_18271)
);

NOR2xp33_ASAP7_75t_L g18272 ( 
.A(n_18199),
.B(n_4126),
.Y(n_18272)
);

BUFx2_ASAP7_75t_L g18273 ( 
.A(n_18203),
.Y(n_18273)
);

AOI22xp33_ASAP7_75t_L g18274 ( 
.A1(n_18193),
.A2(n_4130),
.B1(n_4128),
.B2(n_4129),
.Y(n_18274)
);

NOR3xp33_ASAP7_75t_L g18275 ( 
.A(n_18213),
.B(n_4129),
.C(n_4130),
.Y(n_18275)
);

OAI211xp5_ASAP7_75t_SL g18276 ( 
.A1(n_18160),
.A2(n_4133),
.B(n_4131),
.C(n_4132),
.Y(n_18276)
);

NAND3xp33_ASAP7_75t_SL g18277 ( 
.A(n_18153),
.B(n_4131),
.C(n_4132),
.Y(n_18277)
);

OAI22xp5_ASAP7_75t_L g18278 ( 
.A1(n_18188),
.A2(n_4135),
.B1(n_4133),
.B2(n_4134),
.Y(n_18278)
);

XOR2x2_ASAP7_75t_L g18279 ( 
.A(n_18186),
.B(n_4134),
.Y(n_18279)
);

NOR3xp33_ASAP7_75t_L g18280 ( 
.A(n_18166),
.B(n_4136),
.C(n_4137),
.Y(n_18280)
);

INVx1_ASAP7_75t_L g18281 ( 
.A(n_18211),
.Y(n_18281)
);

AND4x1_ASAP7_75t_L g18282 ( 
.A(n_18144),
.B(n_4139),
.C(n_4140),
.D(n_4138),
.Y(n_18282)
);

NAND4xp25_ASAP7_75t_L g18283 ( 
.A(n_18188),
.B(n_4140),
.C(n_4137),
.D(n_4138),
.Y(n_18283)
);

AOI22xp5_ASAP7_75t_L g18284 ( 
.A1(n_18188),
.A2(n_4143),
.B1(n_4141),
.B2(n_4142),
.Y(n_18284)
);

OAI21xp33_ASAP7_75t_L g18285 ( 
.A1(n_18188),
.A2(n_4142),
.B(n_4144),
.Y(n_18285)
);

AND2x4_ASAP7_75t_L g18286 ( 
.A(n_18211),
.B(n_4560),
.Y(n_18286)
);

NAND4xp25_ASAP7_75t_L g18287 ( 
.A(n_18188),
.B(n_4147),
.C(n_4145),
.D(n_4146),
.Y(n_18287)
);

AOI221xp5_ASAP7_75t_L g18288 ( 
.A1(n_18188),
.A2(n_4147),
.B1(n_4145),
.B2(n_4146),
.C(n_4148),
.Y(n_18288)
);

OAI221xp5_ASAP7_75t_L g18289 ( 
.A1(n_18206),
.A2(n_4150),
.B1(n_4148),
.B2(n_4149),
.C(n_4151),
.Y(n_18289)
);

NAND5xp2_ASAP7_75t_L g18290 ( 
.A(n_18188),
.B(n_4151),
.C(n_4153),
.D(n_4150),
.E(n_4152),
.Y(n_18290)
);

AOI22xp33_ASAP7_75t_L g18291 ( 
.A1(n_18178),
.A2(n_4154),
.B1(n_4149),
.B2(n_4153),
.Y(n_18291)
);

AOI211x1_ASAP7_75t_L g18292 ( 
.A1(n_18166),
.A2(n_4156),
.B(n_4154),
.C(n_4155),
.Y(n_18292)
);

NAND4xp25_ASAP7_75t_L g18293 ( 
.A(n_18188),
.B(n_4157),
.C(n_4155),
.D(n_4156),
.Y(n_18293)
);

INVx2_ASAP7_75t_L g18294 ( 
.A(n_18184),
.Y(n_18294)
);

INVx1_ASAP7_75t_L g18295 ( 
.A(n_18211),
.Y(n_18295)
);

NAND4xp25_ASAP7_75t_SL g18296 ( 
.A(n_18179),
.B(n_4160),
.C(n_4158),
.D(n_4159),
.Y(n_18296)
);

AOI21xp5_ASAP7_75t_L g18297 ( 
.A1(n_18148),
.A2(n_4160),
.B(n_4161),
.Y(n_18297)
);

OAI211xp5_ASAP7_75t_L g18298 ( 
.A1(n_18188),
.A2(n_4163),
.B(n_4161),
.C(n_4162),
.Y(n_18298)
);

NAND3xp33_ASAP7_75t_SL g18299 ( 
.A(n_18153),
.B(n_4162),
.C(n_4163),
.Y(n_18299)
);

INVx3_ASAP7_75t_L g18300 ( 
.A(n_18178),
.Y(n_18300)
);

INVx2_ASAP7_75t_SL g18301 ( 
.A(n_18202),
.Y(n_18301)
);

INVx1_ASAP7_75t_L g18302 ( 
.A(n_18211),
.Y(n_18302)
);

NOR3xp33_ASAP7_75t_SL g18303 ( 
.A(n_18159),
.B(n_4164),
.C(n_4166),
.Y(n_18303)
);

NOR2xp33_ASAP7_75t_L g18304 ( 
.A(n_18188),
.B(n_4164),
.Y(n_18304)
);

OR4x1_ASAP7_75t_L g18305 ( 
.A(n_18170),
.B(n_4168),
.C(n_4166),
.D(n_4167),
.Y(n_18305)
);

OA211x2_ASAP7_75t_L g18306 ( 
.A1(n_18188),
.A2(n_4169),
.B(n_4167),
.C(n_4168),
.Y(n_18306)
);

NAND3xp33_ASAP7_75t_SL g18307 ( 
.A(n_18153),
.B(n_4169),
.C(n_4170),
.Y(n_18307)
);

NAND4xp25_ASAP7_75t_L g18308 ( 
.A(n_18188),
.B(n_4172),
.C(n_4170),
.D(n_4171),
.Y(n_18308)
);

NOR4xp25_ASAP7_75t_L g18309 ( 
.A(n_18160),
.B(n_4175),
.C(n_4173),
.D(n_4174),
.Y(n_18309)
);

OAI22xp5_ASAP7_75t_L g18310 ( 
.A1(n_18188),
.A2(n_4176),
.B1(n_4173),
.B2(n_4175),
.Y(n_18310)
);

NOR2x1p5_ASAP7_75t_L g18311 ( 
.A(n_18300),
.B(n_4176),
.Y(n_18311)
);

AOI21xp5_ASAP7_75t_L g18312 ( 
.A1(n_18229),
.A2(n_4177),
.B(n_4178),
.Y(n_18312)
);

INVx5_ASAP7_75t_L g18313 ( 
.A(n_18300),
.Y(n_18313)
);

AOI22xp5_ASAP7_75t_L g18314 ( 
.A1(n_18304),
.A2(n_4180),
.B1(n_4178),
.B2(n_4179),
.Y(n_18314)
);

INVx1_ASAP7_75t_L g18315 ( 
.A(n_18242),
.Y(n_18315)
);

NAND2xp5_ASAP7_75t_L g18316 ( 
.A(n_18227),
.B(n_4562),
.Y(n_18316)
);

NAND3xp33_ASAP7_75t_L g18317 ( 
.A(n_18238),
.B(n_4179),
.C(n_4181),
.Y(n_18317)
);

INVx1_ASAP7_75t_L g18318 ( 
.A(n_18253),
.Y(n_18318)
);

AOI22xp5_ASAP7_75t_L g18319 ( 
.A1(n_18296),
.A2(n_18226),
.B1(n_18299),
.B2(n_18277),
.Y(n_18319)
);

NAND2xp5_ASAP7_75t_L g18320 ( 
.A(n_18233),
.B(n_4563),
.Y(n_18320)
);

INVx2_ASAP7_75t_L g18321 ( 
.A(n_18305),
.Y(n_18321)
);

AOI22xp5_ASAP7_75t_L g18322 ( 
.A1(n_18307),
.A2(n_4183),
.B1(n_4181),
.B2(n_4182),
.Y(n_18322)
);

INVxp67_ASAP7_75t_SL g18323 ( 
.A(n_18244),
.Y(n_18323)
);

INVx1_ASAP7_75t_L g18324 ( 
.A(n_18279),
.Y(n_18324)
);

NAND2xp5_ASAP7_75t_L g18325 ( 
.A(n_18219),
.B(n_4564),
.Y(n_18325)
);

AOI22xp5_ASAP7_75t_L g18326 ( 
.A1(n_18275),
.A2(n_4184),
.B1(n_4182),
.B2(n_4183),
.Y(n_18326)
);

AND2x2_ASAP7_75t_L g18327 ( 
.A(n_18228),
.B(n_4185),
.Y(n_18327)
);

INVx1_ASAP7_75t_L g18328 ( 
.A(n_18303),
.Y(n_18328)
);

AOI22xp5_ASAP7_75t_L g18329 ( 
.A1(n_18280),
.A2(n_4188),
.B1(n_4185),
.B2(n_4187),
.Y(n_18329)
);

AOI22xp5_ASAP7_75t_L g18330 ( 
.A1(n_18276),
.A2(n_4189),
.B1(n_4187),
.B2(n_4188),
.Y(n_18330)
);

NOR2xp33_ASAP7_75t_L g18331 ( 
.A(n_18248),
.B(n_18294),
.Y(n_18331)
);

INVx1_ASAP7_75t_L g18332 ( 
.A(n_18268),
.Y(n_18332)
);

INVx2_ASAP7_75t_L g18333 ( 
.A(n_18286),
.Y(n_18333)
);

OAI22xp5_ASAP7_75t_L g18334 ( 
.A1(n_18271),
.A2(n_4191),
.B1(n_4192),
.B2(n_4190),
.Y(n_18334)
);

NAND2xp5_ASAP7_75t_L g18335 ( 
.A(n_18286),
.B(n_4576),
.Y(n_18335)
);

AOI22xp5_ASAP7_75t_L g18336 ( 
.A1(n_18265),
.A2(n_4192),
.B1(n_4189),
.B2(n_4190),
.Y(n_18336)
);

AOI22xp5_ASAP7_75t_L g18337 ( 
.A1(n_18255),
.A2(n_4195),
.B1(n_4193),
.B2(n_4194),
.Y(n_18337)
);

HB1xp67_ASAP7_75t_L g18338 ( 
.A(n_18262),
.Y(n_18338)
);

INVx1_ASAP7_75t_L g18339 ( 
.A(n_18306),
.Y(n_18339)
);

INVx2_ASAP7_75t_L g18340 ( 
.A(n_18234),
.Y(n_18340)
);

INVx2_ASAP7_75t_L g18341 ( 
.A(n_18234),
.Y(n_18341)
);

NOR2x1_ASAP7_75t_L g18342 ( 
.A(n_18230),
.B(n_4194),
.Y(n_18342)
);

NOR2xp67_ASAP7_75t_L g18343 ( 
.A(n_18301),
.B(n_4559),
.Y(n_18343)
);

NAND2xp5_ASAP7_75t_L g18344 ( 
.A(n_18240),
.B(n_4560),
.Y(n_18344)
);

AND3x4_ASAP7_75t_L g18345 ( 
.A(n_18223),
.B(n_4193),
.C(n_4195),
.Y(n_18345)
);

NOR3xp33_ASAP7_75t_L g18346 ( 
.A(n_18235),
.B(n_4196),
.C(n_4197),
.Y(n_18346)
);

NAND2xp5_ASAP7_75t_L g18347 ( 
.A(n_18272),
.B(n_18292),
.Y(n_18347)
);

AOI222xp33_ASAP7_75t_L g18348 ( 
.A1(n_18273),
.A2(n_4198),
.B1(n_4200),
.B2(n_4196),
.C1(n_4197),
.C2(n_4199),
.Y(n_18348)
);

OAI22x1_ASAP7_75t_L g18349 ( 
.A1(n_18245),
.A2(n_4200),
.B1(n_4198),
.B2(n_4199),
.Y(n_18349)
);

INVx2_ASAP7_75t_L g18350 ( 
.A(n_18250),
.Y(n_18350)
);

CKINVDCx20_ASAP7_75t_R g18351 ( 
.A(n_18266),
.Y(n_18351)
);

NAND5xp2_ASAP7_75t_L g18352 ( 
.A(n_18256),
.B(n_4203),
.C(n_4201),
.D(n_4202),
.E(n_4204),
.Y(n_18352)
);

AOI21xp5_ASAP7_75t_L g18353 ( 
.A1(n_18281),
.A2(n_4201),
.B(n_4202),
.Y(n_18353)
);

AOI21xp5_ASAP7_75t_L g18354 ( 
.A1(n_18295),
.A2(n_4203),
.B(n_4204),
.Y(n_18354)
);

INVxp67_ASAP7_75t_L g18355 ( 
.A(n_18302),
.Y(n_18355)
);

INVx2_ASAP7_75t_SL g18356 ( 
.A(n_18282),
.Y(n_18356)
);

OAI22xp5_ASAP7_75t_L g18357 ( 
.A1(n_18289),
.A2(n_4207),
.B1(n_4208),
.B2(n_4206),
.Y(n_18357)
);

INVxp33_ASAP7_75t_L g18358 ( 
.A(n_18283),
.Y(n_18358)
);

A2O1A1Ixp33_ASAP7_75t_L g18359 ( 
.A1(n_18285),
.A2(n_18297),
.B(n_18264),
.C(n_18246),
.Y(n_18359)
);

NAND2xp5_ASAP7_75t_L g18360 ( 
.A(n_18309),
.B(n_4583),
.Y(n_18360)
);

NAND2xp5_ASAP7_75t_L g18361 ( 
.A(n_18298),
.B(n_18257),
.Y(n_18361)
);

BUFx2_ASAP7_75t_L g18362 ( 
.A(n_18287),
.Y(n_18362)
);

INVx2_ASAP7_75t_L g18363 ( 
.A(n_18258),
.Y(n_18363)
);

OAI22xp5_ASAP7_75t_L g18364 ( 
.A1(n_18221),
.A2(n_4208),
.B1(n_4209),
.B2(n_4206),
.Y(n_18364)
);

INVx2_ASAP7_75t_L g18365 ( 
.A(n_18267),
.Y(n_18365)
);

OAI22xp5_ASAP7_75t_SL g18366 ( 
.A1(n_18236),
.A2(n_4216),
.B1(n_4224),
.B2(n_4205),
.Y(n_18366)
);

NAND5xp2_ASAP7_75t_L g18367 ( 
.A(n_18249),
.B(n_4210),
.C(n_4205),
.D(n_4209),
.E(n_4211),
.Y(n_18367)
);

INVx2_ASAP7_75t_L g18368 ( 
.A(n_18284),
.Y(n_18368)
);

INVx1_ASAP7_75t_L g18369 ( 
.A(n_18278),
.Y(n_18369)
);

INVx2_ASAP7_75t_L g18370 ( 
.A(n_18232),
.Y(n_18370)
);

INVx2_ASAP7_75t_L g18371 ( 
.A(n_18260),
.Y(n_18371)
);

AOI22xp5_ASAP7_75t_L g18372 ( 
.A1(n_18225),
.A2(n_4212),
.B1(n_4210),
.B2(n_4211),
.Y(n_18372)
);

NAND2xp5_ASAP7_75t_L g18373 ( 
.A(n_18261),
.B(n_4563),
.Y(n_18373)
);

INVxp67_ASAP7_75t_SL g18374 ( 
.A(n_18252),
.Y(n_18374)
);

AOI32xp33_ASAP7_75t_L g18375 ( 
.A1(n_18254),
.A2(n_4214),
.A3(n_4212),
.B1(n_4213),
.B2(n_4215),
.Y(n_18375)
);

INVx2_ASAP7_75t_L g18376 ( 
.A(n_18270),
.Y(n_18376)
);

INVx1_ASAP7_75t_L g18377 ( 
.A(n_18310),
.Y(n_18377)
);

AOI22x1_ASAP7_75t_L g18378 ( 
.A1(n_18224),
.A2(n_4217),
.B1(n_4215),
.B2(n_4216),
.Y(n_18378)
);

INVx2_ASAP7_75t_L g18379 ( 
.A(n_18243),
.Y(n_18379)
);

AOI222xp33_ASAP7_75t_L g18380 ( 
.A1(n_18269),
.A2(n_4220),
.B1(n_4222),
.B2(n_4218),
.C1(n_4219),
.C2(n_4221),
.Y(n_18380)
);

NAND2xp5_ASAP7_75t_L g18381 ( 
.A(n_18288),
.B(n_4577),
.Y(n_18381)
);

NAND2x1_ASAP7_75t_SL g18382 ( 
.A(n_18259),
.B(n_4218),
.Y(n_18382)
);

OR3x1_ASAP7_75t_L g18383 ( 
.A(n_18241),
.B(n_4219),
.C(n_4221),
.Y(n_18383)
);

NAND4xp25_ASAP7_75t_SL g18384 ( 
.A(n_18274),
.B(n_4230),
.C(n_4239),
.D(n_4222),
.Y(n_18384)
);

INVx1_ASAP7_75t_L g18385 ( 
.A(n_18293),
.Y(n_18385)
);

OAI21xp33_ASAP7_75t_L g18386 ( 
.A1(n_18290),
.A2(n_4223),
.B(n_4224),
.Y(n_18386)
);

OAI22xp5_ASAP7_75t_L g18387 ( 
.A1(n_18263),
.A2(n_4226),
.B1(n_4227),
.B2(n_4225),
.Y(n_18387)
);

INVx1_ASAP7_75t_L g18388 ( 
.A(n_18308),
.Y(n_18388)
);

AOI211xp5_ASAP7_75t_L g18389 ( 
.A1(n_18222),
.A2(n_18237),
.B(n_18239),
.C(n_18251),
.Y(n_18389)
);

AOI22xp33_ASAP7_75t_L g18390 ( 
.A1(n_18231),
.A2(n_4226),
.B1(n_4223),
.B2(n_4225),
.Y(n_18390)
);

NAND4xp75_ASAP7_75t_L g18391 ( 
.A(n_18218),
.B(n_4229),
.C(n_4227),
.D(n_4228),
.Y(n_18391)
);

INVx1_ASAP7_75t_L g18392 ( 
.A(n_18247),
.Y(n_18392)
);

AOI211xp5_ASAP7_75t_L g18393 ( 
.A1(n_18220),
.A2(n_4232),
.B(n_4228),
.C(n_4231),
.Y(n_18393)
);

INVx1_ASAP7_75t_L g18394 ( 
.A(n_18320),
.Y(n_18394)
);

XNOR2x1_ASAP7_75t_L g18395 ( 
.A(n_18345),
.B(n_18291),
.Y(n_18395)
);

INVx2_ASAP7_75t_L g18396 ( 
.A(n_18311),
.Y(n_18396)
);

NAND4xp75_ASAP7_75t_L g18397 ( 
.A(n_18331),
.B(n_4233),
.C(n_4231),
.D(n_4232),
.Y(n_18397)
);

INVx2_ASAP7_75t_L g18398 ( 
.A(n_18349),
.Y(n_18398)
);

AOI22xp5_ASAP7_75t_L g18399 ( 
.A1(n_18386),
.A2(n_4235),
.B1(n_4233),
.B2(n_4234),
.Y(n_18399)
);

INVx3_ASAP7_75t_L g18400 ( 
.A(n_18313),
.Y(n_18400)
);

INVx2_ASAP7_75t_L g18401 ( 
.A(n_18342),
.Y(n_18401)
);

NAND2xp5_ASAP7_75t_L g18402 ( 
.A(n_18372),
.B(n_4236),
.Y(n_18402)
);

INVx1_ASAP7_75t_L g18403 ( 
.A(n_18325),
.Y(n_18403)
);

BUFx2_ASAP7_75t_L g18404 ( 
.A(n_18382),
.Y(n_18404)
);

NAND2xp5_ASAP7_75t_L g18405 ( 
.A(n_18330),
.B(n_18336),
.Y(n_18405)
);

NAND2xp5_ASAP7_75t_L g18406 ( 
.A(n_18313),
.B(n_4236),
.Y(n_18406)
);

AOI21xp5_ASAP7_75t_L g18407 ( 
.A1(n_18374),
.A2(n_18355),
.B(n_18339),
.Y(n_18407)
);

INVx2_ASAP7_75t_L g18408 ( 
.A(n_18378),
.Y(n_18408)
);

XNOR2xp5_ASAP7_75t_L g18409 ( 
.A(n_18383),
.B(n_4238),
.Y(n_18409)
);

AOI22xp5_ASAP7_75t_L g18410 ( 
.A1(n_18384),
.A2(n_4240),
.B1(n_4238),
.B2(n_4239),
.Y(n_18410)
);

INVx1_ASAP7_75t_L g18411 ( 
.A(n_18360),
.Y(n_18411)
);

INVx1_ASAP7_75t_L g18412 ( 
.A(n_18373),
.Y(n_18412)
);

INVx2_ASAP7_75t_L g18413 ( 
.A(n_18391),
.Y(n_18413)
);

INVx2_ASAP7_75t_L g18414 ( 
.A(n_18316),
.Y(n_18414)
);

INVx1_ASAP7_75t_L g18415 ( 
.A(n_18344),
.Y(n_18415)
);

INVx2_ASAP7_75t_L g18416 ( 
.A(n_18335),
.Y(n_18416)
);

INVx1_ASAP7_75t_L g18417 ( 
.A(n_18343),
.Y(n_18417)
);

AOI22xp5_ASAP7_75t_L g18418 ( 
.A1(n_18351),
.A2(n_4242),
.B1(n_4240),
.B2(n_4241),
.Y(n_18418)
);

INVx3_ASAP7_75t_L g18419 ( 
.A(n_18313),
.Y(n_18419)
);

INVx2_ASAP7_75t_L g18420 ( 
.A(n_18317),
.Y(n_18420)
);

O2A1O1Ixp33_ASAP7_75t_SL g18421 ( 
.A1(n_18359),
.A2(n_4244),
.B(n_4241),
.C(n_4243),
.Y(n_18421)
);

INVx2_ASAP7_75t_L g18422 ( 
.A(n_18333),
.Y(n_18422)
);

OA22x2_ASAP7_75t_L g18423 ( 
.A1(n_18322),
.A2(n_4245),
.B1(n_4243),
.B2(n_4244),
.Y(n_18423)
);

INVx5_ASAP7_75t_L g18424 ( 
.A(n_18356),
.Y(n_18424)
);

OAI22xp5_ASAP7_75t_SL g18425 ( 
.A1(n_18321),
.A2(n_4247),
.B1(n_4245),
.B2(n_4246),
.Y(n_18425)
);

NAND2xp5_ASAP7_75t_L g18426 ( 
.A(n_18390),
.B(n_18357),
.Y(n_18426)
);

OAI22x1_ASAP7_75t_L g18427 ( 
.A1(n_18340),
.A2(n_4248),
.B1(n_4249),
.B2(n_4247),
.Y(n_18427)
);

INVx1_ASAP7_75t_L g18428 ( 
.A(n_18381),
.Y(n_18428)
);

OR2x2_ASAP7_75t_L g18429 ( 
.A(n_18352),
.B(n_4246),
.Y(n_18429)
);

CKINVDCx20_ASAP7_75t_R g18430 ( 
.A(n_18362),
.Y(n_18430)
);

INVx1_ASAP7_75t_L g18431 ( 
.A(n_18361),
.Y(n_18431)
);

INVx1_ASAP7_75t_L g18432 ( 
.A(n_18392),
.Y(n_18432)
);

XNOR2x1_ASAP7_75t_L g18433 ( 
.A(n_18350),
.B(n_4248),
.Y(n_18433)
);

INVx3_ASAP7_75t_L g18434 ( 
.A(n_18341),
.Y(n_18434)
);

AOI22xp5_ASAP7_75t_L g18435 ( 
.A1(n_18334),
.A2(n_4251),
.B1(n_4249),
.B2(n_4250),
.Y(n_18435)
);

INVx2_ASAP7_75t_L g18436 ( 
.A(n_18337),
.Y(n_18436)
);

INVx1_ASAP7_75t_L g18437 ( 
.A(n_18347),
.Y(n_18437)
);

XNOR2x1_ASAP7_75t_L g18438 ( 
.A(n_18363),
.B(n_4250),
.Y(n_18438)
);

AND2x4_ASAP7_75t_L g18439 ( 
.A(n_18328),
.B(n_4251),
.Y(n_18439)
);

OAI22xp5_ASAP7_75t_L g18440 ( 
.A1(n_18329),
.A2(n_4254),
.B1(n_4252),
.B2(n_4253),
.Y(n_18440)
);

NAND2xp5_ASAP7_75t_L g18441 ( 
.A(n_18393),
.B(n_18380),
.Y(n_18441)
);

INVx5_ASAP7_75t_L g18442 ( 
.A(n_18365),
.Y(n_18442)
);

NAND3x1_ASAP7_75t_L g18443 ( 
.A(n_18315),
.B(n_4252),
.C(n_4254),
.Y(n_18443)
);

INVx2_ASAP7_75t_L g18444 ( 
.A(n_18314),
.Y(n_18444)
);

XOR2xp5_ASAP7_75t_L g18445 ( 
.A(n_18358),
.B(n_4257),
.Y(n_18445)
);

NAND2xp5_ASAP7_75t_SL g18446 ( 
.A(n_18346),
.B(n_4256),
.Y(n_18446)
);

OAI222xp33_ASAP7_75t_L g18447 ( 
.A1(n_18409),
.A2(n_18319),
.B1(n_18388),
.B2(n_18385),
.C1(n_18377),
.C2(n_18369),
.Y(n_18447)
);

NOR3xp33_ASAP7_75t_SL g18448 ( 
.A(n_18407),
.B(n_18324),
.C(n_18332),
.Y(n_18448)
);

NAND5xp2_ASAP7_75t_L g18449 ( 
.A(n_18432),
.B(n_18389),
.C(n_18318),
.D(n_18323),
.E(n_18326),
.Y(n_18449)
);

HB1xp67_ASAP7_75t_L g18450 ( 
.A(n_18400),
.Y(n_18450)
);

AO21x1_ASAP7_75t_L g18451 ( 
.A1(n_18417),
.A2(n_18376),
.B(n_18370),
.Y(n_18451)
);

OAI22xp5_ASAP7_75t_SL g18452 ( 
.A1(n_18413),
.A2(n_18371),
.B1(n_18379),
.B2(n_18368),
.Y(n_18452)
);

AOI22xp33_ASAP7_75t_L g18453 ( 
.A1(n_18419),
.A2(n_18338),
.B1(n_18387),
.B2(n_18364),
.Y(n_18453)
);

INVx1_ASAP7_75t_L g18454 ( 
.A(n_18402),
.Y(n_18454)
);

INVx1_ASAP7_75t_L g18455 ( 
.A(n_18446),
.Y(n_18455)
);

OAI22xp5_ASAP7_75t_L g18456 ( 
.A1(n_18399),
.A2(n_18410),
.B1(n_18435),
.B2(n_18429),
.Y(n_18456)
);

INVx1_ASAP7_75t_L g18457 ( 
.A(n_18395),
.Y(n_18457)
);

INVxp67_ASAP7_75t_L g18458 ( 
.A(n_18422),
.Y(n_18458)
);

CKINVDCx20_ASAP7_75t_R g18459 ( 
.A(n_18430),
.Y(n_18459)
);

INVxp67_ASAP7_75t_SL g18460 ( 
.A(n_18408),
.Y(n_18460)
);

INVx1_ASAP7_75t_L g18461 ( 
.A(n_18396),
.Y(n_18461)
);

OAI221xp5_ASAP7_75t_L g18462 ( 
.A1(n_18434),
.A2(n_18312),
.B1(n_18354),
.B2(n_18353),
.C(n_18375),
.Y(n_18462)
);

OAI22xp5_ASAP7_75t_L g18463 ( 
.A1(n_18424),
.A2(n_18366),
.B1(n_18367),
.B2(n_18327),
.Y(n_18463)
);

AOI21xp5_ASAP7_75t_L g18464 ( 
.A1(n_18426),
.A2(n_18348),
.B(n_4260),
.Y(n_18464)
);

AO21x2_ASAP7_75t_L g18465 ( 
.A1(n_18411),
.A2(n_4257),
.B(n_4259),
.Y(n_18465)
);

INVx1_ASAP7_75t_L g18466 ( 
.A(n_18405),
.Y(n_18466)
);

HB1xp67_ASAP7_75t_L g18467 ( 
.A(n_18424),
.Y(n_18467)
);

INVx2_ASAP7_75t_L g18468 ( 
.A(n_18438),
.Y(n_18468)
);

AOI21xp5_ASAP7_75t_L g18469 ( 
.A1(n_18441),
.A2(n_4262),
.B(n_4261),
.Y(n_18469)
);

INVx2_ASAP7_75t_L g18470 ( 
.A(n_18433),
.Y(n_18470)
);

INVx2_ASAP7_75t_L g18471 ( 
.A(n_18397),
.Y(n_18471)
);

OAI22xp5_ASAP7_75t_L g18472 ( 
.A1(n_18442),
.A2(n_4263),
.B1(n_4259),
.B2(n_4261),
.Y(n_18472)
);

AO22x2_ASAP7_75t_L g18473 ( 
.A1(n_18401),
.A2(n_4265),
.B1(n_4263),
.B2(n_4264),
.Y(n_18473)
);

INVx1_ASAP7_75t_L g18474 ( 
.A(n_18404),
.Y(n_18474)
);

INVx1_ASAP7_75t_SL g18475 ( 
.A(n_18442),
.Y(n_18475)
);

AOI22xp5_ASAP7_75t_L g18476 ( 
.A1(n_18440),
.A2(n_4274),
.B1(n_4282),
.B2(n_4265),
.Y(n_18476)
);

NOR2xp67_ASAP7_75t_L g18477 ( 
.A(n_18398),
.B(n_4267),
.Y(n_18477)
);

OR2x2_ASAP7_75t_L g18478 ( 
.A(n_18420),
.B(n_4269),
.Y(n_18478)
);

INVx1_ASAP7_75t_L g18479 ( 
.A(n_18423),
.Y(n_18479)
);

XOR2xp5_ASAP7_75t_L g18480 ( 
.A(n_18437),
.B(n_18431),
.Y(n_18480)
);

AOI22xp33_ASAP7_75t_L g18481 ( 
.A1(n_18416),
.A2(n_4575),
.B1(n_4582),
.B2(n_4571),
.Y(n_18481)
);

NAND3x1_ASAP7_75t_L g18482 ( 
.A(n_18412),
.B(n_4268),
.C(n_4269),
.Y(n_18482)
);

INVxp67_ASAP7_75t_SL g18483 ( 
.A(n_18444),
.Y(n_18483)
);

AND2x2_ASAP7_75t_L g18484 ( 
.A(n_18414),
.B(n_4271),
.Y(n_18484)
);

AND2x4_ASAP7_75t_L g18485 ( 
.A(n_18436),
.B(n_4271),
.Y(n_18485)
);

INVx1_ASAP7_75t_L g18486 ( 
.A(n_18415),
.Y(n_18486)
);

INVx1_ASAP7_75t_L g18487 ( 
.A(n_18467),
.Y(n_18487)
);

INVx1_ASAP7_75t_L g18488 ( 
.A(n_18450),
.Y(n_18488)
);

AOI22xp5_ASAP7_75t_L g18489 ( 
.A1(n_18459),
.A2(n_18475),
.B1(n_18458),
.B2(n_18452),
.Y(n_18489)
);

OAI22xp33_ASAP7_75t_L g18490 ( 
.A1(n_18476),
.A2(n_18403),
.B1(n_18394),
.B2(n_18428),
.Y(n_18490)
);

AOI22xp33_ASAP7_75t_L g18491 ( 
.A1(n_18461),
.A2(n_18425),
.B1(n_18445),
.B2(n_18427),
.Y(n_18491)
);

INVx1_ASAP7_75t_L g18492 ( 
.A(n_18451),
.Y(n_18492)
);

NAND2xp5_ASAP7_75t_L g18493 ( 
.A(n_18464),
.B(n_18421),
.Y(n_18493)
);

NAND2xp5_ASAP7_75t_L g18494 ( 
.A(n_18483),
.B(n_18443),
.Y(n_18494)
);

OAI31xp33_ASAP7_75t_L g18495 ( 
.A1(n_18463),
.A2(n_18447),
.A3(n_18474),
.B(n_18480),
.Y(n_18495)
);

INVx1_ASAP7_75t_L g18496 ( 
.A(n_18479),
.Y(n_18496)
);

OAI22xp33_ASAP7_75t_L g18497 ( 
.A1(n_18466),
.A2(n_18418),
.B1(n_18406),
.B2(n_18439),
.Y(n_18497)
);

INVxp67_ASAP7_75t_L g18498 ( 
.A(n_18460),
.Y(n_18498)
);

HB1xp67_ASAP7_75t_L g18499 ( 
.A(n_18477),
.Y(n_18499)
);

INVx1_ASAP7_75t_SL g18500 ( 
.A(n_18471),
.Y(n_18500)
);

AOI22xp5_ASAP7_75t_L g18501 ( 
.A1(n_18457),
.A2(n_4273),
.B1(n_4274),
.B2(n_4272),
.Y(n_18501)
);

AOI22xp33_ASAP7_75t_L g18502 ( 
.A1(n_18486),
.A2(n_4273),
.B1(n_4270),
.B2(n_4272),
.Y(n_18502)
);

INVx1_ASAP7_75t_L g18503 ( 
.A(n_18456),
.Y(n_18503)
);

INVx1_ASAP7_75t_L g18504 ( 
.A(n_18462),
.Y(n_18504)
);

INVx1_ASAP7_75t_L g18505 ( 
.A(n_18468),
.Y(n_18505)
);

INVx1_ASAP7_75t_L g18506 ( 
.A(n_18470),
.Y(n_18506)
);

AOI22xp5_ASAP7_75t_L g18507 ( 
.A1(n_18455),
.A2(n_4277),
.B1(n_4278),
.B2(n_4276),
.Y(n_18507)
);

NAND2xp5_ASAP7_75t_L g18508 ( 
.A(n_18453),
.B(n_4276),
.Y(n_18508)
);

AOI22xp33_ASAP7_75t_L g18509 ( 
.A1(n_18454),
.A2(n_4279),
.B1(n_4275),
.B2(n_4277),
.Y(n_18509)
);

INVx1_ASAP7_75t_L g18510 ( 
.A(n_18448),
.Y(n_18510)
);

AND2x2_ASAP7_75t_L g18511 ( 
.A(n_18469),
.B(n_4275),
.Y(n_18511)
);

INVx3_ASAP7_75t_L g18512 ( 
.A(n_18449),
.Y(n_18512)
);

AND2x2_ASAP7_75t_L g18513 ( 
.A(n_18465),
.B(n_4280),
.Y(n_18513)
);

AOI22xp5_ASAP7_75t_L g18514 ( 
.A1(n_18482),
.A2(n_4282),
.B1(n_4283),
.B2(n_4281),
.Y(n_18514)
);

AOI22xp5_ASAP7_75t_L g18515 ( 
.A1(n_18472),
.A2(n_4283),
.B1(n_4284),
.B2(n_4281),
.Y(n_18515)
);

AOI22xp5_ASAP7_75t_L g18516 ( 
.A1(n_18485),
.A2(n_4286),
.B1(n_4287),
.B2(n_4285),
.Y(n_18516)
);

OAI22x1_ASAP7_75t_L g18517 ( 
.A1(n_18478),
.A2(n_18484),
.B1(n_18481),
.B2(n_18473),
.Y(n_18517)
);

AOI22xp5_ASAP7_75t_L g18518 ( 
.A1(n_18473),
.A2(n_4287),
.B1(n_4288),
.B2(n_4286),
.Y(n_18518)
);

AOI22xp33_ASAP7_75t_SL g18519 ( 
.A1(n_18467),
.A2(n_4289),
.B1(n_4290),
.B2(n_4288),
.Y(n_18519)
);

AOI22xp5_ASAP7_75t_L g18520 ( 
.A1(n_18459),
.A2(n_4290),
.B1(n_4291),
.B2(n_4289),
.Y(n_18520)
);

OAI22xp5_ASAP7_75t_L g18521 ( 
.A1(n_18489),
.A2(n_4292),
.B1(n_4280),
.B2(n_4291),
.Y(n_18521)
);

AOI22xp33_ASAP7_75t_L g18522 ( 
.A1(n_18488),
.A2(n_4295),
.B1(n_4293),
.B2(n_4294),
.Y(n_18522)
);

NAND2x1p5_ASAP7_75t_L g18523 ( 
.A(n_18487),
.B(n_4293),
.Y(n_18523)
);

OAI22xp33_ASAP7_75t_L g18524 ( 
.A1(n_18492),
.A2(n_4296),
.B1(n_4294),
.B2(n_4295),
.Y(n_18524)
);

OA21x2_ASAP7_75t_L g18525 ( 
.A1(n_18494),
.A2(n_4304),
.B(n_4296),
.Y(n_18525)
);

INVx1_ASAP7_75t_L g18526 ( 
.A(n_18499),
.Y(n_18526)
);

NOR2xp33_ASAP7_75t_R g18527 ( 
.A(n_18512),
.B(n_4297),
.Y(n_18527)
);

NAND2xp5_ASAP7_75t_L g18528 ( 
.A(n_18513),
.B(n_4297),
.Y(n_18528)
);

A2O1A1Ixp33_ASAP7_75t_L g18529 ( 
.A1(n_18495),
.A2(n_4300),
.B(n_4298),
.C(n_4299),
.Y(n_18529)
);

OAI22x1_ASAP7_75t_L g18530 ( 
.A1(n_18498),
.A2(n_4300),
.B1(n_4298),
.B2(n_4299),
.Y(n_18530)
);

XOR2xp5_ASAP7_75t_L g18531 ( 
.A(n_18503),
.B(n_4301),
.Y(n_18531)
);

AND2x2_ASAP7_75t_SL g18532 ( 
.A(n_18496),
.B(n_18491),
.Y(n_18532)
);

NAND2xp5_ASAP7_75t_L g18533 ( 
.A(n_18512),
.B(n_4301),
.Y(n_18533)
);

OAI22xp5_ASAP7_75t_L g18534 ( 
.A1(n_18515),
.A2(n_4304),
.B1(n_4302),
.B2(n_4303),
.Y(n_18534)
);

NAND2xp5_ASAP7_75t_L g18535 ( 
.A(n_18505),
.B(n_4303),
.Y(n_18535)
);

INVx1_ASAP7_75t_L g18536 ( 
.A(n_18517),
.Y(n_18536)
);

OAI22xp5_ASAP7_75t_SL g18537 ( 
.A1(n_18500),
.A2(n_4307),
.B1(n_4305),
.B2(n_4306),
.Y(n_18537)
);

NAND3xp33_ASAP7_75t_SL g18538 ( 
.A(n_18510),
.B(n_4305),
.C(n_4306),
.Y(n_18538)
);

XNOR2x2_ASAP7_75t_L g18539 ( 
.A(n_18506),
.B(n_4307),
.Y(n_18539)
);

OAI21xp5_ASAP7_75t_L g18540 ( 
.A1(n_18504),
.A2(n_4309),
.B(n_4310),
.Y(n_18540)
);

OAI21xp5_ASAP7_75t_L g18541 ( 
.A1(n_18497),
.A2(n_4311),
.B(n_4312),
.Y(n_18541)
);

OAI22xp5_ASAP7_75t_L g18542 ( 
.A1(n_18508),
.A2(n_4314),
.B1(n_4312),
.B2(n_4313),
.Y(n_18542)
);

OAI21xp5_ASAP7_75t_L g18543 ( 
.A1(n_18493),
.A2(n_4313),
.B(n_4315),
.Y(n_18543)
);

OA21x2_ASAP7_75t_L g18544 ( 
.A1(n_18511),
.A2(n_4323),
.B(n_4315),
.Y(n_18544)
);

OA21x2_ASAP7_75t_L g18545 ( 
.A1(n_18518),
.A2(n_18514),
.B(n_18516),
.Y(n_18545)
);

HB1xp67_ASAP7_75t_L g18546 ( 
.A(n_18490),
.Y(n_18546)
);

NAND2xp5_ASAP7_75t_L g18547 ( 
.A(n_18519),
.B(n_4316),
.Y(n_18547)
);

INVx2_ASAP7_75t_L g18548 ( 
.A(n_18501),
.Y(n_18548)
);

CKINVDCx20_ASAP7_75t_R g18549 ( 
.A(n_18520),
.Y(n_18549)
);

OAI22xp5_ASAP7_75t_L g18550 ( 
.A1(n_18547),
.A2(n_18509),
.B1(n_18507),
.B2(n_18502),
.Y(n_18550)
);

OAI221xp5_ASAP7_75t_R g18551 ( 
.A1(n_18549),
.A2(n_18532),
.B1(n_18546),
.B2(n_18536),
.C(n_18545),
.Y(n_18551)
);

OR3x2_ASAP7_75t_L g18552 ( 
.A(n_18526),
.B(n_4316),
.C(n_4317),
.Y(n_18552)
);

HB1xp67_ASAP7_75t_L g18553 ( 
.A(n_18539),
.Y(n_18553)
);

OAI22xp5_ASAP7_75t_SL g18554 ( 
.A1(n_18548),
.A2(n_4320),
.B1(n_4321),
.B2(n_4319),
.Y(n_18554)
);

CKINVDCx20_ASAP7_75t_R g18555 ( 
.A(n_18528),
.Y(n_18555)
);

HB1xp67_ASAP7_75t_L g18556 ( 
.A(n_18544),
.Y(n_18556)
);

AOI22xp5_ASAP7_75t_L g18557 ( 
.A1(n_18534),
.A2(n_4322),
.B1(n_4318),
.B2(n_4319),
.Y(n_18557)
);

AND2x2_ASAP7_75t_L g18558 ( 
.A(n_18529),
.B(n_18527),
.Y(n_18558)
);

HB1xp67_ASAP7_75t_L g18559 ( 
.A(n_18538),
.Y(n_18559)
);

HB1xp67_ASAP7_75t_L g18560 ( 
.A(n_18523),
.Y(n_18560)
);

OAI22x1_ASAP7_75t_L g18561 ( 
.A1(n_18525),
.A2(n_18531),
.B1(n_18533),
.B2(n_18542),
.Y(n_18561)
);

OAI322xp33_ASAP7_75t_L g18562 ( 
.A1(n_18524),
.A2(n_4326),
.A3(n_4325),
.B1(n_4323),
.B2(n_4318),
.C1(n_4322),
.C2(n_4324),
.Y(n_18562)
);

OAI22x1_ASAP7_75t_L g18563 ( 
.A1(n_18535),
.A2(n_4326),
.B1(n_4324),
.B2(n_4325),
.Y(n_18563)
);

XNOR2x1_ASAP7_75t_L g18564 ( 
.A(n_18521),
.B(n_4561),
.Y(n_18564)
);

AOI22xp33_ASAP7_75t_L g18565 ( 
.A1(n_18537),
.A2(n_4329),
.B1(n_4327),
.B2(n_4328),
.Y(n_18565)
);

AND2x4_ASAP7_75t_L g18566 ( 
.A(n_18541),
.B(n_4329),
.Y(n_18566)
);

INVx2_ASAP7_75t_L g18567 ( 
.A(n_18552),
.Y(n_18567)
);

INVx1_ASAP7_75t_L g18568 ( 
.A(n_18556),
.Y(n_18568)
);

INVx1_ASAP7_75t_L g18569 ( 
.A(n_18560),
.Y(n_18569)
);

OAI21xp5_ASAP7_75t_L g18570 ( 
.A1(n_18559),
.A2(n_18540),
.B(n_18543),
.Y(n_18570)
);

AOI21xp5_ASAP7_75t_L g18571 ( 
.A1(n_18553),
.A2(n_18530),
.B(n_18522),
.Y(n_18571)
);

OAI21xp5_ASAP7_75t_L g18572 ( 
.A1(n_18550),
.A2(n_4328),
.B(n_4330),
.Y(n_18572)
);

AOI22xp5_ASAP7_75t_L g18573 ( 
.A1(n_18555),
.A2(n_4332),
.B1(n_4330),
.B2(n_4331),
.Y(n_18573)
);

BUFx2_ASAP7_75t_L g18574 ( 
.A(n_18558),
.Y(n_18574)
);

OAI22xp5_ASAP7_75t_L g18575 ( 
.A1(n_18564),
.A2(n_4333),
.B1(n_4331),
.B2(n_4332),
.Y(n_18575)
);

OAI22xp5_ASAP7_75t_L g18576 ( 
.A1(n_18565),
.A2(n_4335),
.B1(n_4333),
.B2(n_4334),
.Y(n_18576)
);

NAND2xp5_ASAP7_75t_SL g18577 ( 
.A(n_18561),
.B(n_4334),
.Y(n_18577)
);

AOI22xp5_ASAP7_75t_L g18578 ( 
.A1(n_18566),
.A2(n_4337),
.B1(n_4335),
.B2(n_4336),
.Y(n_18578)
);

OAI22xp5_ASAP7_75t_SL g18579 ( 
.A1(n_18568),
.A2(n_18569),
.B1(n_18567),
.B2(n_18574),
.Y(n_18579)
);

AOI21xp5_ASAP7_75t_L g18580 ( 
.A1(n_18571),
.A2(n_18570),
.B(n_18551),
.Y(n_18580)
);

BUFx3_ASAP7_75t_L g18581 ( 
.A(n_18576),
.Y(n_18581)
);

AOI21xp5_ASAP7_75t_L g18582 ( 
.A1(n_18577),
.A2(n_18557),
.B(n_18575),
.Y(n_18582)
);

OAI22xp5_ASAP7_75t_L g18583 ( 
.A1(n_18578),
.A2(n_18554),
.B1(n_18562),
.B2(n_18563),
.Y(n_18583)
);

OAI22xp5_ASAP7_75t_L g18584 ( 
.A1(n_18579),
.A2(n_18572),
.B1(n_18573),
.B2(n_4339),
.Y(n_18584)
);

OAI21xp5_ASAP7_75t_L g18585 ( 
.A1(n_18580),
.A2(n_4557),
.B(n_4556),
.Y(n_18585)
);

NOR2xp33_ASAP7_75t_L g18586 ( 
.A(n_18581),
.B(n_4336),
.Y(n_18586)
);

AOI22xp5_ASAP7_75t_L g18587 ( 
.A1(n_18583),
.A2(n_4340),
.B1(n_4341),
.B2(n_4339),
.Y(n_18587)
);

XNOR2xp5_ASAP7_75t_L g18588 ( 
.A(n_18582),
.B(n_4558),
.Y(n_18588)
);

NAND2xp5_ASAP7_75t_L g18589 ( 
.A(n_18580),
.B(n_4558),
.Y(n_18589)
);

INVx1_ASAP7_75t_L g18590 ( 
.A(n_18584),
.Y(n_18590)
);

AOI21xp5_ASAP7_75t_L g18591 ( 
.A1(n_18589),
.A2(n_4338),
.B(n_4340),
.Y(n_18591)
);

AOI22xp33_ASAP7_75t_L g18592 ( 
.A1(n_18585),
.A2(n_4342),
.B1(n_4338),
.B2(n_4341),
.Y(n_18592)
);

AOI22xp33_ASAP7_75t_L g18593 ( 
.A1(n_18588),
.A2(n_4345),
.B1(n_4343),
.B2(n_4344),
.Y(n_18593)
);

OAI21xp5_ASAP7_75t_L g18594 ( 
.A1(n_18590),
.A2(n_18591),
.B(n_18592),
.Y(n_18594)
);

NAND2xp5_ASAP7_75t_L g18595 ( 
.A(n_18593),
.B(n_18586),
.Y(n_18595)
);

INVxp67_ASAP7_75t_SL g18596 ( 
.A(n_18590),
.Y(n_18596)
);

OAI221xp5_ASAP7_75t_R g18597 ( 
.A1(n_18596),
.A2(n_18587),
.B1(n_4348),
.B2(n_4344),
.C(n_4347),
.Y(n_18597)
);

AOI22xp5_ASAP7_75t_SL g18598 ( 
.A1(n_18594),
.A2(n_4349),
.B1(n_4347),
.B2(n_4348),
.Y(n_18598)
);

INVxp67_ASAP7_75t_L g18599 ( 
.A(n_18595),
.Y(n_18599)
);

OR2x2_ASAP7_75t_L g18600 ( 
.A(n_18599),
.B(n_4349),
.Y(n_18600)
);

OA21x2_ASAP7_75t_L g18601 ( 
.A1(n_18597),
.A2(n_4350),
.B(n_4351),
.Y(n_18601)
);

INVx2_ASAP7_75t_L g18602 ( 
.A(n_18598),
.Y(n_18602)
);

AOI22xp5_ASAP7_75t_L g18603 ( 
.A1(n_18602),
.A2(n_4353),
.B1(n_4351),
.B2(n_4352),
.Y(n_18603)
);

OAI22xp5_ASAP7_75t_L g18604 ( 
.A1(n_18601),
.A2(n_4354),
.B1(n_4355),
.B2(n_4353),
.Y(n_18604)
);

AOI22xp5_ASAP7_75t_L g18605 ( 
.A1(n_18600),
.A2(n_4356),
.B1(n_4352),
.B2(n_4355),
.Y(n_18605)
);

AOI22xp5_ASAP7_75t_L g18606 ( 
.A1(n_18604),
.A2(n_4358),
.B1(n_4356),
.B2(n_4357),
.Y(n_18606)
);

AOI211xp5_ASAP7_75t_L g18607 ( 
.A1(n_18606),
.A2(n_18605),
.B(n_18603),
.C(n_4359),
.Y(n_18607)
);


endmodule