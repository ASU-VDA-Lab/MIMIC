module fake_jpeg_6429_n_300 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_42),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_53),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_4),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_61),
.B(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_18),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_4),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_33),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_70),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_99),
.Y(n_115)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_78),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_84),
.B1(n_93),
.B2(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_88),
.B(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_32),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_39),
.B1(n_29),
.B2(n_27),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_101),
.B1(n_107),
.B2(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_63),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_21),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_46),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_8),
.Y(n_129)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_116),
.Y(n_149)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_75),
.B(n_69),
.C(n_99),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_51),
.B1(n_66),
.B2(n_57),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_135),
.B1(n_138),
.B2(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_125),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_46),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_127),
.Y(n_164)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_129),
.Y(n_172)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_139),
.Y(n_146)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_10),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_86),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_54),
.C(n_63),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_82),
.A3(n_98),
.B1(n_70),
.B2(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_12),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_83),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_79),
.B1(n_100),
.B2(n_74),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_105),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_152),
.B(n_161),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_74),
.B1(n_85),
.B2(n_82),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_140),
.B1(n_115),
.B2(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_103),
.B1(n_85),
.B2(n_91),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_157),
.B1(n_142),
.B2(n_131),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_81),
.B(n_87),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_143),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_77),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_71),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_122),
.B(n_57),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_95),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_109),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_102),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_72),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_130),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_151),
.B1(n_54),
.B2(n_149),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_131),
.B1(n_139),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_182),
.A2(n_196),
.B1(n_198),
.B2(n_202),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_189),
.B1(n_192),
.B2(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_190),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_105),
.B1(n_67),
.B2(n_130),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_153),
.A2(n_150),
.B1(n_145),
.B2(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_90),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_203),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_204),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_145),
.B1(n_174),
.B2(n_168),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_144),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_147),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_164),
.B1(n_167),
.B2(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_132),
.B1(n_116),
.B2(n_112),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_146),
.B1(n_175),
.B2(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_136),
.B1(n_111),
.B2(n_92),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_173),
.B1(n_158),
.B2(n_162),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_169),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_214),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_172),
.B1(n_177),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_197),
.B(n_196),
.C(n_206),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_92),
.B(n_13),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_160),
.B1(n_158),
.B2(n_165),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_224),
.A2(n_229),
.B(n_191),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_151),
.B(n_148),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_186),
.B(n_178),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_201),
.C(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.C(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_201),
.C(n_179),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_243),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_247),
.B(n_213),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_202),
.C(n_182),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_192),
.A3(n_180),
.B1(n_178),
.B2(n_181),
.C1(n_73),
.C2(n_92),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_222),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_255),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_223),
.B1(n_217),
.B2(n_227),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_241),
.B1(n_236),
.B2(n_218),
.Y(n_264)
);

AOI321xp33_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_259),
.A3(n_225),
.B1(n_210),
.B2(n_247),
.C(n_218),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_258),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_216),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_210),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_217),
.C(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_268),
.B1(n_269),
.B2(n_223),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_233),
.C(n_234),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_270),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_236),
.B1(n_219),
.B2(n_232),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_223),
.B1(n_242),
.B2(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_12),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_281),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_259),
.C(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_275),
.C(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_261),
.C(n_253),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_255),
.C(n_166),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_264),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_13),
.B(n_14),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_13),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_291),
.B(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_279),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_283),
.B1(n_282),
.B2(n_288),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_16),
.B1(n_17),
.B2(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_283),
.C(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_291),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.C(n_16),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_298),
.Y(n_300)
);


endmodule