module fake_jpeg_19988_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_53),
.B1(n_37),
.B2(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_41),
.C(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_30),
.B1(n_21),
.B2(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_18),
.B1(n_22),
.B2(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_78),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_87),
.C(n_95),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_74),
.B1(n_27),
.B2(n_29),
.Y(n_130)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_75),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_37),
.B1(n_22),
.B2(n_38),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_40),
.B1(n_21),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_98),
.B1(n_102),
.B2(n_20),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_38),
.B(n_31),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_77),
.A2(n_24),
.B(n_2),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_93),
.B1(n_35),
.B2(n_27),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_86),
.B1(n_103),
.B2(n_27),
.Y(n_128)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_54),
.B1(n_55),
.B2(n_50),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_41),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_48),
.A2(n_20),
.B1(n_24),
.B2(n_41),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_116),
.B1(n_128),
.B2(n_130),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_35),
.B1(n_29),
.B2(n_26),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_121),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_35),
.C(n_28),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_36),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_125),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_36),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_93),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_1),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_112),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_69),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_146),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_66),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_143),
.Y(n_191)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_140),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_67),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_70),
.B(n_82),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_151),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_80),
.C(n_3),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_1),
.C(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_83),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_78),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_72),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_3),
.B(n_4),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_88),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_68),
.B1(n_96),
.B2(n_94),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_94),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_149),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_130),
.B1(n_125),
.B2(n_120),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_174),
.B1(n_178),
.B2(n_180),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_126),
.B(n_125),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_171),
.B(n_185),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_126),
.B(n_105),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_121),
.C(n_108),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_146),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_134),
.B1(n_106),
.B2(n_95),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_142),
.B1(n_154),
.B2(n_135),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_143),
.B(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_140),
.A2(n_134),
.B1(n_105),
.B2(n_117),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_107),
.B1(n_28),
.B2(n_17),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_28),
.B1(n_29),
.B2(n_26),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_153),
.B1(n_152),
.B2(n_160),
.Y(n_199)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_119),
.A3(n_81),
.B1(n_73),
.B2(n_26),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_158),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_202),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_137),
.B(n_148),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_199),
.B1(n_164),
.B2(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_136),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_211),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_171),
.B1(n_165),
.B2(n_179),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_138),
.B(n_147),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_199),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_229),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_201),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_187),
.B1(n_181),
.B2(n_178),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_232),
.B1(n_235),
.B2(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_184),
.B1(n_165),
.B2(n_170),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_185),
.B1(n_167),
.B2(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_17),
.B1(n_138),
.B2(n_6),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_119),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_17),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_240),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_221),
.B1(n_216),
.B2(n_228),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_204),
.C(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_247),
.C(n_249),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_248),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_207),
.B1(n_209),
.B2(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_233),
.B1(n_227),
.B2(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_217),
.C(n_200),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_206),
.C(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_213),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_254),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_195),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_250),
.B1(n_244),
.B2(n_210),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_221),
.B1(n_232),
.B2(n_219),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_261),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_216),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_223),
.C(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_251),
.C(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_208),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_203),
.B1(n_215),
.B2(n_251),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_272),
.A2(n_258),
.B1(n_256),
.B2(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_262),
.C(n_256),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_4),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_6),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_274),
.C(n_7),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_280),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_281),
.B(n_282),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_265),
.B(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

XOR2x2_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_286),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_275),
.B(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_285),
.C(n_288),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_282),
.B1(n_9),
.B2(n_10),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

OAI311xp33_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_6),
.A3(n_9),
.B1(n_10),
.C1(n_11),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_292),
.B(n_10),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_12),
.B(n_13),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_12),
.B(n_14),
.Y(n_297)
);


endmodule