module fake_aes_6970_n_1157 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1157);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1157;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_771;
wire n_696;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_703;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_928;
wire n_938;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_881;
wire n_806;
wire n_539;
wire n_1066;
wire n_1055;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_639;
wire n_376;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g264 ( .A(n_234), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_74), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_51), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_96), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_81), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_239), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_244), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_229), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_102), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_129), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_216), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_110), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_78), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_103), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_52), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_232), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_164), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_177), .Y(n_281) );
INVxp33_ASAP7_75t_L g282 ( .A(n_65), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_182), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_92), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_94), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_87), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_133), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_236), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_2), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_14), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_86), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_126), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_37), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_261), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_83), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_130), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_167), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_50), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_57), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_77), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_17), .Y(n_303) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_57), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_114), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_262), .Y(n_306) );
INVxp33_ASAP7_75t_SL g307 ( .A(n_128), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_171), .Y(n_308) );
BUFx2_ASAP7_75t_SL g309 ( .A(n_176), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_225), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_48), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_105), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_72), .Y(n_313) );
INVxp33_ASAP7_75t_SL g314 ( .A(n_112), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_11), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_127), .Y(n_317) );
INVxp33_ASAP7_75t_SL g318 ( .A(n_184), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_30), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_190), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_194), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_101), .Y(n_322) );
INVxp33_ASAP7_75t_SL g323 ( .A(n_27), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_260), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_185), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_211), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_75), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_85), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_44), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_27), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_7), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_16), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_32), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_115), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_53), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_146), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_205), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_64), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_9), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_98), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_49), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_131), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_189), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_246), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_157), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_36), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_49), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_152), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_42), .Y(n_350) );
INVxp33_ASAP7_75t_SL g351 ( .A(n_97), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_82), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_259), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_69), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_80), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_33), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_203), .Y(n_357) );
CKINVDCx14_ASAP7_75t_R g358 ( .A(n_77), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_137), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_50), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_66), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_119), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_16), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_46), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_30), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_150), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_52), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_142), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_123), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_1), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_60), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_104), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_230), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_8), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_139), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_220), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_81), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_214), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_51), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_29), .Y(n_380) );
CKINVDCx14_ASAP7_75t_R g381 ( .A(n_255), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_93), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_121), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_213), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_162), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_12), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_47), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_43), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_113), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_175), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_180), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_73), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_297), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_296), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_296), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_298), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_297), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_340), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_297), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_324), .A2(n_88), .B(n_84), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_298), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_340), .B(n_0), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_297), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_279), .Y(n_406) );
AND2x6_ASAP7_75t_L g407 ( .A(n_305), .B(n_89), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_305), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_306), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_349), .B(n_3), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_306), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_390), .A2(n_3), .B(n_4), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_297), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_349), .B(n_4), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_391), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_391), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_363), .B(n_5), .Y(n_420) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_329), .B(n_90), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_319), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_324), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_341), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_319), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_405), .B(n_424), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_405), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_409), .B(n_302), .C(n_301), .Y(n_428) );
BUFx8_ASAP7_75t_SL g429 ( .A(n_405), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_399), .B(n_304), .Y(n_433) );
AND2x6_ASAP7_75t_L g434 ( .A(n_403), .B(n_264), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_409), .B(n_345), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_399), .B(n_282), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_424), .B(n_331), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_400), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_409), .B(n_289), .Y(n_441) );
INVx8_ASAP7_75t_L g442 ( .A(n_407), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_396), .B(n_345), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_403), .A2(n_323), .B1(n_333), .B2(n_281), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_400), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_396), .B(n_366), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_403), .B(n_331), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_397), .B(n_366), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_394), .A2(n_323), .B1(n_281), .B2(n_312), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_395), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_395), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_400), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_400), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_420), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_397), .B(n_271), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_423), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_402), .B(n_377), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_400), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_406), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_400), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_402), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_408), .B(n_267), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_423), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_408), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_427), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_458), .B(n_416), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_426), .B(n_406), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_456), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_426), .B(n_416), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_426), .B(n_411), .Y(n_477) );
INVxp33_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_435), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_452), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_430), .A2(n_410), .B(n_413), .C(n_411), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_456), .Y(n_485) );
INVx8_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_430), .B(n_271), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_452), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_444), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_462), .B(n_420), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_453), .Y(n_492) );
INVx4_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_461), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_466), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_454), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_449), .B(n_394), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_467), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_467), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_434), .A2(n_407), .B1(n_412), .B2(n_410), .Y(n_503) );
NAND2x2_ASAP7_75t_L g504 ( .A(n_433), .B(n_307), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_470), .A2(n_413), .B(n_419), .C(n_418), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_434), .A2(n_421), .B1(n_418), .B2(n_419), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_442), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_462), .B(n_274), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_470), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_438), .B(n_278), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_438), .B(n_449), .Y(n_513) );
AND2x6_ASAP7_75t_SL g514 ( .A(n_439), .B(n_300), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_434), .A2(n_407), .B1(n_412), .B2(n_421), .Y(n_515) );
OR2x6_ASAP7_75t_L g516 ( .A(n_442), .B(n_309), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_449), .B(n_274), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_449), .B(n_308), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_434), .B(n_401), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_439), .B(n_308), .Y(n_523) );
AO22x1_ASAP7_75t_L g524 ( .A1(n_434), .A2(n_407), .B1(n_314), .B2(n_318), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_430), .B(n_325), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_433), .Y(n_526) );
CKINVDCx11_ASAP7_75t_R g527 ( .A(n_439), .Y(n_527) );
BUFx8_ASAP7_75t_L g528 ( .A(n_434), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_444), .B(n_311), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_439), .B(n_412), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_436), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_430), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_434), .A2(n_407), .B1(n_412), .B2(n_314), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_431), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_466), .Y(n_537) );
BUFx12f_ASAP7_75t_L g538 ( .A(n_431), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_451), .B(n_311), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_441), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_431), .B(n_338), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_436), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_431), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_437), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_437), .Y(n_545) );
AND3x2_ASAP7_75t_SL g546 ( .A(n_451), .B(n_365), .C(n_347), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_468), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_460), .B(n_285), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_437), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_437), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_443), .Y(n_551) );
AND2x6_ASAP7_75t_L g552 ( .A(n_468), .B(n_269), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_473), .B(n_459), .Y(n_553) );
CKINVDCx6p67_ASAP7_75t_R g554 ( .A(n_471), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_473), .B(n_459), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_483), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_479), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_539), .A2(n_300), .B1(n_342), .B2(n_312), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_551), .A2(n_326), .B1(n_327), .B2(n_283), .Y(n_560) );
OR2x6_ASAP7_75t_L g561 ( .A(n_486), .B(n_459), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_479), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_474), .B(n_459), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_473), .B(n_443), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_528), .B(n_283), .Y(n_566) );
BUFx12f_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_542), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_486), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_473), .A2(n_532), .B1(n_547), .B2(n_487), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_513), .B(n_448), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_538), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_528), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_526), .Y(n_575) );
INVx4_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
AOI21xp5_ASAP7_75t_SL g577 ( .A1(n_521), .A2(n_412), .B(n_448), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_531), .B(n_374), .C(n_334), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_486), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_476), .B(n_450), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_514), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_535), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_490), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_500), .A2(n_401), .B(n_450), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_497), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_497), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_516), .B(n_326), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_472), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_472), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_499), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_412), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_493), .B(n_301), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_480), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_498), .A2(n_428), .B1(n_318), .B2(n_351), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_499), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_498), .A2(n_428), .B1(n_351), .B2(n_307), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_481), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_481), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_508), .Y(n_605) );
O2A1O1Ixp5_ASAP7_75t_L g606 ( .A1(n_524), .A2(n_337), .B(n_384), .C(n_299), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_516), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
INVx6_ASAP7_75t_SL g609 ( .A(n_516), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_511), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_482), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_516), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_514), .Y(n_613) );
AND3x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_342), .C(n_313), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_506), .A2(n_327), .B1(n_381), .B2(n_321), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_477), .B(n_328), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_512), .Y(n_617) );
AO22x1_ASAP7_75t_L g618 ( .A1(n_478), .A2(n_350), .B1(n_354), .B2(n_328), .Y(n_618) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_537), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_484), .A2(n_401), .B(n_272), .Y(n_620) );
BUFx3_ASAP7_75t_L g621 ( .A(n_508), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_482), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_537), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_552), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_519), .B(n_350), .Y(n_625) );
INVx4_ASAP7_75t_L g626 ( .A(n_493), .Y(n_626) );
INVx3_ASAP7_75t_SL g627 ( .A(n_498), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_529), .B(n_354), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_511), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_492), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_540), .B(n_355), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_506), .A2(n_364), .B1(n_355), .B2(n_339), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_535), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_496), .Y(n_634) );
INVx4_ASAP7_75t_L g635 ( .A(n_493), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_492), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_529), .B(n_364), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_500), .A2(n_446), .B(n_445), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_520), .B(n_392), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_517), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_523), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_504), .A2(n_379), .B1(n_303), .B2(n_343), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_517), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_505), .A2(n_266), .B(n_268), .C(n_265), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_493), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_501), .A2(n_446), .B(n_445), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_496), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_496), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_494), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_475), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_530), .A2(n_290), .B1(n_291), .B2(n_276), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_509), .B(n_294), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_552), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_475), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_552), .B(n_530), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_475), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_485), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_485), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_543), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_548), .B(n_316), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_642), .A2(n_515), .B(n_534), .C(n_503), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_617), .B(n_546), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_617), .B(n_546), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_554), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_572), .B(n_552), .Y(n_665) );
INVx8_ASAP7_75t_L g666 ( .A(n_580), .Y(n_666) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_560), .Y(n_667) );
NAND2xp33_ASAP7_75t_L g668 ( .A(n_580), .B(n_496), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_578), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_572), .A2(n_552), .B1(n_504), .B2(n_521), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_568), .Y(n_671) );
INVx6_ASAP7_75t_L g672 ( .A(n_580), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_628), .B(n_552), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_628), .B(n_524), .Y(n_675) );
OAI21x1_ASAP7_75t_L g676 ( .A1(n_588), .A2(n_502), .B(n_501), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_580), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_572), .A2(n_521), .B1(n_495), .B2(n_485), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_556), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_575), .Y(n_680) );
CKINVDCx14_ASAP7_75t_R g681 ( .A(n_567), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_557), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_557), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_637), .B(n_422), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_565), .A2(n_570), .B1(n_592), .B2(n_598), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_562), .Y(n_686) );
INVx6_ASAP7_75t_L g687 ( .A(n_580), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_616), .B(n_495), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_562), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_584), .A2(n_522), .B1(n_330), .B2(n_348), .Y(n_690) );
AO31x2_ASAP7_75t_L g691 ( .A1(n_593), .A2(n_398), .A3(n_404), .B(n_393), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_644), .A2(n_336), .B(n_356), .C(n_352), .Y(n_692) );
INVx4_ASAP7_75t_L g693 ( .A(n_592), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_616), .A2(n_522), .B1(n_361), .B2(n_367), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_637), .B(n_422), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_571), .B(n_502), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_566), .A2(n_332), .B1(n_365), .B2(n_347), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_597), .A2(n_370), .B1(n_371), .B2(n_360), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_559), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_600), .A2(n_380), .B1(n_388), .B2(n_387), .C(n_386), .Y(n_700) );
BUFx2_ASAP7_75t_SL g701 ( .A(n_576), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g702 ( .A(n_567), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_641), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_594), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_615), .A2(n_332), .B1(n_423), .B2(n_425), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_558), .A2(n_425), .B1(n_423), .B2(n_525), .C(n_488), .Y(n_706) );
BUFx12f_ASAP7_75t_L g707 ( .A(n_582), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_652), .A2(n_541), .B1(n_518), .B2(n_510), .C(n_273), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_597), .A2(n_309), .B1(n_543), .B2(n_533), .Y(n_709) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_627), .A2(n_362), .B1(n_275), .B2(n_277), .C1(n_280), .C2(n_284), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_599), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_559), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_603), .A2(n_543), .B1(n_545), .B2(n_533), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_575), .A2(n_343), .B1(n_344), .B2(n_338), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_604), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_611), .A2(n_543), .B1(n_549), .B2(n_545), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_579), .A2(n_510), .B1(n_518), .B2(n_270), .C(n_385), .Y(n_717) );
OAI21x1_ASAP7_75t_L g718 ( .A1(n_620), .A2(n_544), .B(n_550), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_622), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_553), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_598), .A2(n_507), .B1(n_536), .B2(n_496), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_553), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_581), .A2(n_550), .B(n_549), .Y(n_723) );
AO31x2_ASAP7_75t_L g724 ( .A1(n_630), .A2(n_398), .A3(n_404), .B(n_393), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_636), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_576), .B(n_507), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_571), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_627), .B(n_344), .Y(n_728) );
INVx3_ASAP7_75t_L g729 ( .A(n_626), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_587), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_649), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_602), .B(n_357), .Y(n_732) );
BUFx4_ASAP7_75t_R g733 ( .A(n_609), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_651), .A2(n_544), .B1(n_536), .B2(n_287), .Y(n_734) );
BUFx4f_ASAP7_75t_SL g735 ( .A(n_609), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_563), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_660), .A2(n_375), .B1(n_288), .B2(n_292), .C(n_293), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_638), .A2(n_544), .B(n_295), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_553), .A2(n_536), .B1(n_310), .B2(n_315), .Y(n_739) );
BUFx12f_ASAP7_75t_L g740 ( .A(n_582), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_625), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_587), .Y(n_742) );
INVx4_ASAP7_75t_SL g743 ( .A(n_559), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_639), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_577), .A2(n_317), .B(n_286), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_589), .A2(n_382), .B1(n_359), .B2(n_322), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_590), .Y(n_747) );
INVx4_ASAP7_75t_SL g748 ( .A(n_559), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_586), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_555), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_590), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_576), .B(n_320), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_626), .B(n_335), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_646), .A2(n_353), .B(n_346), .Y(n_754) );
CKINVDCx12_ASAP7_75t_R g755 ( .A(n_561), .Y(n_755) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_613), .A2(n_368), .B1(n_369), .B2(n_372), .C1(n_383), .C2(n_376), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_591), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_596), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_596), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_601), .Y(n_760) );
BUFx4_ASAP7_75t_R g761 ( .A(n_605), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_601), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_607), .A2(n_378), .B1(n_389), .B2(n_373), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_632), .B(n_5), .Y(n_764) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_569), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_614), .B(n_631), .Y(n_766) );
CKINVDCx11_ASAP7_75t_R g767 ( .A(n_569), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_610), .B(n_6), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_612), .A2(n_398), .B1(n_404), .B2(n_393), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_563), .Y(n_770) );
BUFx2_ASAP7_75t_R g771 ( .A(n_563), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_612), .A2(n_398), .B1(n_404), .B2(n_393), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_662), .A2(n_655), .B1(n_624), .B2(n_653), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_677), .B(n_574), .Y(n_774) );
INVx5_ASAP7_75t_SL g775 ( .A(n_726), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_680), .B(n_573), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_671), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g778 ( .A1(n_744), .A2(n_618), .B1(n_624), .B2(n_653), .C1(n_573), .C2(n_629), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_663), .A2(n_643), .B1(n_640), .B2(n_564), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_766), .B(n_585), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_684), .B(n_640), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_703), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_667), .A2(n_643), .B1(n_654), .B2(n_650), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_682), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_705), .A2(n_657), .B1(n_658), .B2(n_656), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_695), .B(n_577), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_669), .Y(n_787) );
BUFx4f_ASAP7_75t_SL g788 ( .A(n_664), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_693), .A2(n_635), .B1(n_645), .B2(n_626), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_700), .A2(n_606), .B1(n_585), .B2(n_595), .C(n_608), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_679), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_661), .A2(n_619), .B(n_595), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_705), .A2(n_585), .B1(n_608), .B2(n_595), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_685), .A2(n_608), .B1(n_659), .B2(n_633), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_675), .A2(n_633), .B1(n_659), .B2(n_645), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_682), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_693), .B(n_635), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_741), .A2(n_645), .B1(n_635), .B2(n_623), .C(n_583), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_673), .A2(n_569), .B1(n_561), .B2(n_605), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_714), .B(n_6), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_761), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_704), .Y(n_802) );
OAI31xp33_ASAP7_75t_SL g803 ( .A1(n_697), .A2(n_414), .A3(n_9), .B(n_7), .Y(n_803) );
AOI21x1_ASAP7_75t_L g804 ( .A1(n_745), .A2(n_414), .B(n_561), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_681), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_702), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_676), .A2(n_414), .B(n_445), .Y(n_807) );
AO31x2_ASAP7_75t_L g808 ( .A1(n_683), .A2(n_414), .A3(n_447), .B(n_446), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_692), .A2(n_623), .B1(n_583), .B2(n_621), .C(n_378), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_767), .Y(n_810) );
CKINVDCx6p67_ASAP7_75t_R g811 ( .A(n_674), .Y(n_811) );
BUFx4f_ASAP7_75t_SL g812 ( .A(n_749), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_764), .A2(n_583), .B1(n_621), .B2(n_623), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_674), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_697), .A2(n_583), .B1(n_623), .B2(n_647), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_732), .B(n_8), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_670), .A2(n_648), .B1(n_647), .B2(n_569), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_728), .B(n_10), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_694), .A2(n_378), .B1(n_389), .B2(n_648), .C(n_634), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_711), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_718), .A2(n_457), .B(n_447), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_670), .B(n_13), .Y(n_822) );
OAI211xp5_ASAP7_75t_SL g823 ( .A1(n_756), .A2(n_447), .B(n_457), .C(n_463), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_746), .A2(n_561), .B1(n_634), .B2(n_389), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_701), .A2(n_634), .B1(n_389), .B2(n_415), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_735), .A2(n_634), .B1(n_417), .B2(n_415), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_737), .A2(n_417), .B1(n_415), .B2(n_457), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_746), .A2(n_417), .B1(n_415), .B2(n_463), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_698), .A2(n_417), .B1(n_415), .B2(n_440), .Y(n_829) );
AOI222xp33_ASAP7_75t_L g830 ( .A1(n_717), .A2(n_415), .B1(n_417), .B2(n_18), .C1(n_19), .C2(n_20), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_678), .A2(n_415), .B1(n_417), .B2(n_18), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_666), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_688), .A2(n_15), .B1(n_17), .B2(n_21), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_710), .B(n_21), .Y(n_834) );
OR2x2_ASAP7_75t_SL g835 ( .A(n_672), .B(n_22), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_715), .Y(n_836) );
NAND2x1_ASAP7_75t_L g837 ( .A(n_672), .B(n_417), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_720), .A2(n_465), .B1(n_455), .B2(n_440), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_719), .B(n_22), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_720), .A2(n_465), .B1(n_455), .B2(n_440), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_707), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_740), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_690), .B(n_23), .Y(n_843) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_666), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_722), .A2(n_465), .B1(n_455), .B2(n_440), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_678), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_846) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_765), .B(n_440), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_722), .A2(n_465), .B1(n_455), .B2(n_440), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_725), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_750), .A2(n_465), .B1(n_455), .B2(n_31), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_739), .A2(n_26), .B1(n_28), .B2(n_31), .Y(n_851) );
INVx6_ASAP7_75t_L g852 ( .A(n_666), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_750), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_731), .A2(n_665), .B1(n_690), .B2(n_753), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_677), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_855) );
INVx1_ASAP7_75t_SL g856 ( .A(n_771), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_683), .Y(n_857) );
INVx2_ASAP7_75t_SL g858 ( .A(n_672), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_752), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_755), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_860) );
OAI221xp5_ASAP7_75t_SL g861 ( .A1(n_706), .A2(n_44), .B1(n_45), .B2(n_46), .C(n_47), .Y(n_861) );
OAI211xp5_ASAP7_75t_SL g862 ( .A1(n_736), .A2(n_45), .B(n_48), .C(n_53), .Y(n_862) );
INVx6_ASAP7_75t_L g863 ( .A(n_743), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_757), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_743), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_758), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_760), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_708), .A2(n_58), .B1(n_59), .B2(n_61), .C(n_62), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_770), .Y(n_869) );
BUFx12f_ASAP7_75t_L g870 ( .A(n_687), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_733), .B(n_63), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_739), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_768), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_709), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_874) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_734), .A2(n_68), .B1(n_70), .B2(n_71), .C1(n_72), .C2(n_73), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_726), .A2(n_70), .B1(n_71), .B2(n_74), .Y(n_876) );
CKINVDCx14_ASAP7_75t_R g877 ( .A(n_687), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_834), .B(n_686), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_784), .Y(n_879) );
NOR2x1p5_ASAP7_75t_L g880 ( .A(n_810), .B(n_729), .Y(n_880) );
INVxp67_ASAP7_75t_L g881 ( .A(n_791), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_782), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_803), .A2(n_709), .B1(n_734), .B2(n_763), .C(n_772), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_861), .A2(n_763), .B1(n_769), .B2(n_723), .C(n_762), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_777), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_786), .A2(n_727), .B1(n_762), .B2(n_686), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_780), .B(n_761), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_854), .A2(n_713), .B1(n_716), .B2(n_687), .C(n_699), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_871), .A2(n_730), .B1(n_759), .B2(n_689), .Y(n_889) );
OAI22xp5_ASAP7_75t_SL g890 ( .A1(n_805), .A2(n_712), .B1(n_765), .B2(n_751), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_802), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g892 ( .A1(n_854), .A2(n_712), .B1(n_727), .B2(n_747), .C(n_742), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_835), .A2(n_747), .B1(n_696), .B2(n_765), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_781), .B(n_75), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_871), .A2(n_721), .B1(n_696), .B2(n_668), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_820), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_868), .A2(n_765), .B1(n_754), .B2(n_724), .C(n_691), .Y(n_897) );
OA21x2_ASAP7_75t_L g898 ( .A1(n_821), .A2(n_738), .B(n_724), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_787), .B(n_76), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_796), .Y(n_900) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_875), .B(n_724), .C(n_691), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_857), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_836), .Y(n_903) );
INVxp67_ASAP7_75t_L g904 ( .A(n_801), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_846), .A2(n_691), .B1(n_79), .B2(n_748), .C(n_99), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_843), .A2(n_748), .B1(n_691), .B2(n_100), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_830), .A2(n_91), .B1(n_95), .B2(n_106), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_779), .A2(n_107), .B1(n_108), .B2(n_109), .C(n_111), .Y(n_908) );
INVx4_ASAP7_75t_L g909 ( .A(n_852), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_849), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_800), .B(n_116), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_818), .B(n_117), .Y(n_912) );
AND2x6_ASAP7_75t_L g913 ( .A(n_775), .B(n_118), .Y(n_913) );
INVx3_ASAP7_75t_L g914 ( .A(n_852), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_864), .Y(n_915) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_779), .A2(n_120), .B1(n_122), .B2(n_124), .C(n_125), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_816), .A2(n_132), .B1(n_134), .B2(n_135), .Y(n_917) );
INVx1_ASAP7_75t_SL g918 ( .A(n_812), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_776), .B(n_136), .Y(n_919) );
OAI21xp5_ASAP7_75t_L g920 ( .A1(n_792), .A2(n_138), .B(n_140), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g921 ( .A1(n_828), .A2(n_141), .B(n_143), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_788), .B(n_144), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_839), .Y(n_923) );
AOI211xp5_ASAP7_75t_SL g924 ( .A1(n_865), .A2(n_145), .B(n_147), .C(n_148), .Y(n_924) );
OAI33xp33_ASAP7_75t_L g925 ( .A1(n_844), .A2(n_149), .A3(n_151), .B1(n_153), .B2(n_154), .B3(n_155), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_822), .A2(n_156), .B1(n_158), .B2(n_159), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_847), .A2(n_160), .B(n_161), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_877), .B(n_163), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_775), .B(n_165), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_793), .A2(n_166), .B1(n_168), .B2(n_169), .C(n_170), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_873), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_851), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_832), .B(n_778), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_793), .A2(n_178), .B1(n_179), .B2(n_181), .C(n_183), .Y(n_934) );
INVx3_ASAP7_75t_L g935 ( .A(n_852), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g936 ( .A1(n_824), .A2(n_186), .B(n_187), .C(n_188), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_794), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_870), .Y(n_938) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_863), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_785), .B(n_195), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_797), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_859), .B(n_199), .Y(n_942) );
AOI21xp5_ASAP7_75t_L g943 ( .A1(n_794), .A2(n_200), .B(n_202), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_862), .A2(n_204), .B1(n_206), .B2(n_207), .Y(n_944) );
BUFx3_ASAP7_75t_L g945 ( .A(n_811), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_872), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_946) );
AO31x2_ASAP7_75t_L g947 ( .A1(n_831), .A2(n_212), .A3(n_215), .B(n_217), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_876), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_785), .A2(n_218), .B1(n_219), .B2(n_222), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_855), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_860), .A2(n_223), .B1(n_224), .B2(n_226), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_833), .A2(n_227), .B1(n_228), .B2(n_231), .C(n_233), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_808), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_814), .B(n_237), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_874), .A2(n_238), .B1(n_240), .B2(n_241), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_808), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_815), .A2(n_242), .B1(n_243), .B2(n_245), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_808), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_859), .A2(n_247), .B(n_248), .C(n_249), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_869), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_815), .A2(n_250), .B1(n_251), .B2(n_252), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_853), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_807), .A2(n_253), .B(n_254), .Y(n_963) );
AOI31xp33_ASAP7_75t_L g964 ( .A1(n_856), .A2(n_256), .A3(n_257), .B(n_258), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_866), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_866), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_882), .B(n_773), .Y(n_967) );
AND2x4_ASAP7_75t_SL g968 ( .A(n_909), .B(n_774), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_899), .B(n_867), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_953), .B(n_774), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_885), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_923), .A2(n_867), .B1(n_874), .B2(n_783), .C(n_850), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_956), .B(n_795), .Y(n_973) );
AOI33xp33_ASAP7_75t_L g974 ( .A1(n_891), .A2(n_850), .A3(n_783), .B1(n_795), .B2(n_827), .B3(n_789), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_896), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_928), .B(n_858), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_903), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_910), .B(n_817), .Y(n_978) );
INVx1_ASAP7_75t_SL g979 ( .A(n_938), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_920), .A2(n_804), .B(n_799), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_881), .B(n_817), .Y(n_981) );
OAI21xp33_ASAP7_75t_SL g982 ( .A1(n_964), .A2(n_798), .B(n_813), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_948), .A2(n_790), .B1(n_827), .B2(n_823), .C(n_809), .Y(n_983) );
AOI33xp33_ASAP7_75t_L g984 ( .A1(n_960), .A2(n_829), .A3(n_813), .B1(n_826), .B2(n_825), .B3(n_819), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_958), .Y(n_985) );
INVx1_ASAP7_75t_SL g986 ( .A(n_918), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_915), .Y(n_987) );
INVx1_ASAP7_75t_SL g988 ( .A(n_945), .Y(n_988) );
OAI33xp33_ASAP7_75t_L g989 ( .A1(n_950), .A2(n_842), .A3(n_841), .B1(n_806), .B2(n_863), .B3(n_829), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_900), .B(n_837), .Y(n_990) );
AND4x1_ASAP7_75t_L g991 ( .A(n_922), .B(n_838), .C(n_840), .D(n_845), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_902), .B(n_848), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_879), .Y(n_993) );
AOI32xp33_ASAP7_75t_L g994 ( .A1(n_887), .A2(n_848), .A3(n_911), .B1(n_893), .B2(n_942), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_933), .B(n_962), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_907), .A2(n_887), .B1(n_889), .B2(n_883), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_909), .B(n_912), .Y(n_997) );
OAI33xp33_ASAP7_75t_L g998 ( .A1(n_951), .A2(n_904), .A3(n_966), .B1(n_965), .B2(n_932), .B3(n_890), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_906), .A2(n_944), .B1(n_926), .B2(n_895), .C(n_917), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_880), .B(n_935), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_901), .A2(n_951), .B1(n_904), .B2(n_925), .C(n_897), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_925), .A2(n_905), .B1(n_888), .B2(n_886), .C(n_892), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_954), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_939), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_914), .B(n_929), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_898), .Y(n_1006) );
NAND2xp5_ASAP7_75t_SL g1007 ( .A(n_886), .B(n_921), .Y(n_1007) );
INVx4_ASAP7_75t_L g1008 ( .A(n_913), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_939), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_939), .B(n_919), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g1011 ( .A(n_924), .B(n_926), .C(n_917), .D(n_955), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_963), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_939), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_947), .B(n_940), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_913), .Y(n_1015) );
OAI31xp33_ASAP7_75t_SL g1016 ( .A1(n_959), .A2(n_949), .A3(n_908), .B(n_916), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_913), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_913), .A2(n_884), .B1(n_952), .B2(n_946), .Y(n_1018) );
INVx4_ASAP7_75t_L g1019 ( .A(n_963), .Y(n_1019) );
NAND2xp33_ASAP7_75t_SL g1020 ( .A(n_931), .B(n_946), .Y(n_1020) );
OAI221xp5_ASAP7_75t_L g1021 ( .A1(n_931), .A2(n_930), .B1(n_934), .B2(n_941), .C(n_936), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_947), .Y(n_1022) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_947), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_943), .B(n_937), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_927), .B(n_957), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_961), .B(n_881), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_894), .B(n_878), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_894), .B(n_878), .Y(n_1028) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_900), .Y(n_1029) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_900), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1029), .B(n_985), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_971), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_973), .B(n_1023), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_975), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_995), .B(n_977), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_968), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_987), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1022), .B(n_1030), .Y(n_1038) );
INVx6_ASAP7_75t_L g1039 ( .A(n_1008), .Y(n_1039) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_1008), .B(n_1015), .Y(n_1040) );
INVxp33_ASAP7_75t_L g1041 ( .A(n_997), .Y(n_1041) );
INVx3_ASAP7_75t_L g1042 ( .A(n_970), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1022), .B(n_970), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_982), .A2(n_1018), .B(n_1011), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_993), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_970), .B(n_1006), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1006), .B(n_1028), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1027), .B(n_967), .Y(n_1048) );
AND2x4_ASAP7_75t_L g1049 ( .A(n_1015), .B(n_1017), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_978), .B(n_981), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_992), .B(n_990), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_1010), .B(n_1009), .Y(n_1052) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_979), .B(n_986), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1012), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1019), .Y(n_1055) );
OR2x2_ASAP7_75t_L g1056 ( .A(n_1014), .B(n_1026), .Y(n_1056) );
AOI221x1_ASAP7_75t_L g1057 ( .A1(n_1020), .A2(n_1003), .B1(n_1004), .B2(n_1013), .C(n_996), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1019), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_969), .B(n_1019), .Y(n_1059) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_1020), .A2(n_1007), .B(n_999), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1005), .B(n_980), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_980), .B(n_1001), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_968), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_976), .B(n_972), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1007), .B(n_1002), .Y(n_1065) );
NOR2x1_ASAP7_75t_L g1066 ( .A(n_1000), .B(n_988), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1025), .Y(n_1067) );
INVx1_ASAP7_75t_SL g1068 ( .A(n_1025), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1025), .B(n_974), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1024), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_1021), .B(n_989), .Y(n_1071) );
NOR2x1_ASAP7_75t_L g1072 ( .A(n_991), .B(n_998), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_998), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_984), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_983), .A2(n_994), .B1(n_1016), .B2(n_984), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1029), .B(n_1030), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1029), .B(n_985), .Y(n_1077) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_1036), .Y(n_1078) );
AOI21xp5_ASAP7_75t_L g1079 ( .A1(n_1060), .A2(n_1044), .B(n_1057), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1032), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1075), .A2(n_1036), .B1(n_1063), .B2(n_1071), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1047), .B(n_1059), .Y(n_1082) );
INVxp67_ASAP7_75t_L g1083 ( .A(n_1066), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1032), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1034), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1034), .Y(n_1086) );
AOI211x1_ASAP7_75t_L g1087 ( .A1(n_1065), .A2(n_1074), .B(n_1064), .C(n_1035), .Y(n_1087) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_1039), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1048), .B(n_1065), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1050), .B(n_1047), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1051), .B(n_1050), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_1067), .B(n_1068), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1070), .B(n_1069), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1070), .B(n_1069), .Y(n_1094) );
INVx3_ASAP7_75t_L g1095 ( .A(n_1039), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1056), .B(n_1051), .Y(n_1096) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_1063), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_1041), .B(n_1072), .Y(n_1098) );
AND2x4_ASAP7_75t_SL g1099 ( .A(n_1040), .B(n_1042), .Y(n_1099) );
INVx3_ASAP7_75t_L g1100 ( .A(n_1039), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1045), .B(n_1037), .Y(n_1101) );
NAND3xp33_ASAP7_75t_SL g1102 ( .A(n_1053), .B(n_1062), .C(n_1073), .Y(n_1102) );
AND2x4_ASAP7_75t_L g1103 ( .A(n_1067), .B(n_1049), .Y(n_1103) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_1073), .B(n_1056), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1096), .B(n_1076), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1080), .Y(n_1106) );
INVx1_ASAP7_75t_SL g1107 ( .A(n_1078), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1084), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1104), .B(n_1059), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1082), .B(n_1061), .Y(n_1110) );
XOR2x2_ASAP7_75t_L g1111 ( .A(n_1087), .B(n_1049), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1091), .B(n_1038), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1090), .B(n_1031), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1093), .B(n_1033), .Y(n_1114) );
INVx1_ASAP7_75t_SL g1115 ( .A(n_1097), .Y(n_1115) );
NAND4xp25_ASAP7_75t_L g1116 ( .A(n_1079), .B(n_1049), .C(n_1052), .D(n_1058), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1101), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1094), .B(n_1052), .Y(n_1118) );
XOR2x2_ASAP7_75t_L g1119 ( .A(n_1081), .B(n_1031), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1103), .B(n_1046), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1085), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1122 ( .A1(n_1083), .A2(n_1039), .B1(n_1040), .B2(n_1042), .Y(n_1122) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_1099), .Y(n_1123) );
XNOR2xp5_ASAP7_75t_L g1124 ( .A(n_1089), .B(n_1040), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g1125 ( .A(n_1098), .Y(n_1125) );
INVx2_ASAP7_75t_SL g1126 ( .A(n_1099), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1086), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_1102), .A2(n_1043), .B1(n_1046), .B2(n_1077), .Y(n_1128) );
NAND2xp33_ASAP7_75t_L g1129 ( .A(n_1088), .B(n_1055), .Y(n_1129) );
NOR3x1_ASAP7_75t_L g1130 ( .A(n_1088), .B(n_1054), .C(n_1055), .Y(n_1130) );
INVx1_ASAP7_75t_SL g1131 ( .A(n_1095), .Y(n_1131) );
NOR2x1_ASAP7_75t_L g1132 ( .A(n_1116), .B(n_1107), .Y(n_1132) );
AOI21xp5_ASAP7_75t_L g1133 ( .A1(n_1119), .A2(n_1111), .B(n_1129), .Y(n_1133) );
NOR3xp33_ASAP7_75t_L g1134 ( .A(n_1125), .B(n_1122), .C(n_1115), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1110), .B(n_1120), .Y(n_1135) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_1123), .Y(n_1136) );
OA22x2_ASAP7_75t_L g1137 ( .A1(n_1123), .A2(n_1126), .B1(n_1124), .B2(n_1128), .Y(n_1137) );
AOI221x1_ASAP7_75t_L g1138 ( .A1(n_1133), .A2(n_1117), .B1(n_1109), .B2(n_1106), .C(n_1121), .Y(n_1138) );
AOI22xp33_ASAP7_75t_SL g1139 ( .A1(n_1137), .A2(n_1100), .B1(n_1095), .B2(n_1131), .Y(n_1139) );
AOI21xp5_ASAP7_75t_L g1140 ( .A1(n_1132), .A2(n_1105), .B(n_1118), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1136), .Y(n_1141) );
NAND4xp25_ASAP7_75t_L g1142 ( .A(n_1134), .B(n_1130), .C(n_1100), .D(n_1092), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1141), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_1139), .A2(n_1112), .B1(n_1113), .B2(n_1135), .Y(n_1144) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_1142), .A2(n_1140), .B1(n_1138), .B2(n_1114), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1143), .Y(n_1146) );
NOR3xp33_ASAP7_75t_L g1147 ( .A(n_1144), .B(n_1127), .C(n_1108), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1145), .B(n_1127), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1146), .Y(n_1149) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_1148), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1149), .Y(n_1151) );
INVxp67_ASAP7_75t_SL g1152 ( .A(n_1150), .Y(n_1152) );
HB1xp67_ASAP7_75t_L g1153 ( .A(n_1151), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1151), .Y(n_1154) );
XNOR2xp5_ASAP7_75t_L g1155 ( .A(n_1152), .B(n_1147), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1153), .Y(n_1156) );
AOI21xp5_ASAP7_75t_L g1157 ( .A1(n_1156), .A2(n_1155), .B(n_1154), .Y(n_1157) );
endmodule