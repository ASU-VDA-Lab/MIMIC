module fake_jpeg_13193_n_587 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_587);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_587;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_64),
.Y(n_185)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_65),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_80),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_90),
.Y(n_137)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_8),
.C(n_16),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_24),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_35),
.B(n_8),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_108),
.B(n_53),
.Y(n_156)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_26),
.B(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_14),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_115),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_35),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_117),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_32),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_84),
.A2(n_45),
.B1(n_25),
.B2(n_33),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_131),
.A2(n_134),
.B(n_135),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_58),
.A2(n_45),
.B1(n_33),
.B2(n_50),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_33),
.B1(n_50),
.B2(n_53),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_145),
.B1(n_151),
.B2(n_167),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g241 ( 
.A(n_138),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_140),
.B(n_144),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_54),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_48),
.B1(n_51),
.B2(n_44),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_53),
.B1(n_51),
.B2(n_48),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_19),
.B1(n_44),
.B2(n_30),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_49),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_102),
.A2(n_55),
.B1(n_54),
.B2(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_37),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_181),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_80),
.A2(n_19),
.B1(n_30),
.B2(n_38),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_56),
.A2(n_24),
.B1(n_36),
.B2(n_38),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_75),
.A2(n_55),
.B1(n_40),
.B2(n_37),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_82),
.A2(n_49),
.B1(n_47),
.B2(n_52),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_72),
.B(n_40),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_66),
.A2(n_36),
.B1(n_47),
.B2(n_52),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_94),
.B1(n_76),
.B2(n_78),
.Y(n_202)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_137),
.B(n_57),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_218),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_88),
.B1(n_74),
.B2(n_109),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_194),
.A2(n_133),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_134),
.A2(n_69),
.B1(n_71),
.B2(n_91),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_195),
.A2(n_212),
.B1(n_224),
.B2(n_237),
.Y(n_281)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_196),
.Y(n_280)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_198),
.Y(n_291)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_202),
.A2(n_243),
.B1(n_135),
.B2(n_151),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_100),
.B1(n_106),
.B2(n_104),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_169),
.B(n_65),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_204),
.B(n_211),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_223),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_206),
.Y(n_315)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

BUFx24_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_122),
.A2(n_89),
.B1(n_49),
.B2(n_57),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_210),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_113),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_136),
.A2(n_79),
.B1(n_81),
.B2(n_112),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_130),
.A2(n_185),
.B1(n_132),
.B2(n_49),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_213),
.A2(n_215),
.B1(n_256),
.B2(n_257),
.Y(n_267)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_130),
.A2(n_49),
.B1(n_103),
.B2(n_111),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_123),
.B(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_220),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_10),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_167),
.A2(n_105),
.B1(n_113),
.B2(n_115),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_228),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_156),
.B(n_8),
.C(n_17),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_230),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_146),
.B(n_9),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_232),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_158),
.B(n_68),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_147),
.B(n_7),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_242),
.Y(n_277)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_235),
.Y(n_305)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_131),
.A2(n_99),
.B1(n_9),
.B2(n_12),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_142),
.Y(n_238)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_153),
.B(n_0),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_186),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_125),
.B1(n_155),
.B2(n_143),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_126),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_172),
.B(n_17),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_2),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_121),
.B(n_17),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_241),
.Y(n_270)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_128),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_252),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_190),
.A2(n_14),
.B1(n_9),
.B2(n_3),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_253),
.A2(n_143),
.B1(n_129),
.B2(n_180),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_254),
.Y(n_304)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_255),
.Y(n_317)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_259),
.B1(n_206),
.B2(n_254),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_185),
.A2(n_152),
.B1(n_191),
.B2(n_184),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_260),
.A2(n_4),
.B1(n_6),
.B2(n_214),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_273),
.B1(n_308),
.B2(n_194),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_220),
.B(n_1),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_269),
.B(n_287),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_270),
.B(n_279),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_209),
.B(n_176),
.C(n_154),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_276),
.C(n_253),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_208),
.B(n_125),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_283),
.A2(n_301),
.B1(n_302),
.B2(n_260),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_118),
.B(n_157),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_284),
.A2(n_287),
.B(n_260),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_225),
.A2(n_155),
.B1(n_129),
.B2(n_157),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_285),
.A2(n_296),
.B1(n_238),
.B2(n_245),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_222),
.A2(n_9),
.B(n_3),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_200),
.A2(n_154),
.B1(n_133),
.B2(n_180),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_294),
.B1(n_288),
.B2(n_302),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_199),
.A2(n_212),
.B1(n_242),
.B2(n_224),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_237),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_200),
.A2(n_222),
.B1(n_202),
.B2(n_194),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_2),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_279),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_323),
.B1(n_336),
.B2(n_339),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_277),
.B(n_236),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_326),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_197),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_320),
.B(n_331),
.C(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_194),
.B1(n_244),
.B2(n_226),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_295),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_324),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_298),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_277),
.B(n_239),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_303),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_327),
.B(n_349),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_250),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_257),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_235),
.C(n_251),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_358),
.Y(n_363)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_228),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_261),
.B(n_290),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_271),
.A2(n_226),
.B1(n_255),
.B2(n_217),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_278),
.B(n_216),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_352),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_301),
.A2(n_234),
.B1(n_240),
.B2(n_196),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_281),
.A2(n_256),
.B1(n_260),
.B2(n_227),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_340),
.A2(n_341),
.B1(n_304),
.B2(n_306),
.Y(n_385)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_344),
.A2(n_294),
.B1(n_300),
.B2(n_267),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_269),
.B(n_282),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_347),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_269),
.B(n_207),
.C(n_6),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_273),
.A2(n_6),
.B1(n_207),
.B2(n_281),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_348),
.A2(n_317),
.B1(n_289),
.B2(n_314),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_6),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_263),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_353),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_297),
.B(n_288),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_270),
.B(n_310),
.CI(n_284),
.CON(n_353),
.SN(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_303),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_354),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_357),
.A2(n_283),
.B1(n_286),
.B2(n_313),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_262),
.B(n_291),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_359),
.B(n_361),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_262),
.B(n_265),
.C(n_289),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_275),
.Y(n_394)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_265),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_291),
.B(n_317),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_362),
.A2(n_275),
.B(n_300),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_374),
.C(n_325),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_368),
.A2(n_382),
.B1(n_343),
.B2(n_402),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_362),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_354),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_293),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_362),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_379),
.B(n_384),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_348),
.B1(n_322),
.B2(n_321),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_324),
.B1(n_342),
.B2(n_329),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_275),
.B(n_314),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_387),
.A2(n_359),
.B(n_327),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_341),
.A2(n_306),
.B1(n_309),
.B2(n_304),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_388),
.A2(n_389),
.B1(n_393),
.B2(n_339),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_340),
.A2(n_309),
.B1(n_299),
.B2(n_286),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_391),
.A2(n_402),
.B1(n_333),
.B2(n_351),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_318),
.A2(n_313),
.B1(n_312),
.B2(n_280),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_360),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_319),
.B(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_396),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_326),
.B(n_305),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_275),
.B(n_312),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_280),
.B(n_272),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_323),
.A2(n_272),
.B1(n_266),
.B2(n_292),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_352),
.C(n_359),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_407),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_345),
.C(n_334),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_409),
.A2(n_423),
.B(n_429),
.Y(n_447)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_412),
.Y(n_446)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_337),
.C(n_356),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_416),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_414),
.A2(n_388),
.B1(n_393),
.B2(n_389),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_356),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_336),
.C(n_331),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_353),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_418),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_363),
.B(n_332),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_419),
.B(n_366),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_420),
.A2(n_430),
.B1(n_432),
.B2(n_391),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_347),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_378),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_367),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_425),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_398),
.A2(n_355),
.B(n_353),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_372),
.C(n_374),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_396),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_367),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_427),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_401),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_433),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_344),
.B(n_361),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_431),
.A2(n_436),
.B(n_376),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_346),
.B1(n_343),
.B2(n_350),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_377),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_397),
.B(n_346),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_434),
.B(n_437),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_R g457 ( 
.A(n_435),
.B(n_378),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_377),
.Y(n_437)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_431),
.A2(n_372),
.B1(n_390),
.B2(n_386),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_441),
.A2(n_445),
.B1(n_456),
.B2(n_429),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_399),
.B(n_387),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_442),
.A2(n_424),
.B(n_466),
.Y(n_479)
);

OA21x2_ASAP7_75t_SL g443 ( 
.A1(n_427),
.A2(n_392),
.B(n_383),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_443),
.B(n_454),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_417),
.A2(n_390),
.B1(n_371),
.B2(n_379),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_448),
.A2(n_428),
.B1(n_433),
.B2(n_437),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_459),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_423),
.A2(n_364),
.B(n_380),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_452),
.B(n_424),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_418),
.B(n_375),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_425),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_455),
.B(n_434),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_417),
.A2(n_395),
.B1(n_375),
.B2(n_366),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_413),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_461),
.C(n_465),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_403),
.B(n_400),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_376),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_400),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_468),
.C(n_426),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_266),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_471),
.A2(n_440),
.B(n_464),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_472),
.A2(n_464),
.B1(n_463),
.B2(n_461),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_456),
.B(n_466),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_481),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_490),
.Y(n_503)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_453),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_477),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g516 ( 
.A(n_479),
.B(n_480),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_442),
.A2(n_436),
.B(n_422),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_449),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_446),
.Y(n_484)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_446),
.Y(n_485)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_421),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_486),
.B(n_473),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_469),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_491),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_468),
.C(n_444),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_444),
.C(n_438),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_448),
.A2(n_416),
.B1(n_410),
.B2(n_406),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_462),
.A2(n_410),
.B1(n_405),
.B2(n_408),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_492),
.A2(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_462),
.A2(n_420),
.B1(n_412),
.B2(n_411),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_447),
.A2(n_430),
.B1(n_432),
.B2(n_366),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_447),
.B(n_292),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_495),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_452),
.A2(n_315),
.B1(n_441),
.B2(n_451),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_504),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_465),
.C(n_438),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_501),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_467),
.C(n_439),
.Y(n_501)
);

BUFx12f_ASAP7_75t_SL g502 ( 
.A(n_471),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_517),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_507),
.A2(n_518),
.B1(n_474),
.B2(n_494),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_490),
.B(n_439),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_476),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_458),
.C(n_315),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_515),
.C(n_495),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_475),
.B(n_473),
.C(n_491),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_472),
.A2(n_478),
.B1(n_485),
.B2(n_484),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_525),
.Y(n_538)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_504),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_515),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_498),
.B(n_479),
.C(n_478),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_534),
.C(n_519),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_480),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_535),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_510),
.A2(n_470),
.B1(n_483),
.B2(n_488),
.Y(n_529)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_505),
.A2(n_474),
.B(n_470),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_505),
.A2(n_482),
.B1(n_477),
.B2(n_474),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_536),
.Y(n_540)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_533),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_496),
.C(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_512),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_492),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_518),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_534),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_543),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_550),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_500),
.C(n_503),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_500),
.C(n_503),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_508),
.C(n_541),
.Y(n_563)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_546),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_530),
.A2(n_497),
.B1(n_513),
.B2(n_512),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_526),
.A2(n_516),
.B1(n_497),
.B2(n_502),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_551),
.A2(n_520),
.B1(n_516),
.B2(n_506),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_559),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_542),
.A2(n_527),
.B(n_513),
.Y(n_556)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_523),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_557),
.B(n_561),
.Y(n_571)
);

MAJx2_ASAP7_75t_L g559 ( 
.A(n_543),
.B(n_523),
.C(n_527),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_552),
.A2(n_509),
.B1(n_524),
.B2(n_537),
.Y(n_560)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_560),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_551),
.A2(n_528),
.B(n_509),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_544),
.B(n_536),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_562),
.B(n_563),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_549),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_564),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_558),
.B(n_539),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_570),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_553),
.B(n_540),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_548),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_SL g578 ( 
.A(n_573),
.B(n_556),
.C(n_547),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_563),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_574),
.Y(n_580)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_545),
.B(n_554),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_575),
.A2(n_577),
.B(n_578),
.Y(n_579)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_571),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_576),
.A2(n_567),
.B(n_569),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_572),
.B(n_547),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_582),
.B(n_583),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_580),
.B(n_566),
.C(n_559),
.Y(n_583)
);

BUFx24_ASAP7_75t_SL g585 ( 
.A(n_584),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_585),
.A2(n_560),
.B(n_579),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_586),
.B(n_566),
.Y(n_587)
);


endmodule