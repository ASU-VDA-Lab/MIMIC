module fake_netlist_6_3027_n_1254 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1254);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1254;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_46),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_39),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_36),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_86),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_90),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_9),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_146),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_56),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_28),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_85),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_66),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_83),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_20),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_75),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_64),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_80),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_166),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_131),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_141),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_96),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_110),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_67),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_54),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_20),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_162),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_24),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_177),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_87),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_143),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_76),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_158),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_52),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_109),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_144),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_120),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_134),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_97),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_95),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_31),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_72),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_149),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_126),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_98),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_163),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_51),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_165),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_122),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_49),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_171),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_82),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_160),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_147),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_152),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_164),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_142),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_172),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_178),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_91),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_57),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_32),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_48),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_136),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_47),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_224),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_R g303 ( 
.A(n_252),
.B(n_0),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_242),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_248),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_278),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_1),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_264),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_200),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_204),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_188),
.B(n_2),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_208),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_214),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_186),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_223),
.B(n_2),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_211),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_180),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_249),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_213),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_230),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_241),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_258),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_243),
.B(n_3),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_262),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_201),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_263),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_183),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_249),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_185),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_3),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_207),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_209),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_187),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_210),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_272),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_189),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_192),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_284),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_199),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_287),
.B(n_5),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_199),
.B(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_202),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_202),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_294),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_194),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_275),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_196),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_197),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_203),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_298),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_217),
.Y(n_377)
);

BUFx2_ASAP7_75t_SL g378 ( 
.A(n_280),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_280),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_220),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_179),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_283),
.Y(n_383)
);

BUFx6f_ASAP7_75t_SL g384 ( 
.A(n_286),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_212),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_228),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_233),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_245),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_251),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_179),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_310),
.B(n_181),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_181),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_190),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_190),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_314),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_182),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_193),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_339),
.A2(n_371),
.B1(n_326),
.B2(n_302),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_308),
.B(n_253),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_308),
.B(n_261),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_343),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_288),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_312),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_191),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_191),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_382),
.B(n_306),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_332),
.B(n_198),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_361),
.A2(n_296),
.B(n_205),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_370),
.B(n_198),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_366),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_240),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_373),
.B(n_240),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_319),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_351),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_374),
.B(n_206),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_377),
.B(n_269),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_238),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_323),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_380),
.B(n_267),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_269),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_317),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_317),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_346),
.B(n_270),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_325),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_381),
.B(n_215),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_327),
.B(n_286),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_325),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_328),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_321),
.B(n_330),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_328),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_329),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_402),
.B(n_331),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_457),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_402),
.A2(n_303),
.B1(n_365),
.B2(n_316),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_422),
.A2(n_316),
.B1(n_360),
.B2(n_376),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_414),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_399),
.B(n_414),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_327),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_393),
.B(n_321),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_404),
.B(n_357),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_420),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_404),
.B(n_357),
.Y(n_485)
);

AND3x1_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_369),
.C(n_307),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_457),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_453),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_453),
.A2(n_300),
.B1(n_347),
.B2(n_342),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_450),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_457),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

NOR2x1p5_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_368),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_453),
.B(n_424),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_404),
.A2(n_350),
.B1(n_320),
.B2(n_311),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_398),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_407),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_393),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_445),
.B(n_330),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_403),
.B(n_315),
.C(n_311),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_394),
.B(n_352),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_441),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_445),
.B(n_334),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_450),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_396),
.B(n_355),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_334),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_396),
.B(n_385),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_406),
.B(n_329),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_335),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_447),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_406),
.A2(n_445),
.B1(n_452),
.B2(n_411),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_424),
.A2(n_301),
.B(n_337),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_445),
.B(n_335),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_418),
.B(n_425),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_305),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_519),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_504),
.B(n_445),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_411),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_406),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_475),
.B(n_410),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_491),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_450),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_531),
.B(n_413),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_437),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_514),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

AO22x2_ASAP7_75t_L g545 ( 
.A1(n_461),
.A2(n_339),
.B1(n_397),
.B2(n_433),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_496),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_527),
.A2(n_424),
.B(n_439),
.C(n_437),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_496),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_324),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_413),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_514),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_485),
.B(n_426),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_492),
.B(n_437),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_503),
.B(n_436),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_492),
.B(n_426),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_517),
.B(n_439),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_523),
.A2(n_479),
.B1(n_497),
.B2(n_517),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_525),
.B(n_443),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_498),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_439),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_509),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_523),
.A2(n_458),
.B1(n_443),
.B2(n_453),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_446),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_525),
.B(n_395),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_480),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_523),
.A2(n_479),
.B1(n_497),
.B2(n_485),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_510),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_523),
.B(n_446),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_395),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_498),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_523),
.B(n_446),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_487),
.B(n_418),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_506),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_397),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_493),
.B(n_425),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_525),
.B(n_433),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_486),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_495),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_479),
.B(n_429),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_411),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_530),
.B(n_423),
.Y(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_479),
.A2(n_453),
.B1(n_429),
.B2(n_438),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_421),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_525),
.B(n_405),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_479),
.B(n_432),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_520),
.B(n_405),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_489),
.B(n_403),
.C(n_421),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_524),
.B(n_470),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_479),
.B(n_432),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_483),
.B(n_438),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_435),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_478),
.A2(n_304),
.B1(n_435),
.B2(n_338),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_500),
.B(n_405),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_483),
.B(n_408),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_483),
.B(n_408),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_476),
.B(n_336),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_512),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_500),
.B(n_408),
.Y(n_605)
);

O2A1O1Ixp5_ASAP7_75t_L g606 ( 
.A1(n_529),
.A2(n_522),
.B(n_528),
.C(n_512),
.Y(n_606)
);

BUFx8_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_464),
.B(n_441),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_522),
.B(n_408),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_528),
.B(n_408),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_408),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_499),
.B(n_408),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_500),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_500),
.B(n_419),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_484),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_500),
.B(n_419),
.Y(n_617)
);

BUFx6f_ASAP7_75t_SL g618 ( 
.A(n_476),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_503),
.B(n_336),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_476),
.A2(n_344),
.B1(n_338),
.B2(n_376),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_508),
.B(n_419),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_511),
.B(n_344),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_476),
.B(n_368),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_476),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_464),
.B(n_419),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_497),
.A2(n_292),
.B1(n_289),
.B2(n_285),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_497),
.A2(n_283),
.B1(n_441),
.B2(n_447),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_419),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_464),
.B(n_419),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_508),
.B(n_283),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_588),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_497),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_533),
.B(n_270),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_540),
.B(n_463),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_575),
.B(n_463),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_583),
.A2(n_502),
.B(n_516),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_572),
.B(n_274),
.C(n_273),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_502),
.B(n_516),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_596),
.A2(n_502),
.B(n_518),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_532),
.B(n_384),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_579),
.B(n_466),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_535),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_542),
.B(n_273),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_537),
.B(n_384),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_595),
.A2(n_481),
.B(n_466),
.C(n_467),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_595),
.A2(n_534),
.B1(n_535),
.B2(n_612),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_585),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_606),
.A2(n_529),
.B(n_471),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_543),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_538),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_551),
.B(n_467),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_591),
.A2(n_502),
.B(n_518),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_SL g656 ( 
.A(n_549),
.B(n_276),
.C(n_274),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_534),
.B(n_471),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_538),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_537),
.B(n_384),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_587),
.B(n_442),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_547),
.A2(n_481),
.B(n_477),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_569),
.A2(n_477),
.B(n_526),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_553),
.B(n_526),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_561),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_664)
);

O2A1O1Ixp5_ASAP7_75t_L g665 ( 
.A1(n_593),
.A2(n_473),
.B(n_468),
.C(n_469),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_562),
.B(n_484),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_556),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_564),
.B(n_276),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_585),
.B(n_442),
.Y(n_671)
);

CKINVDCx10_ASAP7_75t_R g672 ( 
.A(n_618),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_554),
.B(n_279),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_550),
.B(n_279),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_490),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_568),
.B(n_490),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_585),
.B(n_444),
.Y(n_677)
);

AO21x1_ASAP7_75t_L g678 ( 
.A1(n_593),
.A2(n_473),
.B(n_469),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_557),
.B(n_281),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_565),
.A2(n_501),
.B(n_494),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_620),
.B(n_341),
.C(n_340),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_570),
.B(n_494),
.Y(n_682)
);

OA22x2_ASAP7_75t_L g683 ( 
.A1(n_577),
.A2(n_541),
.B1(n_581),
.B2(n_544),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_539),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_624),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_541),
.B(n_281),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_546),
.B(n_501),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_546),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_548),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_571),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_548),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_560),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_556),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_600),
.A2(n_505),
.B(n_434),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_590),
.B(n_598),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_444),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_560),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_591),
.A2(n_415),
.B(n_419),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_589),
.B(n_282),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_582),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_608),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_576),
.B(n_505),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_L g704 ( 
.A1(n_622),
.A2(n_599),
.B(n_619),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_625),
.A2(n_455),
.B(n_449),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_597),
.B(n_449),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_559),
.B(n_282),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_559),
.B(n_285),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_566),
.B(n_289),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_588),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_566),
.B(n_292),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_580),
.B(n_226),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_573),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_449),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_628),
.A2(n_455),
.B(n_434),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_629),
.A2(n_455),
.B(n_434),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_558),
.A2(n_460),
.B1(n_459),
.B2(n_456),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_555),
.B(n_460),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_584),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_231),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_574),
.B(n_604),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_584),
.Y(n_722)
);

AOI21x1_ASAP7_75t_L g723 ( 
.A1(n_600),
.A2(n_431),
.B(n_416),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_627),
.A2(n_459),
.B(n_456),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_567),
.B(n_451),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_608),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_613),
.A2(n_431),
.B(n_427),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_617),
.A2(n_431),
.B(n_427),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_447),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_706),
.A2(n_602),
.B(n_601),
.Y(n_730)
);

AOI222xp33_ASAP7_75t_L g731 ( 
.A1(n_695),
.A2(n_545),
.B1(n_286),
.B2(n_623),
.C1(n_349),
.C2(n_353),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_669),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_648),
.B(n_603),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_674),
.B(n_611),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_594),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_626),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_683),
.A2(n_545),
.B1(n_618),
.B2(n_615),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_699),
.A2(n_545),
.B1(n_607),
.B2(n_345),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_702),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_632),
.A2(n_605),
.B(n_614),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_706),
.A2(n_605),
.B(n_614),
.Y(n_741)
);

NOR3xp33_ASAP7_75t_L g742 ( 
.A(n_704),
.B(n_451),
.C(n_454),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_647),
.A2(n_586),
.B1(n_616),
.B2(n_610),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_SL g744 ( 
.A1(n_686),
.A2(n_234),
.B1(n_236),
.B2(n_244),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_721),
.A2(n_609),
.B(n_621),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_721),
.A2(n_621),
.B(n_616),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_660),
.B(n_416),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_696),
.B(n_454),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_700),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_672),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_643),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_671),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_656),
.B(n_607),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_642),
.A2(n_630),
.B(n_265),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_694),
.A2(n_440),
.B(n_430),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_633),
.A2(n_440),
.B(n_430),
.C(n_428),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_642),
.A2(n_259),
.B(n_247),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_643),
.B(n_607),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_SL g760 ( 
.A1(n_641),
.A2(n_428),
.B(n_448),
.C(n_260),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_643),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_649),
.Y(n_762)
);

NOR2x1_ASAP7_75t_SL g763 ( 
.A(n_631),
.B(n_447),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_712),
.A2(n_256),
.B(n_250),
.C(n_268),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_653),
.Y(n_765)
);

NOR2x1_ASAP7_75t_L g766 ( 
.A(n_638),
.B(n_448),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_636),
.A2(n_266),
.B(n_257),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_667),
.B(n_246),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_649),
.B(n_448),
.Y(n_769)
);

O2A1O1Ixp5_ASAP7_75t_L g770 ( 
.A1(n_668),
.A2(n_283),
.B(n_255),
.C(n_254),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_681),
.B(n_720),
.C(n_659),
.Y(n_771)
);

AO32x1_ASAP7_75t_L g772 ( 
.A1(n_717),
.A2(n_283),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_772)
);

BUFx8_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_671),
.B(n_283),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_689),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_645),
.B(n_6),
.C(n_10),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_639),
.A2(n_77),
.B(n_173),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_683),
.B(n_6),
.Y(n_778)
);

OA22x2_ASAP7_75t_L g779 ( 
.A1(n_713),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_649),
.B(n_55),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_685),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_702),
.B(n_58),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_702),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_691),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_R g785 ( 
.A(n_685),
.B(n_59),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_644),
.A2(n_11),
.B(n_13),
.Y(n_786)
);

BUFx8_ASAP7_75t_L g787 ( 
.A(n_685),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_640),
.A2(n_92),
.B(n_170),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_726),
.A2(n_634),
.B1(n_635),
.B2(n_637),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_657),
.A2(n_89),
.B(n_168),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_692),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_725),
.B(n_15),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_701),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_725),
.B(n_16),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_677),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_734),
.A2(n_680),
.B(n_661),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_752),
.B(n_673),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_748),
.B(n_652),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_755),
.A2(n_730),
.B(n_740),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_751),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_736),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_733),
.B(n_679),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_771),
.A2(n_662),
.B(n_680),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_735),
.B(n_707),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_746),
.A2(n_665),
.B(n_661),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_735),
.B(n_708),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_768),
.B(n_658),
.Y(n_808)
);

OAI22x1_ASAP7_75t_L g809 ( 
.A1(n_771),
.A2(n_711),
.B1(n_709),
.B2(n_697),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_789),
.A2(n_726),
.B(n_687),
.Y(n_810)
);

AO31x2_ASAP7_75t_L g811 ( 
.A1(n_743),
.A2(n_678),
.A3(n_717),
.B(n_705),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_741),
.A2(n_651),
.B(n_745),
.Y(n_812)
);

OAI22xp33_ASAP7_75t_L g813 ( 
.A1(n_776),
.A2(n_724),
.B1(n_684),
.B2(n_726),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_777),
.A2(n_651),
.B(n_723),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_750),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_732),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_754),
.A2(n_687),
.B(n_703),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_792),
.B(n_714),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_788),
.A2(n_655),
.B(n_715),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_795),
.B(n_714),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_SL g821 ( 
.A1(n_776),
.A2(n_786),
.B(n_760),
.C(n_780),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_786),
.A2(n_724),
.B(n_646),
.C(n_662),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_770),
.A2(n_727),
.B(n_654),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_790),
.A2(n_716),
.B(n_698),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_758),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_737),
.B(n_637),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_742),
.B(n_703),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_787),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_767),
.A2(n_729),
.B(n_676),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_794),
.B(n_719),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_796),
.B(n_666),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_764),
.A2(n_682),
.B(n_675),
.C(n_729),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_773),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_749),
.B(n_722),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_747),
.A2(n_710),
.B(n_670),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_781),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_774),
.B(n_664),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_783),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_762),
.B(n_631),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_757),
.A2(n_690),
.B(n_728),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_787),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_783),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_766),
.A2(n_663),
.B(n_710),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_SL g844 ( 
.A1(n_778),
.A2(n_663),
.B(n_17),
.C(n_18),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_775),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_762),
.A2(n_670),
.B1(n_17),
.B2(n_18),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_731),
.B(n_16),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_784),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_848)
);

AOI221x1_ASAP7_75t_L g849 ( 
.A1(n_738),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_849)
);

AO31x2_ASAP7_75t_L g850 ( 
.A1(n_763),
.A2(n_25),
.A3(n_26),
.B(n_27),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_791),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_731),
.B(n_793),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_847),
.A2(n_738),
.B1(n_773),
.B2(n_744),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_839),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_807),
.A2(n_744),
.B1(n_753),
.B2(n_759),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_807),
.A2(n_802),
.B1(n_837),
.B2(n_809),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_SL g857 ( 
.A1(n_802),
.A2(n_779),
.B1(n_785),
.B2(n_782),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_802),
.A2(n_769),
.B1(n_765),
.B2(n_761),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_838),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_838),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_836),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_852),
.A2(n_769),
.B1(n_761),
.B2(n_751),
.Y(n_862)
);

INVx6_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

INVx6_ASAP7_75t_SL g864 ( 
.A(n_839),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_834),
.Y(n_865)
);

CKINVDCx6p67_ASAP7_75t_R g866 ( 
.A(n_841),
.Y(n_866)
);

BUFx4f_ASAP7_75t_SL g867 ( 
.A(n_841),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_816),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_842),
.Y(n_869)
);

CKINVDCx6p67_ASAP7_75t_R g870 ( 
.A(n_828),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_825),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_805),
.A2(n_849),
.B1(n_808),
.B2(n_799),
.Y(n_872)
);

INVx6_ASAP7_75t_L g873 ( 
.A(n_830),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_827),
.A2(n_756),
.B(n_769),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_828),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_842),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_803),
.A2(n_762),
.B1(n_739),
.B2(n_761),
.Y(n_877)
);

INVx6_ASAP7_75t_L g878 ( 
.A(n_798),
.Y(n_878)
);

CKINVDCx6p67_ASAP7_75t_R g879 ( 
.A(n_815),
.Y(n_879)
);

CKINVDCx6p67_ASAP7_75t_R g880 ( 
.A(n_815),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_845),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_831),
.B(n_739),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_831),
.A2(n_751),
.B1(n_772),
.B2(n_31),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_818),
.B(n_28),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_801),
.Y(n_885)
);

INVx6_ASAP7_75t_L g886 ( 
.A(n_813),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_826),
.A2(n_833),
.B1(n_846),
.B2(n_820),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_844),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_844),
.Y(n_889)
);

CKINVDCx14_ASAP7_75t_R g890 ( 
.A(n_821),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_804),
.A2(n_772),
.B1(n_33),
.B2(n_34),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_850),
.Y(n_892)
);

CKINVDCx14_ASAP7_75t_R g893 ( 
.A(n_821),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_850),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_812),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_806),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_813),
.A2(n_772),
.B1(n_33),
.B2(n_34),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_843),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_797),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_810),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_850),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_840),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_850),
.Y(n_903)
);

INVx5_ASAP7_75t_L g904 ( 
.A(n_832),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_822),
.B(n_37),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_823),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_SL g907 ( 
.A1(n_848),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_907)
);

BUFx12f_ASAP7_75t_L g908 ( 
.A(n_848),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_851),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_800),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_851),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_896),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_894),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_886),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_892),
.B(n_811),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_898),
.B(n_811),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_872),
.B(n_822),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_898),
.Y(n_919)
);

INVx6_ASAP7_75t_L g920 ( 
.A(n_854),
.Y(n_920)
);

AO31x2_ASAP7_75t_L g921 ( 
.A1(n_903),
.A2(n_817),
.A3(n_835),
.B(n_811),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_874),
.A2(n_832),
.B(n_814),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_910),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_910),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_868),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_868),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_871),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_895),
.B(n_811),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_871),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_881),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_889),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_881),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_909),
.B(n_829),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_886),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_911),
.A2(n_819),
.B(n_824),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_886),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_905),
.A2(n_824),
.B(n_115),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_886),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_890),
.B(n_42),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_904),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_890),
.B(n_43),
.Y(n_941)
);

INVx4_ASAP7_75t_SL g942 ( 
.A(n_888),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_904),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_904),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_908),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_904),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_904),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_893),
.Y(n_948)
);

AND3x1_ASAP7_75t_L g949 ( 
.A(n_939),
.B(n_855),
.C(n_856),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_916),
.B(n_893),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_923),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_912),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_918),
.B(n_907),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_916),
.B(n_883),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_918),
.A2(n_908),
.B1(n_853),
.B2(n_902),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_923),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_912),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_916),
.B(n_878),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_916),
.B(n_878),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_935),
.A2(n_897),
.B(n_862),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_922),
.B(n_888),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_916),
.B(n_878),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_945),
.A2(n_906),
.B(n_857),
.C(n_900),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_914),
.B(n_891),
.Y(n_964)
);

AOI221xp5_ASAP7_75t_L g965 ( 
.A1(n_939),
.A2(n_899),
.B1(n_887),
.B2(n_884),
.C(n_865),
.Y(n_965)
);

AOI221xp5_ASAP7_75t_L g966 ( 
.A1(n_941),
.A2(n_900),
.B1(n_882),
.B2(n_877),
.C(n_861),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_920),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_923),
.Y(n_968)
);

INVx6_ASAP7_75t_L g969 ( 
.A(n_914),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_932),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_932),
.B(n_878),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_928),
.B(n_873),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_923),
.B(n_854),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_931),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_922),
.A2(n_885),
.B(n_869),
.C(n_873),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_917),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_941),
.A2(n_858),
.B(n_861),
.C(n_860),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_917),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_923),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_923),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_912),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_913),
.B(n_885),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_945),
.Y(n_984)
);

NAND4xp25_ASAP7_75t_SL g985 ( 
.A(n_948),
.B(n_879),
.C(n_880),
.D(n_866),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_915),
.B(n_873),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_915),
.B(n_873),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_945),
.A2(n_866),
.B1(n_875),
.B2(n_879),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_912),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_971),
.B(n_913),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_976),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_956),
.B(n_923),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_976),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_915),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_971),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_952),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_970),
.B(n_981),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_880),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_970),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_986),
.B(n_928),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_986),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_981),
.B(n_921),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_987),
.B(n_972),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_978),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_978),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_952),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_974),
.Y(n_1007)
);

NAND4xp25_ASAP7_75t_L g1008 ( 
.A(n_965),
.B(n_948),
.C(n_934),
.D(n_936),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_974),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_987),
.B(n_928),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_987),
.B(n_923),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_951),
.B(n_921),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_952),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_957),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_957),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_972),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1003),
.B(n_951),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_993),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_993),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_995),
.B(n_957),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_990),
.B(n_951),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1006),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1007),
.B(n_982),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1003),
.B(n_951),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1006),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_990),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1009),
.B(n_982),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_SL g1028 ( 
.A1(n_1008),
.A2(n_955),
.B1(n_965),
.B2(n_949),
.C(n_963),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_999),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1011),
.B(n_979),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1011),
.B(n_979),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_998),
.A2(n_953),
.B1(n_964),
.B2(n_961),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1013),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1013),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1014),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_992),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_996),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_996),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1014),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.Y(n_1040)
);

AND2x4_ASAP7_75t_SL g1041 ( 
.A(n_1032),
.B(n_950),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1036),
.B(n_992),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1029),
.B(n_1016),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1036),
.B(n_992),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1026),
.B(n_1001),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1026),
.B(n_997),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1017),
.B(n_994),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1037),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1018),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1051),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_1017),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_1040),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1047),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1047),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_1043),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1050),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1050),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_1053),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1056),
.B(n_1046),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1057),
.B(n_1049),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_1049),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1055),
.A2(n_1041),
.B1(n_949),
.B2(n_985),
.Y(n_1064)
);

AOI321xp33_ASAP7_75t_L g1065 ( 
.A1(n_1064),
.A2(n_1028),
.A3(n_955),
.B1(n_1054),
.B2(n_966),
.C(n_977),
.Y(n_1065)
);

NAND4xp25_ASAP7_75t_L g1066 ( 
.A(n_1060),
.B(n_1028),
.C(n_988),
.D(n_1054),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1061),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1062),
.B(n_1054),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_SL g1069 ( 
.A1(n_1063),
.A2(n_1052),
.B(n_977),
.C(n_1059),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1064),
.B(n_1041),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1060),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1060),
.B(n_1052),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1060),
.B(n_1053),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_1045),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1061),
.Y(n_1075)
);

OR3x2_ASAP7_75t_L g1076 ( 
.A(n_1061),
.B(n_867),
.C(n_985),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1071),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1067),
.B(n_875),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1073),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1075),
.A2(n_1072),
.B(n_1068),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1073),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1074),
.B(n_1042),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1066),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_1070),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1076),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_SL g1086 ( 
.A1(n_1069),
.A2(n_1058),
.B(n_1048),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1065),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_1071),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1072),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1073),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1076),
.A2(n_961),
.B1(n_1044),
.B2(n_1042),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_1071),
.Y(n_1092)
);

NOR3x1_ASAP7_75t_L g1093 ( 
.A(n_1084),
.B(n_870),
.C(n_1021),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1087),
.B(n_1045),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1083),
.A2(n_961),
.B1(n_1044),
.B2(n_966),
.Y(n_1095)
);

AOI222xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1088),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.C1(n_46),
.C2(n_50),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1081),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1077),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1079),
.Y(n_1099)
);

NAND4xp25_ASAP7_75t_SL g1100 ( 
.A(n_1086),
.B(n_870),
.C(n_1048),
.D(n_954),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1077),
.Y(n_1101)
);

AO22x2_ASAP7_75t_L g1102 ( 
.A1(n_1090),
.A2(n_942),
.B1(n_1018),
.B2(n_1019),
.Y(n_1102)
);

XOR2x2_ASAP7_75t_L g1103 ( 
.A(n_1078),
.B(n_50),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1081),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1082),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1088),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1082),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1092),
.A2(n_1020),
.B(n_1023),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1092),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1089),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1085),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_1106),
.A2(n_1109),
.B(n_1099),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1098),
.Y(n_1113)
);

NAND4xp25_ASAP7_75t_L g1114 ( 
.A(n_1094),
.B(n_1080),
.C(n_1091),
.D(n_975),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1099),
.B(n_1020),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1101),
.B(n_967),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1097),
.B(n_1104),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1105),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_1110),
.B(n_876),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1107),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_1102),
.B(n_1019),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1103),
.B(n_51),
.Y(n_1122)
);

AND3x4_ASAP7_75t_L g1123 ( 
.A(n_1111),
.B(n_956),
.C(n_968),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1094),
.B(n_1021),
.Y(n_1124)
);

XNOR2xp5_ASAP7_75t_L g1125 ( 
.A(n_1095),
.B(n_1102),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_1108),
.A2(n_1023),
.B(n_1027),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1093),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1100),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1117),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1122),
.B(n_1096),
.Y(n_1130)
);

NOR4xp25_ASAP7_75t_L g1131 ( 
.A(n_1112),
.B(n_1100),
.C(n_1096),
.D(n_1027),
.Y(n_1131)
);

AOI222xp33_ASAP7_75t_L g1132 ( 
.A1(n_1112),
.A2(n_1113),
.B1(n_1125),
.B2(n_1115),
.C1(n_1118),
.C2(n_1120),
.Y(n_1132)
);

OAI211xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1127),
.A2(n_975),
.B(n_1033),
.C(n_1025),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1128),
.A2(n_954),
.B(n_936),
.Y(n_1134)
);

AOI211xp5_ASAP7_75t_L g1135 ( 
.A1(n_1114),
.A2(n_937),
.B(n_980),
.C(n_854),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1124),
.B(n_1024),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1121),
.Y(n_1137)
);

OAI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1116),
.A2(n_961),
.B1(n_1034),
.B2(n_1039),
.C(n_1035),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1126),
.A2(n_937),
.B(n_964),
.C(n_960),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1123),
.B(n_876),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1119),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1118),
.B(n_1024),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1122),
.B(n_1022),
.Y(n_1143)
);

OAI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1112),
.A2(n_961),
.B1(n_956),
.B2(n_968),
.C(n_1012),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1112),
.A2(n_937),
.B(n_964),
.C(n_960),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1122),
.A2(n_60),
.B(n_61),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1112),
.A2(n_961),
.B(n_933),
.Y(n_1147)
);

AOI321xp33_ASAP7_75t_L g1148 ( 
.A1(n_1112),
.A2(n_954),
.A3(n_973),
.B1(n_950),
.B2(n_938),
.C(n_934),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1112),
.A2(n_933),
.B(n_1038),
.Y(n_1149)
);

OAI211xp5_ASAP7_75t_L g1150 ( 
.A1(n_1112),
.A2(n_885),
.B(n_869),
.C(n_979),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1122),
.A2(n_960),
.B(n_859),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1128),
.A2(n_942),
.B1(n_980),
.B2(n_973),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1131),
.A2(n_1039),
.B1(n_1022),
.B2(n_1025),
.C(n_1035),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1132),
.B(n_1033),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1130),
.B(n_979),
.C(n_869),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1142),
.A2(n_942),
.B1(n_980),
.B2(n_973),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1129),
.A2(n_1034),
.B1(n_1038),
.B2(n_1037),
.C(n_1005),
.Y(n_1157)
);

AOI221x1_ASAP7_75t_L g1158 ( 
.A1(n_1146),
.A2(n_1038),
.B1(n_1037),
.B2(n_1004),
.C(n_991),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1152),
.A2(n_859),
.B(n_860),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1137),
.Y(n_1160)
);

AOI211xp5_ASAP7_75t_L g1161 ( 
.A1(n_1141),
.A2(n_980),
.B(n_854),
.C(n_938),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1143),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1134),
.A2(n_942),
.B1(n_980),
.B2(n_973),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1144),
.A2(n_1136),
.B1(n_1138),
.B2(n_1135),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1140),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1147),
.A2(n_980),
.B1(n_1015),
.B2(n_968),
.C(n_919),
.Y(n_1166)
);

AOI32xp33_ASAP7_75t_L g1167 ( 
.A1(n_1133),
.A2(n_950),
.A3(n_994),
.B1(n_914),
.B2(n_958),
.Y(n_1167)
);

AOI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1150),
.A2(n_980),
.B(n_854),
.C(n_1012),
.Y(n_1168)
);

AOI222xp33_ASAP7_75t_L g1169 ( 
.A1(n_1145),
.A2(n_942),
.B1(n_914),
.B2(n_931),
.C1(n_1015),
.C2(n_925),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1151),
.A2(n_942),
.B1(n_863),
.B2(n_920),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1151),
.A2(n_1149),
.B1(n_1139),
.B2(n_1148),
.C(n_919),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1132),
.B(n_997),
.Y(n_1172)
);

AOI211xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1130),
.A2(n_983),
.B(n_1002),
.C(n_943),
.Y(n_1173)
);

NOR4xp25_ASAP7_75t_L g1174 ( 
.A(n_1130),
.B(n_983),
.C(n_927),
.D(n_925),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1131),
.A2(n_919),
.B1(n_927),
.B2(n_926),
.C(n_929),
.Y(n_1175)
);

NAND4xp25_ASAP7_75t_L g1176 ( 
.A(n_1132),
.B(n_914),
.C(n_959),
.D(n_962),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_942),
.B1(n_863),
.B2(n_920),
.Y(n_1177)
);

OAI211xp5_ASAP7_75t_L g1178 ( 
.A1(n_1160),
.A2(n_1002),
.B(n_943),
.C(n_929),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1165),
.Y(n_1179)
);

XOR2x2_ASAP7_75t_L g1180 ( 
.A(n_1172),
.B(n_63),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1162),
.B(n_1154),
.C(n_1164),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_L g1182 ( 
.A(n_1159),
.B(n_68),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1155),
.B(n_924),
.C(n_926),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1158),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1171),
.A2(n_863),
.B1(n_920),
.B2(n_969),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_L g1186 ( 
.A(n_1175),
.B(n_70),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1174),
.B(n_71),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1156),
.A2(n_863),
.B1(n_920),
.B2(n_969),
.Y(n_1188)
);

XNOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1170),
.B(n_73),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1163),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1167),
.B(n_959),
.Y(n_1191)
);

NOR2x1_ASAP7_75t_L g1192 ( 
.A(n_1173),
.B(n_74),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1161),
.B(n_1010),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1153),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1166),
.B(n_920),
.Y(n_1195)
);

NAND4xp75_ASAP7_75t_L g1196 ( 
.A(n_1157),
.B(n_944),
.C(n_924),
.D(n_1000),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1168),
.B(n_1010),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1169),
.B(n_1000),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1179),
.B(n_962),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_L g1200 ( 
.A(n_1181),
.B(n_935),
.C(n_924),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1180),
.A2(n_1177),
.B1(n_1185),
.B2(n_1195),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1194),
.A2(n_962),
.B(n_958),
.Y(n_1202)
);

OR3x2_ASAP7_75t_L g1203 ( 
.A(n_1184),
.B(n_864),
.C(n_93),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_L g1204 ( 
.A(n_1190),
.B(n_935),
.C(n_958),
.Y(n_1204)
);

OAI211xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1186),
.A2(n_84),
.B(n_94),
.C(n_99),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1197),
.B(n_930),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1192),
.B(n_969),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1182),
.B(n_969),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1187),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1191),
.B(n_930),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1189),
.B(n_930),
.C(n_947),
.Y(n_1211)
);

AND4x1_ASAP7_75t_L g1212 ( 
.A(n_1188),
.B(n_864),
.C(n_101),
.D(n_102),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1193),
.B(n_969),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1209),
.B(n_1191),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1199),
.Y(n_1215)
);

OAI211xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1201),
.A2(n_1183),
.B(n_1178),
.C(n_1198),
.Y(n_1216)
);

INVxp33_ASAP7_75t_SL g1217 ( 
.A(n_1207),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1203),
.A2(n_1196),
.B1(n_864),
.B2(n_944),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1199),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1208),
.B(n_944),
.Y(n_1220)
);

BUFx2_ASAP7_75t_SL g1221 ( 
.A(n_1212),
.Y(n_1221)
);

NOR4xp25_ASAP7_75t_L g1222 ( 
.A(n_1205),
.B(n_100),
.C(n_106),
.D(n_107),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1206),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1202),
.A2(n_947),
.B1(n_946),
.B2(n_940),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1213),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1200),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1211),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1204),
.B(n_947),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1215),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1217),
.A2(n_1210),
.B1(n_947),
.B2(n_946),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1221),
.A2(n_1216),
.B1(n_1214),
.B2(n_1219),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1225),
.A2(n_946),
.B1(n_940),
.B2(n_989),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1225),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1218),
.A2(n_1227),
.B1(n_1223),
.B2(n_1226),
.Y(n_1234)
);

OR3x2_ASAP7_75t_L g1235 ( 
.A(n_1222),
.B(n_111),
.C(n_112),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1220),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1224),
.Y(n_1237)
);

OAI22x1_ASAP7_75t_L g1238 ( 
.A1(n_1228),
.A2(n_946),
.B1(n_940),
.B2(n_989),
.Y(n_1238)
);

AOI311xp33_ASAP7_75t_L g1239 ( 
.A1(n_1233),
.A2(n_113),
.A3(n_117),
.B(n_118),
.C(n_121),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1229),
.A2(n_940),
.B(n_125),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1231),
.B(n_123),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_SL g1242 ( 
.A(n_1236),
.B(n_127),
.Y(n_1242)
);

INVxp33_ASAP7_75t_L g1243 ( 
.A(n_1234),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_1237),
.A2(n_989),
.B1(n_982),
.B2(n_132),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1241),
.B(n_1230),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1240),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1243),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1242),
.A2(n_1238),
.B(n_1235),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1246),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1249),
.A2(n_1247),
.B(n_1245),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1250),
.A2(n_1248),
.B(n_1232),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1251),
.Y(n_1252)
);

OAI221xp5_ASAP7_75t_R g1253 ( 
.A1(n_1252),
.A2(n_1239),
.B1(n_1244),
.B2(n_133),
.C(n_135),
.Y(n_1253)
);

AOI211xp5_ASAP7_75t_L g1254 ( 
.A1(n_1253),
.A2(n_128),
.B(n_130),
.C(n_138),
.Y(n_1254)
);


endmodule