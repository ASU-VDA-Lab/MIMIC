module fake_jpeg_3098_n_541 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_52),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_53),
.B(n_60),
.Y(n_148)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_14),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_32),
.B(n_13),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_28),
.Y(n_102)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_13),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_11),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_11),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_149),
.C(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_29),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_104),
.B(n_90),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_34),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_83),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_34),
.B1(n_44),
.B2(n_25),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_116),
.A2(n_129),
.B1(n_131),
.B2(n_147),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_27),
.B1(n_33),
.B2(n_25),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_44),
.B1(n_35),
.B2(n_29),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_51),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_151),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_34),
.B1(n_44),
.B2(n_35),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_156),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_52),
.B(n_31),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_163),
.A2(n_183),
.B1(n_200),
.B2(n_208),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_48),
.C(n_55),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_168),
.B(n_195),
.C(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_169),
.B(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_186),
.B1(n_206),
.B2(n_105),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_99),
.A2(n_81),
.B1(n_83),
.B2(n_34),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_36),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_41),
.B1(n_36),
.B2(n_34),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_218)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_116),
.A2(n_86),
.B1(n_77),
.B2(n_76),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_68),
.B1(n_65),
.B2(n_95),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_108),
.A2(n_31),
.B1(n_37),
.B2(n_41),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_189),
.A2(n_20),
.B1(n_150),
.B2(n_158),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_108),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_194),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_37),
.B1(n_41),
.B2(n_98),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_157),
.B1(n_132),
.B2(n_90),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_24),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_24),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_157),
.A2(n_24),
.B1(n_38),
.B2(n_89),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_117),
.B(n_38),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_132),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_96),
.B1(n_38),
.B2(n_15),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_209),
.A2(n_210),
.B1(n_160),
.B2(n_137),
.Y(n_240)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_105),
.B1(n_155),
.B2(n_152),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_123),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_234),
.C(n_238),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_119),
.A3(n_132),
.B1(n_124),
.B2(n_136),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_178),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_226),
.B1(n_186),
.B2(n_206),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_120),
.B1(n_122),
.B2(n_141),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_173),
.A2(n_120),
.B1(n_122),
.B2(n_141),
.Y(n_236)
);

AO21x2_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_244),
.B(n_210),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_168),
.B(n_127),
.CI(n_93),
.CON(n_242),
.SN(n_242)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_242),
.A2(n_164),
.B(n_191),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_158),
.B1(n_127),
.B2(n_160),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_201),
.B1(n_175),
.B2(n_165),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_195),
.C(n_172),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_256),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_257),
.B1(n_262),
.B2(n_267),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_195),
.B(n_172),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_251),
.A2(n_254),
.B(n_272),
.Y(n_303)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_183),
.B1(n_205),
.B2(n_178),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_170),
.C(n_176),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_258),
.B(n_270),
.Y(n_287)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_190),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_263),
.Y(n_294)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_171),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_162),
.B1(n_196),
.B2(n_187),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_225),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_233),
.Y(n_290)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_165),
.B1(n_167),
.B2(n_175),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_221),
.B(n_218),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_227),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_280),
.Y(n_306)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_236),
.B1(n_244),
.B2(n_229),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_285),
.A2(n_289),
.B1(n_291),
.B2(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_260),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_288),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_229),
.B1(n_242),
.B2(n_223),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_242),
.B1(n_214),
.B2(n_248),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_299),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_293),
.B(n_177),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_233),
.B1(n_226),
.B2(n_219),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_298),
.A2(n_304),
.B(n_231),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_276),
.B(n_252),
.Y(n_304)
);

OAI211xp5_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_221),
.B(n_218),
.C(n_235),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_262),
.A2(n_240),
.B1(n_235),
.B2(n_241),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_299),
.B1(n_278),
.B2(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_277),
.B(n_241),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_294),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_318),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_262),
.B1(n_278),
.B2(n_252),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_325),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_319),
.B(n_336),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_294),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_256),
.B1(n_270),
.B2(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_249),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_340),
.C(n_341),
.Y(n_355)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

OAI22x1_ASAP7_75t_SL g325 ( 
.A1(n_289),
.A2(n_264),
.B1(n_274),
.B2(n_273),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_251),
.B1(n_271),
.B2(n_269),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_311),
.B1(n_310),
.B2(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_342),
.B(n_303),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_332),
.B(n_182),
.Y(n_376)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_258),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_SL g373 ( 
.A(n_335),
.B(n_243),
.Y(n_373)
);

OAI211xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_280),
.B(n_217),
.C(n_268),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_261),
.B1(n_259),
.B2(n_253),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_338),
.A2(n_297),
.B1(n_310),
.B2(n_311),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_306),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_339),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_185),
.C(n_188),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_204),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_309),
.A2(n_202),
.B(n_197),
.C(n_121),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_331),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_363),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_287),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_356),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_353),
.A2(n_360),
.B1(n_374),
.B2(n_325),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_357),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_295),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_315),
.A2(n_303),
.B(n_308),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_306),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_370),
.C(n_326),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_327),
.A2(n_288),
.B1(n_292),
.B2(n_291),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_327),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_367),
.A2(n_368),
.B1(n_338),
.B2(n_316),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_315),
.A2(n_296),
.B1(n_302),
.B2(n_284),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_296),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_318),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_330),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_377),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_317),
.A2(n_284),
.B1(n_283),
.B2(n_302),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_329),
.A2(n_302),
.B(n_283),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_342),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_376),
.B(n_228),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_243),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_374),
.B1(n_367),
.B2(n_357),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_382),
.B(n_350),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_383),
.A2(n_385),
.B1(n_400),
.B2(n_408),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_320),
.C(n_313),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_387),
.C(n_396),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_346),
.A2(n_314),
.B1(n_333),
.B2(n_343),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_370),
.C(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_366),
.A2(n_314),
.B(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_397),
.Y(n_411)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_351),
.A2(n_345),
.B1(n_322),
.B2(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_355),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_334),
.Y(n_394)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_328),
.C(n_324),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_239),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_401),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_239),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_342),
.B1(n_246),
.B2(n_203),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_247),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_368),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_405),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_348),
.A2(n_342),
.B1(n_246),
.B2(n_216),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_407),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_247),
.C(n_246),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_353),
.A2(n_342),
.B1(n_203),
.B2(n_216),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_348),
.B(n_228),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_364),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_410),
.A2(n_416),
.B1(n_389),
.B2(n_402),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_419),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_354),
.B1(n_375),
.B2(n_362),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_347),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_418),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_382),
.Y(n_418)
);

AOI21xp33_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_362),
.B(n_361),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_395),
.A2(n_347),
.B(n_361),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_424),
.A2(n_390),
.B(n_383),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_427),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_350),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_349),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_437),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_433),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_386),
.B(n_349),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_436),
.B(n_431),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_232),
.Y(n_437)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_434),
.A2(n_389),
.B1(n_400),
.B2(n_408),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_440),
.A2(n_410),
.B1(n_416),
.B2(n_422),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_407),
.C(n_399),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_453),
.C(n_456),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_442),
.A2(n_455),
.B1(n_459),
.B2(n_10),
.Y(n_481)
);

AOI211xp5_ASAP7_75t_L g444 ( 
.A1(n_420),
.A2(n_211),
.B(n_192),
.C(n_220),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_444),
.A2(n_134),
.B1(n_40),
.B2(n_20),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_232),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_447),
.B(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_436),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_184),
.C(n_166),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_207),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_192),
.C(n_152),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_164),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_460),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_220),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_421),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_415),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_220),
.C(n_140),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_412),
.C(n_437),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_462),
.A2(n_477),
.B1(n_444),
.B2(n_449),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_470),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_479),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_430),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_476),
.B(n_20),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_412),
.C(n_413),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_474),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_471),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_428),
.C(n_435),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_140),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_478),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_442),
.A2(n_134),
.B(n_40),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_15),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_15),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_440),
.A2(n_15),
.B1(n_10),
.B2(n_2),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_480),
.B(n_476),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_452),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_468),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_483),
.B(n_492),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_497),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_495),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_464),
.Y(n_487)
);

OAI21x1_ASAP7_75t_SL g514 ( 
.A1(n_487),
.A2(n_489),
.B(n_490),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_458),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_471),
.A2(n_446),
.B(n_439),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_463),
.B(n_456),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_466),
.B(n_461),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_493),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_441),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_453),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_498),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_465),
.A2(n_15),
.B(n_20),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_478),
.B(n_479),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_469),
.B(n_467),
.C(n_466),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_500),
.A2(n_505),
.B(n_509),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_490),
.B(n_485),
.CI(n_487),
.CON(n_502),
.SN(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_506),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_4),
.Y(n_519)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_0),
.B(n_1),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_15),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_0),
.B(n_1),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_497),
.B(n_484),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_510),
.A2(n_511),
.B(n_3),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_494),
.A2(n_499),
.B(n_488),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_SL g512 ( 
.A1(n_494),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_2),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g516 ( 
.A(n_501),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_519),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_517),
.A2(n_508),
.B1(n_512),
.B2(n_507),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_9),
.C(n_6),
.Y(n_520)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_520),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_501),
.A2(n_5),
.B(n_6),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_521),
.A2(n_522),
.B(n_524),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_503),
.A2(n_5),
.B(n_6),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_5),
.C(n_6),
.Y(n_523)
);

MAJx2_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_525),
.C(n_7),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_508),
.B(n_7),
.Y(n_525)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_527),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_530),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_500),
.C(n_8),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_531),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_520),
.B(n_8),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_535),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_534),
.C(n_526),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_528),
.C(n_536),
.Y(n_539)
);

AOI21x1_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_538),
.B(n_7),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_9),
.C(n_227),
.Y(n_541)
);


endmodule