module fake_jpeg_13921_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_53),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_15),
.A2(n_7),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_15),
.B(n_6),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_68),
.Y(n_113)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_92),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_34),
.B1(n_28),
.B2(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_81),
.B(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_28),
.B1(n_29),
.B2(n_21),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_18),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_85),
.A2(n_106),
.B1(n_96),
.B2(n_94),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_28),
.B1(n_29),
.B2(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_89),
.A2(n_104),
.B1(n_0),
.B2(n_1),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_27),
.B1(n_22),
.B2(n_36),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_30),
.B1(n_27),
.B2(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_35),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_44),
.A2(n_18),
.B1(n_33),
.B2(n_36),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_16),
.B1(n_36),
.B2(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_0),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_18),
.B1(n_33),
.B2(n_20),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_33),
.B1(n_20),
.B2(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_105),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_25),
.B1(n_27),
.B2(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_30),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_1),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_70),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_122),
.B(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_31),
.B1(n_8),
.B2(n_9),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_88),
.B1(n_89),
.B2(n_81),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_0),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_137),
.B(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_114),
.B1(n_87),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_84),
.B1(n_109),
.B2(n_108),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_147),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_6),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_145),
.B1(n_102),
.B2(n_82),
.Y(n_168)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_149),
.Y(n_161)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_73),
.A2(n_8),
.B(n_12),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_85),
.B1(n_96),
.B2(n_79),
.Y(n_170)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_76),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_155),
.B(n_78),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_14),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_86),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_160),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_85),
.B1(n_93),
.B2(n_97),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_171),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_82),
.B1(n_102),
.B2(n_111),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_166),
.A2(n_196),
.B1(n_143),
.B2(n_154),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_100),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_191),
.B1(n_193),
.B2(n_195),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_129),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_144),
.C(n_137),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_179),
.C(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_188),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_122),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_142),
.A2(n_96),
.B1(n_111),
.B2(n_74),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_117),
.B(n_116),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_112),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_127),
.A2(n_112),
.B1(n_77),
.B2(n_95),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_118),
.A2(n_77),
.B1(n_95),
.B2(n_108),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_119),
.A2(n_109),
.B1(n_84),
.B2(n_107),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_121),
.A2(n_74),
.B1(n_107),
.B2(n_9),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_107),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_133),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_199),
.B(n_200),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_119),
.B(n_151),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_204),
.A2(n_213),
.B(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_172),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_213),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_207),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_133),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_218),
.C(n_174),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_135),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_215),
.B(n_226),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_164),
.A2(n_153),
.B1(n_151),
.B2(n_123),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_222),
.B1(n_205),
.B2(n_221),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_170),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_115),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_158),
.A2(n_126),
.B1(n_125),
.B2(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_149),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_223),
.B(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_228),
.Y(n_252)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_162),
.A2(n_146),
.B1(n_132),
.B2(n_139),
.Y(n_228)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_139),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_173),
.B(n_131),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_128),
.B1(n_136),
.B2(n_131),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_186),
.B1(n_181),
.B2(n_169),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_9),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_191),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_190),
.B1(n_175),
.B2(n_169),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_2),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_259),
.C(n_263),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_219),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_206),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_189),
.B1(n_193),
.B2(n_170),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_244),
.A2(n_255),
.B(n_270),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_217),
.B1(n_158),
.B2(n_198),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_211),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_203),
.B(n_226),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_159),
.B1(n_192),
.B2(n_168),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_183),
.C(n_192),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_269),
.B1(n_222),
.B2(n_172),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_202),
.C(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_200),
.B(n_185),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_165),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_272),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_215),
.B(n_185),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_160),
.C(n_161),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_228),
.C(n_227),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_SL g270 ( 
.A1(n_204),
.A2(n_160),
.B(n_175),
.Y(n_270)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_160),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_281),
.C(n_285),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_217),
.B1(n_203),
.B2(n_202),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_301),
.B1(n_259),
.B2(n_239),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_231),
.B(n_237),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_235),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_298),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_284),
.A2(n_292),
.B(n_282),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_216),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_296),
.B1(n_243),
.B2(n_248),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_295),
.Y(n_324)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_233),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_293),
.C(n_240),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_234),
.B(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_252),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_245),
.A2(n_228),
.B1(n_210),
.B2(n_201),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_258),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_244),
.A2(n_212),
.B1(n_209),
.B2(n_190),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_305),
.A2(n_306),
.B1(n_293),
.B2(n_325),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_248),
.B1(n_261),
.B2(n_246),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_321),
.Y(n_347)
);

BUFx4f_ASAP7_75t_SL g309 ( 
.A(n_288),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_317),
.C(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_272),
.B1(n_257),
.B2(n_246),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_257),
.B1(n_246),
.B2(n_266),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_271),
.C(n_247),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_271),
.C(n_247),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_250),
.C(n_242),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_291),
.C(n_274),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_292),
.A2(n_275),
.B(n_284),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_321),
.A2(n_280),
.B(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_258),
.B1(n_242),
.B2(n_250),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_301),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_294),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_333),
.B(n_325),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_296),
.B1(n_275),
.B2(n_287),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_346),
.B1(n_323),
.B2(n_315),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_307),
.B(n_290),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_338),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_285),
.C(n_278),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_343),
.C(n_319),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_279),
.Y(n_338)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_306),
.A2(n_297),
.B(n_279),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_273),
.C(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_326),
.A2(n_286),
.B1(n_277),
.B2(n_289),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_349),
.A2(n_356),
.B(n_342),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

AO221x1_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_334),
.B1(n_304),
.B2(n_320),
.C(n_311),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_335),
.A2(n_316),
.B1(n_303),
.B2(n_312),
.Y(n_353)
);

OAI321xp33_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_354),
.A3(n_363),
.B1(n_362),
.B2(n_344),
.C(n_341),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_303),
.B1(n_312),
.B2(n_318),
.Y(n_354)
);

AOI21xp33_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_308),
.B(n_317),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_331),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_330),
.B(n_305),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_358),
.B(n_360),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_320),
.C(n_304),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_371),
.B(n_353),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_SL g366 ( 
.A1(n_359),
.A2(n_332),
.A3(n_336),
.B1(n_347),
.B2(n_329),
.C1(n_346),
.C2(n_339),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_368),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_328),
.C(n_343),
.Y(n_368)
);

NOR3xp33_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_332),
.C(n_313),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_370),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_337),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_347),
.B(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_340),
.B(n_345),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_374),
.A2(n_362),
.B(n_355),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_357),
.Y(n_386)
);

INVx11_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_365),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_377),
.B(n_375),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_363),
.Y(n_378)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_381),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_350),
.B(n_361),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_384),
.A2(n_387),
.B1(n_309),
.B2(n_249),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_386),
.B(n_368),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_348),
.B(n_352),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_393),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_392),
.Y(n_397)
);

AOI322xp5_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_367),
.A3(n_334),
.B1(n_311),
.B2(n_340),
.C1(n_348),
.C2(n_309),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g393 ( 
.A1(n_380),
.A2(n_340),
.A3(n_309),
.B1(n_338),
.B2(n_254),
.C1(n_229),
.C2(n_249),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_395),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_386),
.B(n_172),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_161),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_3),
.C(n_5),
.Y(n_400)
);

AOI321xp33_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_382),
.A3(n_383),
.B1(n_380),
.B2(n_387),
.C(n_378),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_390),
.A2(n_379),
.B(n_229),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_396),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_390),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_401),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_402),
.C(n_394),
.Y(n_406)
);

AOI321xp33_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_407),
.A3(n_401),
.B1(n_404),
.B2(n_3),
.C(n_5),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_408),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_3),
.Y(n_410)
);


endmodule