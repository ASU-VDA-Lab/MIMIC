module fake_jpeg_28559_n_451 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_9),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_66),
.Y(n_108)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_57),
.Y(n_114)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_92),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_93),
.Y(n_131)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_90),
.Y(n_110)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_22),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_47),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_99),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_17),
.B1(n_39),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_86),
.B1(n_28),
.B2(n_41),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_67),
.B1(n_65),
.B2(n_49),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_136),
.B1(n_28),
.B2(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_70),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_135),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_51),
.B(n_19),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_22),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_46),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_48),
.A2(n_17),
.B1(n_41),
.B2(n_29),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_71),
.A2(n_39),
.B(n_38),
.C(n_35),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_33),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_55),
.B(n_19),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_42),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_29),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_188),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_106),
.B(n_0),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_151),
.B(n_166),
.C(n_177),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_42),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_167),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_102),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_156),
.Y(n_234)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_125),
.B1(n_126),
.B2(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

NAND2x1_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_73),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_58),
.B1(n_100),
.B2(n_105),
.Y(n_212)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_68),
.C(n_78),
.Y(n_166)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_170),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_191),
.B1(n_114),
.B2(n_62),
.Y(n_202)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_98),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_173),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_111),
.A2(n_87),
.B1(n_43),
.B2(n_35),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_96),
.B(n_0),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_192),
.Y(n_208)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_180),
.Y(n_223)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_181),
.Y(n_226)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_182),
.A2(n_187),
.B1(n_195),
.B2(n_196),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_190),
.Y(n_227)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

OR2x6_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_145),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_186),
.A2(n_197),
.B(n_134),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_43),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_109),
.B(n_28),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_97),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_102),
.B(n_33),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_119),
.A2(n_92),
.B1(n_81),
.B2(n_80),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_112),
.B1(n_52),
.B2(n_101),
.Y(n_237)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_114),
.A2(n_31),
.B(n_45),
.C(n_46),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_237),
.B1(n_159),
.B2(n_173),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_201),
.A2(n_202),
.B1(n_230),
.B2(n_212),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_118),
.B1(n_77),
.B2(n_126),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_209),
.B1(n_217),
.B2(n_218),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_154),
.A2(n_145),
.B1(n_129),
.B2(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_150),
.A2(n_105),
.B1(n_61),
.B2(n_53),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_53),
.B1(n_61),
.B2(n_137),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_162),
.A2(n_148),
.B(n_116),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_221),
.A2(n_181),
.B(n_173),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_151),
.B(n_31),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_236),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_148),
.B1(n_116),
.B2(n_100),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_195),
.B1(n_196),
.B2(n_181),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_153),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_151),
.B(n_17),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_176),
.C(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_253),
.C(n_273),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_162),
.B(n_176),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_241),
.A2(n_243),
.B(n_215),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_265),
.B1(n_269),
.B2(n_244),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_176),
.B(n_188),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_251),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_177),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_246),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_177),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_157),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_248),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_166),
.Y(n_248)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_201),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_158),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_206),
.A2(n_197),
.B1(n_170),
.B2(n_178),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_262),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_152),
.B(n_149),
.C(n_165),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_257),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_172),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_261),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_259),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_155),
.B(n_180),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_260),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_182),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_206),
.A2(n_163),
.B1(n_160),
.B2(n_156),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_213),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_200),
.A2(n_179),
.B1(n_164),
.B2(n_169),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_266),
.A2(n_211),
.B(n_207),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_234),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_168),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_271),
.Y(n_294)
);

INVx5_ASAP7_75t_SL g269 ( 
.A(n_201),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_229),
.B1(n_205),
.B2(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_208),
.B(n_185),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_187),
.C(n_23),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_239),
.B(n_212),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_296),
.B(n_304),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_202),
.B1(n_212),
.B2(n_237),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_281),
.B1(n_288),
.B2(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_23),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_252),
.B1(n_239),
.B2(n_257),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_280),
.A2(n_301),
.B1(n_305),
.B2(n_267),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_203),
.B1(n_217),
.B2(n_231),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_283),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_232),
.C(n_218),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_291),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_249),
.A2(n_215),
.B1(n_223),
.B2(n_232),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_226),
.B(n_230),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_293),
.Y(n_325)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_241),
.A2(n_226),
.B(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_247),
.B(n_224),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_258),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_243),
.B(n_271),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_255),
.A2(n_220),
.B(n_224),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_242),
.A2(n_216),
.B1(n_204),
.B2(n_213),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_274),
.A2(n_254),
.B1(n_251),
.B2(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_307),
.A2(n_316),
.B1(n_323),
.B2(n_326),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_253),
.C(n_238),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_318),
.C(n_324),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_281),
.B1(n_298),
.B2(n_274),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_273),
.B1(n_262),
.B2(n_256),
.Y(n_310)
);

AOI22x1_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_307),
.B1(n_276),
.B2(n_314),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_274),
.B(n_290),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_265),
.B1(n_253),
.B2(n_261),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_246),
.C(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_256),
.B1(n_240),
.B2(n_272),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_322),
.A2(n_327),
.B1(n_330),
.B2(n_298),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_274),
.A2(n_263),
.B1(n_259),
.B2(n_250),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_240),
.C(n_207),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_277),
.A2(n_250),
.B1(n_211),
.B2(n_233),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_233),
.B1(n_219),
.B2(n_3),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_219),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_333),
.C(n_334),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_302),
.B1(n_290),
.B2(n_279),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_23),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_294),
.B(n_10),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_335),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_23),
.C(n_1),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_23),
.C(n_1),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_279),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_324),
.B(n_276),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_336),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_291),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_353),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_344),
.B1(n_346),
.B2(n_349),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_350),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_343),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_312),
.A2(n_282),
.B1(n_287),
.B2(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_296),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_293),
.B1(n_300),
.B2(n_304),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_352),
.B1(n_326),
.B2(n_321),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_313),
.A2(n_299),
.B1(n_306),
.B2(n_293),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_284),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_284),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_357),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_298),
.B1(n_293),
.B2(n_302),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_356),
.A2(n_358),
.B1(n_360),
.B2(n_317),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_306),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_282),
.B1(n_289),
.B2(n_295),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_313),
.A2(n_289),
.B1(n_287),
.B2(n_1),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_316),
.C(n_314),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_369),
.C(n_372),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_339),
.C(n_353),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_319),
.Y(n_370)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_310),
.C(n_323),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_352),
.Y(n_373)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_310),
.C(n_333),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_4),
.C(n_8),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_378),
.B1(n_380),
.B2(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_379),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_351),
.B1(n_349),
.B2(n_357),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_320),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_337),
.A2(n_317),
.B1(n_287),
.B2(n_334),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_348),
.B1(n_342),
.B2(n_4),
.Y(n_388)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_382),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_371),
.B(n_342),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_389),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_364),
.B(n_341),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_387),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_388),
.A2(n_396),
.B1(n_361),
.B2(n_380),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_370),
.B(n_348),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_2),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_398),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_379),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_393),
.A2(n_363),
.B1(n_375),
.B2(n_381),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_2),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_397),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_2),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_390),
.Y(n_403)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_400),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_408),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_361),
.B(n_376),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_411),
.Y(n_418)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_378),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_407),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_373),
.B1(n_394),
.B2(n_392),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_368),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_368),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_367),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_399),
.A2(n_372),
.B1(n_374),
.B2(n_364),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_413),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_367),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_413),
.C(n_406),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_409),
.B(n_398),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_419),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_387),
.C(n_393),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_383),
.C(n_384),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_424),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_14),
.C(n_10),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_402),
.A2(n_4),
.B(n_10),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_425),
.A2(n_407),
.B1(n_404),
.B2(n_12),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_401),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_429),
.Y(n_436)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_419),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_403),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_434),
.B(n_418),
.Y(n_435)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_421),
.A2(n_423),
.B(n_418),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_432),
.A2(n_427),
.B(n_428),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_424),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_406),
.C(n_11),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_438),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_440),
.C(n_10),
.Y(n_444)
);

INVx11_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_439),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_439),
.A2(n_431),
.B(n_414),
.Y(n_442)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_442),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_444),
.B(n_436),
.C(n_12),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_446),
.A2(n_441),
.B(n_443),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_447),
.A2(n_445),
.B(n_12),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_11),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_14),
.B(n_343),
.Y(n_451)
);


endmodule