module fake_jpeg_2380_n_448 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_18),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_56),
.B(n_85),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_15),
.C(n_13),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_20),
.A2(n_15),
.B(n_9),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_61),
.B(n_99),
.Y(n_177)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_65),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_66),
.Y(n_147)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_9),
.C(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_73),
.Y(n_125)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_18),
.B(n_8),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_78),
.Y(n_162)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_22),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_0),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_95),
.Y(n_129)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_0),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_29),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_102),
.Y(n_142)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_106),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_36),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_33),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_113),
.Y(n_152)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_22),
.Y(n_141)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_42),
.B(n_3),
.C(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_114),
.Y(n_160)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_4),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_41),
.B1(n_43),
.B2(n_49),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_126),
.A2(n_128),
.B1(n_153),
.B2(n_163),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_84),
.A2(n_41),
.B1(n_43),
.B2(n_49),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_60),
.B(n_51),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_135),
.B(n_144),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_52),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_138),
.B(n_141),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_37),
.B1(n_51),
.B2(n_36),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_140),
.A2(n_156),
.B1(n_116),
.B2(n_147),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_175),
.B1(n_128),
.B2(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_69),
.B(n_38),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_75),
.A2(n_41),
.B1(n_38),
.B2(n_42),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_104),
.B1(n_97),
.B2(n_96),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_86),
.B(n_28),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_161),
.B(n_164),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_26),
.B1(n_34),
.B2(n_52),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_37),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_65),
.B(n_37),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_165),
.B(n_169),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_65),
.B(n_3),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_3),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_178),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_70),
.A2(n_32),
.B1(n_5),
.B2(n_7),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_176),
.B(n_179),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_94),
.B(n_4),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_91),
.B(n_5),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_62),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_77),
.B(n_32),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_74),
.B(n_32),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_80),
.A2(n_90),
.B1(n_83),
.B2(n_89),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_186),
.B1(n_132),
.B2(n_170),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_101),
.B(n_107),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_158),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_84),
.B1(n_72),
.B2(n_21),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

BUFx2_ASAP7_75t_SL g267 ( 
.A(n_190),
.Y(n_267)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_193),
.A2(n_220),
.B1(n_232),
.B2(n_247),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_163),
.B1(n_139),
.B2(n_153),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_218),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_146),
.B1(n_160),
.B2(n_177),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_199),
.Y(n_274)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g276 ( 
.A(n_204),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_140),
.A2(n_177),
.B1(n_142),
.B2(n_156),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_133),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_209),
.Y(n_269)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_209),
.B(n_222),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_189),
.B1(n_149),
.B2(n_131),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_210),
.A2(n_229),
.B1(n_237),
.B2(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_138),
.A2(n_134),
.B1(n_121),
.B2(n_120),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_120),
.A2(n_121),
.B1(n_134),
.B2(n_157),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_219),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_262)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_224),
.Y(n_292)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_227),
.Y(n_253)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_145),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_230),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_148),
.A2(n_187),
.B1(n_183),
.B2(n_157),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_236),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_136),
.B1(n_155),
.B2(n_167),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_171),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_234),
.B(n_194),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_148),
.A2(n_187),
.B1(n_183),
.B2(n_174),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_136),
.A2(n_132),
.B(n_137),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_241),
.B(n_217),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_166),
.A2(n_171),
.B1(n_174),
.B2(n_155),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_137),
.A2(n_168),
.B(n_123),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_119),
.A2(n_150),
.B1(n_167),
.B2(n_168),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_150),
.A2(n_152),
.B1(n_146),
.B2(n_160),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_138),
.B(n_160),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_163),
.B1(n_128),
.B2(n_126),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_117),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_251),
.B1(n_194),
.B2(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_235),
.Y(n_268)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_117),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_203),
.B(n_214),
.C(n_196),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_256),
.B(n_283),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_261),
.A2(n_278),
.B1(n_293),
.B2(n_216),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_213),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_275),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_272),
.A2(n_296),
.B(n_276),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_239),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_287),
.B1(n_249),
.B2(n_251),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_200),
.A2(n_241),
.B1(n_247),
.B2(n_220),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_216),
.B1(n_220),
.B2(n_204),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_203),
.B(n_200),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_289),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_207),
.B(n_191),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_247),
.B1(n_240),
.B2(n_216),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_266),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_199),
.B(n_248),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_208),
.B(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_247),
.A2(n_216),
.B1(n_220),
.B2(n_233),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_238),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_289),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_303),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_223),
.B(n_226),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_307),
.B(n_328),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_254),
.B1(n_296),
.B2(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_316),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_254),
.A2(n_212),
.B1(n_224),
.B2(n_278),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_297),
.B(n_260),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_262),
.A2(n_261),
.B1(n_256),
.B2(n_252),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_252),
.B1(n_281),
.B2(n_257),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_269),
.A2(n_264),
.B(n_253),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_311),
.A2(n_267),
.B(n_277),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_313),
.B(n_330),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_258),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_319),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_259),
.A2(n_265),
.B1(n_264),
.B2(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_276),
.A2(n_285),
.B1(n_271),
.B2(n_292),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_259),
.A2(n_265),
.B1(n_286),
.B2(n_271),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_292),
.B1(n_277),
.B2(n_290),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_274),
.Y(n_333)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_274),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_330),
.Y(n_351)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_274),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_279),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_279),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_335),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_354),
.B1(n_347),
.B2(n_337),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_342),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_340),
.A2(n_302),
.B(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_315),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_316),
.C(n_329),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_344),
.B(n_349),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_320),
.B(n_304),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_346),
.B(n_311),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_310),
.Y(n_349)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_352),
.A2(n_307),
.B1(n_306),
.B2(n_312),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_356),
.A2(n_365),
.B1(n_339),
.B2(n_336),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_336),
.A2(n_303),
.B1(n_300),
.B2(n_328),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_361),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_360),
.A2(n_375),
.B(n_340),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_351),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_363),
.Y(n_377)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_332),
.A2(n_312),
.B1(n_304),
.B2(n_322),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_372),
.C(n_374),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_327),
.B1(n_317),
.B2(n_318),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_368),
.A2(n_369),
.B1(n_371),
.B2(n_332),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_331),
.B1(n_323),
.B2(n_324),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_331),
.B1(n_330),
.B2(n_326),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_326),
.C(n_321),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_350),
.C(n_338),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_321),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_344),
.Y(n_376)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_390),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_370),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_392),
.B1(n_369),
.B2(n_353),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_367),
.B(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_350),
.C(n_342),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_389),
.C(n_378),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_336),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_368),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_350),
.C(n_359),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_341),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_356),
.B1(n_366),
.B2(n_345),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_395),
.A2(n_357),
.B1(n_381),
.B2(n_385),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_359),
.Y(n_397)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_384),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_353),
.B(n_355),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_403),
.Y(n_409)
);

NOR3xp33_ASAP7_75t_SL g403 ( 
.A(n_376),
.B(n_341),
.C(n_366),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_362),
.C(n_353),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_382),
.C(n_385),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_407),
.B(n_386),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_416),
.C(n_407),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_389),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_411),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_392),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_417),
.B1(n_418),
.B2(n_381),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_362),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_404),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_395),
.A2(n_402),
.B1(n_394),
.B2(n_400),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_394),
.B(n_399),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_419),
.A2(n_424),
.B(n_421),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_422),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_358),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_413),
.A2(n_402),
.B1(n_400),
.B2(n_396),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_423),
.B(n_425),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_401),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_427),
.B(n_391),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_408),
.C(n_416),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_428),
.B(n_430),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_411),
.C(n_418),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_419),
.B(n_403),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_433),
.B(n_391),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_434),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_429),
.A2(n_424),
.B(n_426),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_436),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_437),
.B(n_438),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_435),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_428),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_444),
.Y(n_445)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_431),
.B(n_439),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_440),
.B1(n_434),
.B2(n_387),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_340),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g448 ( 
.A(n_447),
.Y(n_448)
);


endmodule