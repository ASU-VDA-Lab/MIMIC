module fake_jpeg_7058_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_37),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_46),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_11),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_34),
.B(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_57),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_1),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_92),
.Y(n_119)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_23),
.B1(n_35),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_68),
.B1(n_74),
.B2(n_24),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_35),
.B1(n_19),
.B2(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_67),
.A2(n_73),
.B1(n_80),
.B2(n_89),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_35),
.B1(n_26),
.B2(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_16),
.B1(n_26),
.B2(n_27),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_19),
.B1(n_16),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_19),
.B1(n_27),
.B2(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_105),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_32),
.B1(n_27),
.B2(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_28),
.B1(n_37),
.B2(n_18),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_88),
.B1(n_30),
.B2(n_29),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_91),
.A2(n_106),
.B1(n_24),
.B2(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_1),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_104),
.Y(n_132)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_10),
.Y(n_134)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_1),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_10),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_111),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_121),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_2),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_133),
.B1(n_78),
.B2(n_87),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_24),
.B1(n_52),
.B2(n_4),
.Y(n_133)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_105),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_137),
.Y(n_165)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_24),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_93),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_76),
.B1(n_96),
.B2(n_70),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_86),
.B(n_108),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_155),
.B(n_123),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_86),
.C(n_64),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_154),
.C(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_144),
.A2(n_147),
.B1(n_103),
.B2(n_90),
.Y(n_202)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_152),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_71),
.B1(n_85),
.B2(n_96),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_148),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_158),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_117),
.B1(n_70),
.B2(n_63),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_64),
.C(n_104),
.Y(n_154)
);

OR2x4_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_122),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_77),
.B(n_100),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_92),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_172),
.Y(n_190)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_69),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_117),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_102),
.C(n_101),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_61),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_62),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_126),
.A2(n_120),
.B1(n_135),
.B2(n_121),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_139),
.B1(n_130),
.B2(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_94),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_2),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_107),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_184),
.B1(n_205),
.B2(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_139),
.C(n_130),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_161),
.C(n_169),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_115),
.B1(n_107),
.B2(n_112),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_192),
.B(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_194),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_199),
.B(n_6),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_197),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_141),
.B1(n_112),
.B2(n_111),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_129),
.B(n_141),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_170),
.B(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_178),
.B1(n_159),
.B2(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_215),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_103),
.B1(n_90),
.B2(n_136),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_4),
.C(n_5),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_164),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_150),
.A2(n_178),
.B1(n_167),
.B2(n_144),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_5),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_217),
.A2(n_218),
.B(n_227),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_195),
.A2(n_142),
.B(n_143),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_159),
.B(n_158),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_244),
.C(n_180),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_146),
.B1(n_152),
.B2(n_157),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_6),
.B1(n_8),
.B2(n_206),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_193),
.A2(n_166),
.B(n_8),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_206),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_136),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_179),
.B1(n_184),
.B2(n_189),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_250),
.C(n_267),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_214),
.A3(n_207),
.B1(n_181),
.B2(n_180),
.C1(n_208),
.C2(n_209),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_263),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_213),
.B1(n_183),
.B2(n_215),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_257),
.B(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_182),
.C(n_190),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_201),
.B(n_190),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_258),
.B(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

AO22x1_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_6),
.B1(n_8),
.B2(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_221),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_266),
.B1(n_241),
.B2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_251),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_221),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_229),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_222),
.A2(n_217),
.B1(n_231),
.B2(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_227),
.C(n_231),
.Y(n_267)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_271),
.A2(n_272),
.B1(n_286),
.B2(n_253),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_236),
.B1(n_234),
.B2(n_240),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_266),
.B1(n_252),
.B2(n_258),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_225),
.CI(n_219),
.CON(n_275),
.SN(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_225),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_219),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_265),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_233),
.C(n_229),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_233),
.B(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_247),
.C(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_295),
.C(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_267),
.B1(n_261),
.B2(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_275),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_249),
.B1(n_254),
.B2(n_239),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_299),
.B(n_271),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_246),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_313),
.B(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_278),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_268),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_280),
.C(n_274),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_296),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_306),
.B(n_313),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_320),
.B(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_279),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_270),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_275),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_293),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_277),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_254),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_323),
.C(n_223),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_314),
.B(n_318),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_332),
.C(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_289),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

AOI321xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_331),
.A3(n_276),
.B1(n_289),
.B2(n_295),
.C(n_333),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_272),
.B(n_276),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_237),
.Y(n_338)
);


endmodule