module fake_jpeg_10730_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_90),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_75),
.B1(n_58),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_77),
.B1(n_63),
.B2(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_79),
.B1(n_61),
.B2(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_67),
.B1(n_54),
.B2(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_73),
.B1(n_78),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_66),
.B1(n_59),
.B2(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_80),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_65),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_120),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_70),
.B(n_60),
.C(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_13),
.Y(n_139)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_59),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_55),
.B1(n_53),
.B2(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_128),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_68),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_0),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_126),
.Y(n_145)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_1),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_136),
.B1(n_143),
.B2(n_18),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_14),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_32),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_15),
.B(n_17),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_26),
.B(n_30),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_107),
.B1(n_118),
.B2(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_157),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_21),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_22),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_23),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2x1_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_24),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_165),
.B(n_146),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_31),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_174),
.C(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_147),
.C(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_163),
.B1(n_173),
.B2(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_182),
.B1(n_183),
.B2(n_176),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_180),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_159),
.B1(n_130),
.B2(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_143),
.C(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_185),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_184),
.B1(n_186),
.B2(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_172),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_157),
.C(n_35),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_34),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_164),
.Y(n_195)
);


endmodule