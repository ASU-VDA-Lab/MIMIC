module real_jpeg_33843_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OR2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_25),
.Y(n_43)
);

NAND2x1p5_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_12),
.Y(n_11)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_2),
.B(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_34),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g12 ( 
.A1(n_4),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_35),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_15),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OR2x6_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_21),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);


endmodule