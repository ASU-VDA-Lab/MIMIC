module fake_jpeg_14046_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_7),
.B(n_9),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_0),
.CON(n_65),
.SN(n_65)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_98),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_78),
.Y(n_145)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_49),
.Y(n_161)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_40),
.B(n_23),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_161),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_61),
.A2(n_48),
.B1(n_37),
.B2(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_122),
.B1(n_125),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_23),
.B1(n_37),
.B2(n_48),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_66),
.A2(n_37),
.B1(n_48),
.B2(n_45),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_129),
.A2(n_106),
.B1(n_97),
.B2(n_89),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_45),
.B1(n_50),
.B2(n_40),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_54),
.A2(n_19),
.B1(n_42),
.B2(n_33),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_137),
.A2(n_144),
.B1(n_146),
.B2(n_162),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_70),
.A2(n_45),
.B1(n_50),
.B2(n_65),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_60),
.A2(n_45),
.B1(n_50),
.B2(n_49),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_55),
.A2(n_49),
.B1(n_32),
.B2(n_51),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_39),
.B1(n_105),
.B2(n_92),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_82),
.B(n_19),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_155),
.B(n_156),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_42),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_64),
.A2(n_68),
.B1(n_49),
.B2(n_81),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_164),
.B(n_86),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_79),
.B(n_33),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_168),
.B(n_86),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_114),
.B(n_73),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_171),
.B(n_177),
.Y(n_260)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_24),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_173),
.B(n_175),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_24),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_176),
.B(n_193),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_115),
.A2(n_51),
.B(n_43),
.C(n_25),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_203),
.Y(n_234)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_93),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_183),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_184),
.A2(n_194),
.B1(n_160),
.B2(n_36),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_111),
.B(n_39),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_185),
.B(n_198),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_123),
.B(n_98),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_154),
.C(n_167),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_57),
.B1(n_90),
.B2(n_88),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_233),
.B1(n_146),
.B2(n_162),
.Y(n_243)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_56),
.B1(n_87),
.B2(n_80),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_133),
.B(n_25),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_120),
.A2(n_43),
.B1(n_83),
.B2(n_76),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_215),
.B1(n_216),
.B2(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_200),
.B(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_212),
.Y(n_240)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_113),
.Y(n_210)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_0),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_218),
.Y(n_262)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_221),
.Y(n_246)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_119),
.B(n_0),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_R g252 ( 
.A(n_224),
.B(n_231),
.Y(n_252)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_154),
.B(n_62),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_36),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_230),
.A2(n_232),
.B1(n_120),
.B2(n_128),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_110),
.A2(n_74),
.B1(n_58),
.B2(n_67),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_203),
.B1(n_231),
.B2(n_118),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_241),
.A2(n_265),
.B1(n_187),
.B2(n_208),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_173),
.A2(n_175),
.B1(n_185),
.B2(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_242),
.A2(n_243),
.B1(n_256),
.B2(n_266),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_211),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_201),
.A2(n_128),
.B1(n_148),
.B2(n_124),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_254),
.A2(n_255),
.B1(n_204),
.B2(n_209),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_148),
.B1(n_170),
.B2(n_149),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_110),
.B1(n_140),
.B2(n_163),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_183),
.A2(n_178),
.B1(n_213),
.B2(n_198),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_261),
.A2(n_270),
.B(n_192),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_191),
.A2(n_127),
.B(n_95),
.C(n_78),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_264),
.B(n_172),
.C(n_187),
.Y(n_289)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_194),
.A2(n_150),
.B1(n_166),
.B2(n_140),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_177),
.A2(n_166),
.B1(n_150),
.B2(n_163),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_178),
.A2(n_160),
.B1(n_170),
.B2(n_149),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_267),
.A2(n_277),
.B1(n_233),
.B2(n_235),
.Y(n_305)
);

AOI32xp33_ASAP7_75t_L g270 ( 
.A1(n_178),
.A2(n_127),
.A3(n_72),
.B1(n_71),
.B2(n_91),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_280),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_184),
.A2(n_36),
.B1(n_100),
.B2(n_17),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_183),
.B(n_36),
.C(n_17),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_188),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_289),
.A2(n_298),
.B1(n_332),
.B2(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_251),
.A2(n_190),
.B1(n_227),
.B2(n_182),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_294),
.A2(n_309),
.B(n_310),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_252),
.A2(n_224),
.B(n_214),
.Y(n_295)
);

OAI31xp33_ASAP7_75t_L g351 ( 
.A1(n_295),
.A2(n_266),
.A3(n_280),
.B(n_247),
.Y(n_351)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_262),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_312),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_299),
.B(n_300),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_174),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_270),
.A2(n_218),
.B1(n_220),
.B2(n_181),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_302),
.A2(n_337),
.B(n_257),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_249),
.B(n_210),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_321),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_317),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_252),
.A2(n_180),
.B1(n_189),
.B2(n_216),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_215),
.B1(n_206),
.B2(n_225),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_228),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_308),
.B(n_313),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_240),
.A2(n_217),
.B(n_186),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_246),
.B(n_192),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_314),
.A2(n_284),
.B(n_236),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_244),
.C(n_249),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_315),
.B(n_320),
.C(n_324),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_323),
.B1(n_327),
.B2(n_253),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_261),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_244),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_318),
.A2(n_319),
.B1(n_329),
.B2(n_330),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_277),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_278),
.B(n_17),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_242),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_1),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_325),
.Y(n_349)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_328),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_256),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_239),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_264),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_238),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_332),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_334),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_239),
.B(n_234),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_6),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_8),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_243),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_338),
.B1(n_253),
.B2(n_285),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_248),
.A2(n_11),
.B1(n_13),
.B2(n_10),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_264),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_342),
.B(n_346),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_308),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_309),
.B1(n_290),
.B2(n_292),
.Y(n_394)
);

OAI21xp33_ASAP7_75t_L g411 ( 
.A1(n_351),
.A2(n_263),
.B(n_269),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_335),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_379),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_296),
.A2(n_264),
.B1(n_245),
.B2(n_283),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_353),
.A2(n_373),
.B1(n_318),
.B2(n_328),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_248),
.B1(n_262),
.B2(n_257),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_354),
.A2(n_360),
.B(n_377),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_329),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_264),
.B1(n_247),
.B2(n_285),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_358),
.A2(n_364),
.B1(n_382),
.B2(n_289),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_336),
.A2(n_314),
.B1(n_294),
.B2(n_302),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_380),
.B(n_337),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_295),
.A2(n_286),
.B1(n_275),
.B2(n_276),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_281),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_365),
.B(n_368),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_276),
.C(n_272),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_370),
.C(n_312),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_286),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_369),
.B(n_374),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_272),
.C(n_286),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_371),
.B(n_375),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_296),
.A2(n_263),
.B1(n_273),
.B2(n_257),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_303),
.B(n_250),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_314),
.A2(n_269),
.B1(n_263),
.B2(n_282),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_297),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_314),
.A2(n_284),
.B(n_263),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_338),
.A2(n_330),
.B1(n_307),
.B2(n_310),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_383),
.A2(n_386),
.B1(n_390),
.B2(n_394),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_289),
.B(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_393),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_360),
.A2(n_301),
.B1(n_300),
.B2(n_299),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_372),
.A2(n_353),
.B1(n_367),
.B2(n_346),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_387),
.A2(n_400),
.B(n_417),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_347),
.A2(n_323),
.B1(n_316),
.B2(n_313),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_321),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_397),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_382),
.A2(n_319),
.B1(n_333),
.B2(n_325),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_396),
.A2(n_405),
.B1(n_393),
.B2(n_383),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_339),
.Y(n_398)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_293),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_407),
.C(n_410),
.Y(n_421)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_405),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_345),
.B(n_317),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_403),
.B(n_414),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_404),
.A2(n_406),
.B1(n_419),
.B2(n_340),
.Y(n_449)
);

INVx3_ASAP7_75t_SL g405 ( 
.A(n_358),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_363),
.A2(n_331),
.B1(n_326),
.B2(n_328),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_236),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_355),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_409),
.Y(n_422)
);

HB1xp67_ASAP7_75t_SL g444 ( 
.A(n_411),
.Y(n_444)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_349),
.B(n_304),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_415),
.Y(n_435)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_418),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_350),
.A2(n_304),
.B(n_282),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_258),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_342),
.A2(n_275),
.B1(n_273),
.B2(n_258),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_366),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_434),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_SL g426 ( 
.A1(n_394),
.A2(n_350),
.B(n_351),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_426),
.B(n_427),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_386),
.A2(n_361),
.B1(n_370),
.B2(n_359),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_345),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_451),
.C(n_403),
.Y(n_455)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_366),
.C(n_368),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_433),
.C(n_440),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_374),
.C(n_359),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_378),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_385),
.A2(n_344),
.B1(n_343),
.B2(n_377),
.Y(n_436)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_389),
.B(n_378),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_437),
.B(n_388),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_385),
.A2(n_344),
.B1(n_343),
.B2(n_357),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_439),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_385),
.A2(n_380),
.B1(n_381),
.B2(n_356),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_375),
.C(n_340),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_391),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_418),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_389),
.B(n_402),
.C(n_384),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_448),
.C(n_354),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_384),
.B(n_364),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_449),
.A2(n_405),
.B1(n_396),
.B2(n_390),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_371),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_453),
.A2(n_459),
.B1(n_463),
.B2(n_474),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_471),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_460),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_387),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_476),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_449),
.A2(n_431),
.B1(n_446),
.B2(n_441),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_443),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_446),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_462),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_447),
.B(n_391),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_431),
.A2(n_409),
.B1(n_397),
.B2(n_404),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_443),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_467),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_468),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_408),
.B(n_400),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_469),
.A2(n_442),
.B(n_420),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_450),
.A2(n_417),
.B(n_406),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_470),
.A2(n_472),
.B(n_435),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_437),
.B(n_415),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_SL g472 ( 
.A1(n_444),
.A2(n_408),
.B(n_401),
.C(n_416),
.Y(n_472)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_473),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_444),
.A2(n_414),
.B1(n_413),
.B2(n_398),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_422),
.A2(n_412),
.B1(n_381),
.B2(n_419),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_475),
.A2(n_430),
.B1(n_439),
.B2(n_429),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_376),
.C(n_362),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_421),
.C(n_424),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_422),
.B(n_379),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_480),
.B(n_442),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_453),
.A2(n_438),
.B1(n_429),
.B2(n_436),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_483),
.A2(n_489),
.B1(n_466),
.B2(n_458),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_487),
.A2(n_472),
.B1(n_479),
.B2(n_475),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_459),
.A2(n_435),
.B1(n_427),
.B2(n_426),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_456),
.C(n_457),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_496),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_434),
.C(n_440),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_494),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_425),
.B1(n_448),
.B2(n_445),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_493),
.A2(n_500),
.B1(n_504),
.B2(n_474),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_425),
.C(n_452),
.Y(n_494)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_420),
.Y(n_499)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_478),
.A2(n_348),
.B1(n_362),
.B2(n_273),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_348),
.B(n_11),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_502),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_8),
.C(n_10),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_469),
.A2(n_11),
.B(n_8),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_496),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_458),
.B1(n_473),
.B2(n_463),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_522),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_456),
.C(n_476),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_513),
.C(n_517),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_511),
.A2(n_519),
.B1(n_504),
.B2(n_501),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_479),
.C(n_472),
.Y(n_513)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_515),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_488),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_516),
.B(n_518),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_486),
.C(n_489),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_454),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_471),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_497),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_472),
.C(n_498),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_523),
.C(n_495),
.Y(n_535)
);

FAx1_ASAP7_75t_SL g522 ( 
.A(n_497),
.B(n_472),
.CI(n_491),
.CON(n_522),
.SN(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_493),
.C(n_482),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_532),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_505),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_531),
.Y(n_542)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_484),
.B(n_499),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_530),
.A2(n_534),
.B(n_515),
.Y(n_545)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_537),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_521),
.A2(n_484),
.B(n_513),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_535),
.B(n_487),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_485),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_536),
.A2(n_508),
.B(n_522),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_482),
.C(n_483),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_507),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_522),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_520),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_541),
.B(n_550),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_510),
.C(n_506),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_536),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_544),
.B(n_533),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_545),
.A2(n_525),
.B(n_526),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_528),
.A2(n_519),
.B1(n_485),
.B2(n_500),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_547),
.A2(n_527),
.B1(n_539),
.B2(n_528),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_549),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_502),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_526),
.C(n_537),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_553),
.Y(n_558)
);

AOI21xp33_ASAP7_75t_L g560 ( 
.A1(n_554),
.A2(n_556),
.B(n_557),
.Y(n_560)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_555),
.B(n_546),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_545),
.B(n_552),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_540),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_540),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_562),
.B(n_563),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_558),
.A2(n_552),
.B(n_542),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_R g565 ( 
.A(n_564),
.B(n_542),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_565),
.B(n_560),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_566),
.C(n_538),
.Y(n_568)
);

OAI311xp33_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_531),
.A3(n_547),
.B1(n_539),
.C1(n_532),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_503),
.Y(n_570)
);


endmodule