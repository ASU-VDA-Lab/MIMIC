module fake_jpeg_28125_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_1),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_37),
.B1(n_41),
.B2(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_42),
.B1(n_51),
.B2(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_48),
.B1(n_44),
.B2(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_45),
.B1(n_40),
.B2(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_46),
.B1(n_39),
.B2(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_83),
.Y(n_100)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_71),
.B1(n_65),
.B2(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_87),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_2),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_20),
.A3(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_98),
.B1(n_81),
.B2(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_103),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_83),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_105),
.B(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_23),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_94),
.C(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_7),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_91),
.B(n_95),
.C(n_24),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_112),
.B1(n_10),
.B2(n_11),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_91),
.B(n_19),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_111),
.C(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_113),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_17),
.B(n_18),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_25),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_26),
.Y(n_126)
);


endmodule