module fake_ariane_375_n_2437 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2437);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2437;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_352;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2415;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_374;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2375;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_369;
wire n_240;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g233 ( 
.A(n_109),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_216),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_49),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_130),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_113),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_198),
.Y(n_245)
);

INVx4_ASAP7_75t_R g246 ( 
.A(n_139),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_141),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_43),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_127),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_142),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_63),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_101),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_144),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_37),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_23),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_156),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_103),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_221),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_100),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_138),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_84),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_110),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_217),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_56),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_105),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_189),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_195),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_184),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_157),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_84),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_81),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_7),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_21),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_229),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_218),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_0),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_166),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_83),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_40),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_131),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_93),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_92),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_82),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_27),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_96),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_25),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_199),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_72),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_16),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_231),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_48),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_85),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_103),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_213),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_61),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_165),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_168),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_208),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_107),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_80),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_215),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_78),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_188),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_37),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_115),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_128),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_19),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_94),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_8),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_13),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_64),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_91),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_89),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_59),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_191),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_28),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_34),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_171),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_147),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_78),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_49),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_160),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_31),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_29),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_26),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_211),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_117),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_44),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_62),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_11),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_39),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_3),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_64),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_161),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_83),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_145),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_17),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_88),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_42),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_17),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_42),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_46),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_47),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_121),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_111),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_118),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_73),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_53),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_52),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_58),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_58),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_219),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_135),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_182),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_60),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_48),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_18),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_12),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_97),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_16),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_149),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_192),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_46),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_151),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_159),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_230),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_23),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_175),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_97),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_126),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_65),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_1),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_91),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_90),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_53),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_34),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_98),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_4),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_190),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_106),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_180),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_15),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_173),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_129),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_92),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_183),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_136),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_28),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_96),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_116),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_102),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_33),
.Y(n_427)
);

BUFx10_ASAP7_75t_L g428 ( 
.A(n_57),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_35),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_19),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_26),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_32),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_30),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_57),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_206),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_29),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_55),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_227),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_14),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_68),
.Y(n_440)
);

BUFx2_ASAP7_75t_SL g441 ( 
.A(n_61),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_87),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_22),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_71),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_12),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_47),
.Y(n_446)
);

BUFx5_ASAP7_75t_L g447 ( 
.A(n_112),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_93),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_201),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_203),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_86),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_124),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_35),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_210),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_66),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_202),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_5),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_369),
.B(n_233),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_261),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_369),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_233),
.B(n_1),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_290),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_252),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_252),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_255),
.B(n_2),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_255),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_256),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_298),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_325),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_256),
.B(n_2),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_260),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_403),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_365),
.B(n_3),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_260),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_265),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_265),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_452),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_376),
.B(n_5),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_376),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_266),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_266),
.B(n_6),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_249),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_267),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_258),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_292),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_267),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_269),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_263),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_264),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_303),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_269),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_307),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_273),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_273),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_295),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_308),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_307),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_358),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_364),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_300),
.B(n_7),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_270),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_276),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_277),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_278),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_277),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_294),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_294),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_371),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_280),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_304),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_304),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_316),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_316),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_408),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_335),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_324),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_324),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_411),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_282),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_242),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_330),
.B(n_9),
.Y(n_525)
);

INVx4_ASAP7_75t_R g526 ( 
.A(n_246),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_330),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_334),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_288),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_334),
.B(n_9),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_291),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_424),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_337),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_429),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_307),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_337),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_347),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_347),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_360),
.B(n_10),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_296),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_305),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_243),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_360),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_303),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_433),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_379),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_335),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_437),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_306),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_335),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_362),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_379),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_310),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_387),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_250),
.B(n_10),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_312),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_303),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_236),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_387),
.B(n_11),
.Y(n_559)
);

INVxp33_ASAP7_75t_SL g560 ( 
.A(n_341),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_321),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_236),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_389),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_326),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_389),
.B(n_14),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_415),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_327),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_415),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_329),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_243),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_332),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_236),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_341),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_250),
.B(n_272),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_339),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_362),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_307),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_307),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_422),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_461),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_495),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_524),
.B(n_238),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_485),
.B(n_239),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_471),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_500),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_488),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_535),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_480),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_470),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_459),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_460),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_474),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_579),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_462),
.B(n_362),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_460),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_498),
.Y(n_607)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_493),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_487),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_491),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_458),
.B(n_422),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_499),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_492),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_560),
.B(n_425),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_442),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_580),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_544),
.B(n_234),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_469),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_473),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_425),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_475),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_504),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_477),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_477),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_478),
.B(n_442),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_505),
.B(n_340),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_507),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_479),
.A2(n_456),
.B(n_438),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_512),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_557),
.B(n_234),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_479),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_523),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_529),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_518),
.B(n_438),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_531),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_481),
.A2(n_359),
.B1(n_367),
.B2(n_262),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_540),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_486),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_501),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_486),
.Y(n_647)
);

OA21x2_ASAP7_75t_L g648 ( 
.A1(n_489),
.A2(n_456),
.B(n_381),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_489),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_541),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_549),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_494),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_494),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_496),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_496),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_575),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_497),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_497),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_506),
.Y(n_663)
);

NAND2x1_ASAP7_75t_L g664 ( 
.A(n_526),
.B(n_246),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_508),
.B(n_442),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_508),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_509),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_553),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_509),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_561),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_564),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_510),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_511),
.Y(n_675)
);

CKINVDCx16_ASAP7_75t_R g676 ( 
.A(n_464),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_551),
.B(n_245),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_513),
.B(n_245),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_603),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_643),
.A2(n_641),
.B1(n_616),
.B2(n_481),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_574),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_603),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_666),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_625),
.B(n_522),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_666),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_666),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_584),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_616),
.B(n_677),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_322),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_604),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_584),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_601),
.B(n_578),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_622),
.B(n_567),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_604),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_658),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_584),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_591),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_606),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_590),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_609),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_476),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_625),
.B(n_502),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_476),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_601),
.B(n_617),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_669),
.B(n_586),
.Y(n_708)
);

NAND2x1p5_ASAP7_75t_L g709 ( 
.A(n_664),
.B(n_648),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_658),
.B(n_569),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_658),
.B(n_571),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_666),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_666),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_590),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_669),
.B(n_577),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_621),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_597),
.B(n_322),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_677),
.B(n_513),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_619),
.B(n_514),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_621),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_666),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_658),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_613),
.B(n_547),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_610),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_623),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_623),
.Y(n_726)
);

NAND2x1p5_ASAP7_75t_L g727 ( 
.A(n_664),
.B(n_648),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_613),
.B(n_550),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_619),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_619),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_629),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_622),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_605),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_622),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_602),
.B(n_322),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_611),
.Y(n_736)
);

INVx4_ASAP7_75t_SL g737 ( 
.A(n_622),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_582),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_637),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_605),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_629),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_602),
.B(n_355),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_637),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_622),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_618),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_619),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_631),
.A2(n_467),
.B1(n_525),
.B2(n_472),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_640),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_640),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_645),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_615),
.A2(n_463),
.B1(n_530),
.B2(n_484),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_628),
.B(n_647),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_622),
.B(n_251),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_628),
.B(n_514),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_622),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_542),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_631),
.A2(n_539),
.B1(n_559),
.B2(n_558),
.Y(n_759)
);

INVxp33_ASAP7_75t_SL g760 ( 
.A(n_626),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_608),
.B(n_555),
.Y(n_761)
);

BUFx4f_ASAP7_75t_L g762 ( 
.A(n_649),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_653),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_628),
.B(n_515),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_608),
.B(n_570),
.Y(n_765)
);

INVx8_ASAP7_75t_L g766 ( 
.A(n_617),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_653),
.B(n_355),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_649),
.B(n_251),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_654),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_628),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_649),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_617),
.B(n_570),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_381),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_632),
.B(n_562),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_649),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_634),
.Y(n_777)
);

BUFx8_ASAP7_75t_SL g778 ( 
.A(n_607),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_638),
.A2(n_565),
.B1(n_503),
.B2(n_555),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_639),
.B(n_573),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_629),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_655),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_647),
.B(n_515),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_589),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_617),
.B(n_516),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_647),
.B(n_516),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_649),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_618),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_642),
.A2(n_650),
.B1(n_651),
.B2(n_644),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_618),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_647),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_649),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_665),
.B(n_519),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_649),
.B(n_652),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_652),
.B(n_519),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_660),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_665),
.B(n_520),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_660),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_652),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_652),
.B(n_520),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_643),
.A2(n_300),
.B1(n_353),
.B2(n_309),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_657),
.B(n_527),
.Y(n_802)
);

NOR2x1p5_ASAP7_75t_L g803 ( 
.A(n_668),
.B(n_672),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_657),
.B(n_527),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_662),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_583),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_657),
.Y(n_807)
);

AO22x2_ASAP7_75t_L g808 ( 
.A1(n_620),
.A2(n_575),
.B1(n_533),
.B2(n_536),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_673),
.B(n_528),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_662),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_667),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_667),
.Y(n_812)
);

AND2x6_ASAP7_75t_L g813 ( 
.A(n_670),
.B(n_528),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_670),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_594),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_595),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_657),
.B(n_533),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_648),
.B(n_536),
.Y(n_818)
);

AND2x6_ASAP7_75t_L g819 ( 
.A(n_674),
.B(n_537),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_587),
.B(n_659),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_595),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_674),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

AND2x2_ASAP7_75t_SL g824 ( 
.A(n_633),
.B(n_648),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_659),
.B(n_641),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_648),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_665),
.B(n_537),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_L g828 ( 
.A1(n_678),
.A2(n_309),
.B1(n_385),
.B2(n_353),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_659),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_588),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_627),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_627),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_595),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_583),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_595),
.B(n_538),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_598),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_678),
.B(n_538),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_583),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_816),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_688),
.A2(n_731),
.B(n_781),
.C(n_741),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_825),
.B(n_838),
.Y(n_843)
);

NAND2x1_ASAP7_75t_L g844 ( 
.A(n_813),
.B(n_598),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_825),
.B(n_598),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_816),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_838),
.B(n_598),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_838),
.B(n_587),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_687),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_816),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_687),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_729),
.B(n_630),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_710),
.B(n_635),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_710),
.B(n_676),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_681),
.B(n_630),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_821),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_680),
.A2(n_343),
.B1(n_624),
.B2(n_630),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_681),
.B(n_636),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_729),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_729),
.B(n_636),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_731),
.A2(n_624),
.B(n_656),
.C(n_636),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_730),
.B(n_656),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_723),
.B(n_656),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_723),
.B(n_663),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_728),
.B(n_663),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_L g867 ( 
.A1(n_748),
.A2(n_385),
.B1(n_455),
.B2(n_349),
.C(n_346),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_728),
.B(n_663),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_711),
.B(n_676),
.Y(n_869)
);

NOR2x2_ASAP7_75t_L g870 ( 
.A(n_760),
.B(n_661),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_691),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_708),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_821),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_691),
.Y(n_874)
);

NAND2x1_ASAP7_75t_L g875 ( 
.A(n_813),
.B(n_671),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_718),
.B(n_711),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_766),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_692),
.B(n_671),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_722),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_692),
.B(n_671),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_759),
.B(n_809),
.C(n_789),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_707),
.A2(n_661),
.B1(n_633),
.B2(n_546),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_760),
.B(n_596),
.Y(n_883)
);

BUFx4_ASAP7_75t_L g884 ( 
.A(n_778),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_730),
.B(n_585),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_833),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_766),
.B(n_661),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_707),
.A2(n_633),
.B1(n_546),
.B2(n_552),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_730),
.B(n_747),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_696),
.A2(n_345),
.B1(n_348),
.B2(n_344),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_SL g891 ( 
.A1(n_761),
.A2(n_521),
.B1(n_532),
.B2(n_517),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_764),
.A2(n_552),
.B(n_554),
.C(n_543),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_692),
.B(n_585),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_833),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_747),
.B(n_543),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_764),
.A2(n_563),
.B(n_566),
.C(n_554),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_833),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_741),
.A2(n_455),
.B(n_237),
.C(n_257),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_793),
.B(n_563),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_813),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_793),
.B(n_566),
.Y(n_901)
);

INVx8_ASAP7_75t_L g902 ( 
.A(n_766),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_697),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_807),
.A2(n_633),
.B(n_572),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_836),
.B(n_568),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_679),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_836),
.B(n_568),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_766),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_797),
.B(n_572),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_747),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_707),
.A2(n_633),
.B1(n_581),
.B2(n_576),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_722),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_765),
.B(n_715),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_797),
.B(n_576),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_761),
.B(n_705),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_797),
.B(n_581),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_703),
.A2(n_336),
.B1(n_234),
.B2(n_315),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_827),
.B(n_235),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_696),
.B(n_599),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_682),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_827),
.B(n_240),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_757),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_698),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_752),
.B(n_614),
.Y(n_924)
);

AND2x6_ASAP7_75t_SL g925 ( 
.A(n_774),
.B(n_237),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_813),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_827),
.B(n_286),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_785),
.B(n_241),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_697),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_272),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_785),
.B(n_354),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_703),
.B(n_241),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_781),
.B(n_354),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_703),
.A2(n_706),
.B1(n_826),
.B2(n_808),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_791),
.B(n_281),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_684),
.B(n_646),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_738),
.B(n_244),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_706),
.B(n_675),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_791),
.Y(n_939)
);

AND2x6_ASAP7_75t_SL g940 ( 
.A(n_780),
.B(n_257),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_690),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_706),
.B(n_394),
.Y(n_942)
);

AND2x2_ASAP7_75t_SL g943 ( 
.A(n_820),
.B(n_826),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_815),
.B(n_534),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_840),
.B(n_441),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_L g946 ( 
.A(n_813),
.B(n_281),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_779),
.B(n_545),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_791),
.B(n_281),
.Y(n_948)
);

INVx8_ASAP7_75t_L g949 ( 
.A(n_813),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_753),
.B(n_394),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_753),
.B(n_436),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_819),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_820),
.A2(n_247),
.B1(n_253),
.B2(n_248),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_802),
.A2(n_283),
.B(n_297),
.C(n_259),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_700),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_834),
.B(n_436),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_772),
.B(n_259),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_819),
.A2(n_254),
.B1(n_271),
.B2(n_268),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_738),
.B(n_274),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_SL g960 ( 
.A(n_784),
.B(n_372),
.C(n_357),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_834),
.B(n_451),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_694),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_794),
.A2(n_693),
.B(n_837),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_772),
.B(n_548),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_700),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_834),
.B(n_451),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_772),
.B(n_283),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_695),
.B(n_699),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_818),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_837),
.B(n_373),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_704),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_837),
.B(n_374),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_826),
.A2(n_234),
.B1(n_336),
.B2(n_366),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_704),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_808),
.A2(n_336),
.B1(n_428),
.B2(n_315),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_714),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_701),
.B(n_441),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_683),
.Y(n_978)
);

NAND2x1_ASAP7_75t_L g979 ( 
.A(n_819),
.B(n_588),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_702),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_824),
.B(n_281),
.Y(n_981)
);

BUFx8_ASAP7_75t_L g982 ( 
.A(n_778),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_716),
.B(n_297),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_720),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_725),
.B(n_726),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_824),
.B(n_281),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_739),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_744),
.B(n_302),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_714),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_819),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_770),
.B(n_302),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_749),
.B(n_313),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_750),
.B(n_313),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_751),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_733),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_758),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_733),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_763),
.B(n_769),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_770),
.A2(n_390),
.B1(n_457),
.B2(n_391),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_776),
.B(n_317),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_819),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_740),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_782),
.B(n_317),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_796),
.B(n_318),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_808),
.B(n_318),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_803),
.B(n_338),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_798),
.B(n_338),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_805),
.B(n_346),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_SL g1009 ( 
.A(n_784),
.B(n_336),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_810),
.B(n_349),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_811),
.B(n_363),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_819),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_801),
.B(n_363),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_740),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_767),
.A2(n_319),
.B1(n_303),
.B2(n_428),
.Y(n_1015)
);

OA22x2_ASAP7_75t_L g1016 ( 
.A1(n_891),
.A2(n_812),
.B1(n_822),
.B2(n_814),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_952),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_849),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_906),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_923),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_876),
.B(n_799),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_883),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_872),
.Y(n_1024)
);

BUFx4f_ASAP7_75t_L g1025 ( 
.A(n_902),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_949),
.B(n_799),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_915),
.B(n_724),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_902),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_853),
.B(n_724),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_952),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_920),
.Y(n_1031)
);

BUFx8_ASAP7_75t_SL g1032 ( 
.A(n_884),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_829),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_909),
.B(n_829),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_941),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_SL g1036 ( 
.A(n_938),
.B(n_377),
.C(n_375),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_902),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_SL g1038 ( 
.A1(n_924),
.A2(n_382),
.B1(n_384),
.B2(n_383),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_914),
.B(n_719),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_881),
.A2(n_736),
.B1(n_777),
.B2(n_724),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_902),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_962),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_916),
.A2(n_802),
.B(n_755),
.C(n_786),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_952),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_899),
.B(n_783),
.Y(n_1045)
);

INVxp67_ASAP7_75t_SL g1046 ( 
.A(n_879),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_1009),
.B(n_736),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_901),
.B(n_795),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_936),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_848),
.B(n_800),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_879),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_980),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_982),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_922),
.B(n_736),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_887),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_984),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_887),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_987),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_994),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_887),
.B(n_737),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_996),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_949),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_857),
.B(n_804),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_872),
.Y(n_1064)
);

OR2x4_ASAP7_75t_L g1065 ( 
.A(n_854),
.B(n_777),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_968),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_949),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_851),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_922),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_944),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_944),
.B(n_817),
.Y(n_1071)
);

INVx3_ASAP7_75t_SL g1072 ( 
.A(n_870),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_985),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_847),
.B(n_818),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_887),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_913),
.B(n_777),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_949),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_978),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_851),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_900),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_890),
.B(n_398),
.C(n_386),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_998),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_878),
.Y(n_1083)
);

NOR2x2_ASAP7_75t_L g1084 ( 
.A(n_1006),
.B(n_792),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_880),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_964),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_978),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_1006),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_889),
.A2(n_693),
.B(n_794),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_978),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_905),
.B(n_689),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_978),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_982),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_871),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_982),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_841),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_869),
.B(n_828),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_871),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_877),
.B(n_689),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_877),
.B(n_737),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1006),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_874),
.Y(n_1102)
);

NAND2x1_ASAP7_75t_L g1103 ( 
.A(n_859),
.B(n_712),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_874),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_978),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_925),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_900),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_903),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_940),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_903),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_893),
.B(n_709),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_947),
.B(n_823),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_907),
.B(n_689),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_900),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1006),
.Y(n_1115)
);

CKINVDCx14_ASAP7_75t_R g1116 ( 
.A(n_919),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_957),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_929),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_900),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_900),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_846),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_960),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_943),
.B(n_926),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_SL g1124 ( 
.A(n_867),
.B(n_410),
.C(n_404),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_929),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_845),
.B(n_689),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_850),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_855),
.B(n_689),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_858),
.B(n_689),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_955),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_856),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_908),
.B(n_737),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_945),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_865),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_970),
.B(n_717),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_873),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_957),
.B(n_315),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_918),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_886),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_943),
.B(n_745),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_894),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_972),
.A2(n_735),
.B1(n_717),
.B2(n_767),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_897),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_908),
.B(n_709),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_999),
.B(n_417),
.C(n_412),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_844),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_863),
.B(n_717),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_991),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_926),
.B(n_717),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_991),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_928),
.B(n_712),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_990),
.B(n_1001),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_991),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_967),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_921),
.B(n_727),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_859),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_927),
.B(n_727),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_990),
.B(n_1001),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_864),
.B(n_717),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_R g1161 ( 
.A(n_945),
.B(n_713),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_945),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_866),
.B(n_717),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_R g1164 ( 
.A(n_945),
.B(n_1005),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_967),
.B(n_315),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_SL g1166 ( 
.A(n_977),
.B(n_423),
.C(n_420),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_SL g1167 ( 
.A(n_953),
.B(n_431),
.C(n_427),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_983),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_884),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_928),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_979),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_928),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_868),
.A2(n_831),
.B(n_832),
.C(n_393),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_988),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_965),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_942),
.B(n_735),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_932),
.B(n_1013),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_965),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_R g1179 ( 
.A(n_1012),
.B(n_735),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_859),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1012),
.B(n_712),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_844),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_932),
.B(n_735),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_930),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_992),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1013),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_993),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_971),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_931),
.B(n_735),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_933),
.B(n_713),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_882),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_895),
.B(n_713),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1005),
.B(n_735),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_912),
.B(n_767),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_910),
.B(n_745),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_934),
.B(n_767),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1000),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_870),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1003),
.B(n_440),
.C(n_434),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_950),
.B(n_767),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_895),
.B(n_721),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_885),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1004),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1007),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_842),
.B(n_959),
.C(n_937),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1008),
.B(n_445),
.C(n_444),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_910),
.B(n_767),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1010),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_910),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1011),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_939),
.Y(n_1211)
);

AOI211x1_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_951),
.B(n_904),
.C(n_956),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1018),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1141),
.A2(n_986),
.B(n_981),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1029),
.B(n_975),
.Y(n_1215)
);

AND2x6_ASAP7_75t_L g1216 ( 
.A(n_1017),
.B(n_939),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_889),
.B(n_885),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1021),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1069),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1022),
.A2(n_939),
.B(n_935),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1045),
.A2(n_966),
.B(n_961),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1029),
.B(n_917),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1024),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_SL g1224 ( 
.A(n_1047),
.B(n_448),
.C(n_446),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1020),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1177),
.B(n_973),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1073),
.B(n_1082),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1037),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1032),
.B(n_969),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1097),
.A2(n_861),
.B(n_946),
.C(n_896),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1064),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1031),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1063),
.A2(n_946),
.B(n_896),
.C(n_892),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1141),
.A2(n_986),
.B(n_981),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1091),
.A2(n_948),
.B(n_935),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1113),
.A2(n_948),
.B(n_963),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1055),
.B(n_875),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1126),
.A2(n_860),
.B(n_852),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1054),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1048),
.A2(n_1050),
.B(n_1148),
.Y(n_1240)
);

AND2x2_ASAP7_75t_SL g1241 ( 
.A(n_1134),
.B(n_1015),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1138),
.B(n_319),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_1017),
.B(n_971),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1210),
.B(n_888),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1111),
.B(n_683),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1076),
.B(n_911),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1076),
.B(n_892),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1160),
.A2(n_1163),
.B(n_1033),
.Y(n_1248)
);

AOI21x1_ASAP7_75t_SL g1249 ( 
.A1(n_1039),
.A2(n_860),
.B(n_852),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1089),
.A2(n_979),
.B(n_976),
.Y(n_1250)
);

AO22x2_ASAP7_75t_L g1251 ( 
.A1(n_1112),
.A2(n_989),
.B1(n_1002),
.B2(n_997),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1168),
.B(n_1174),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1074),
.A2(n_862),
.B(n_762),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1192),
.A2(n_862),
.B(n_762),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1018),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1037),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1038),
.A2(n_898),
.A3(n_954),
.B1(n_754),
.B2(n_768),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1195),
.A2(n_762),
.B(n_974),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1123),
.A2(n_976),
.B(n_974),
.Y(n_1259)
);

OAI22x1_ASAP7_75t_L g1260 ( 
.A1(n_1088),
.A2(n_958),
.B1(n_409),
.B2(n_395),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1070),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1185),
.A2(n_342),
.B(n_443),
.C(n_439),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1187),
.B(n_989),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1197),
.B(n_995),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1086),
.B(n_995),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_1040),
.B(n_721),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1156),
.A2(n_768),
.B(n_754),
.Y(n_1267)
);

AOI211x1_ASAP7_75t_L g1268 ( 
.A1(n_1035),
.A2(n_409),
.B(n_443),
.C(n_378),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1123),
.A2(n_1002),
.B(n_997),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1203),
.A2(n_342),
.B(n_407),
.C(n_378),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1200),
.A2(n_792),
.B(n_1014),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1053),
.Y(n_1272)
);

O2A1O1Ixp5_ASAP7_75t_L g1273 ( 
.A1(n_1205),
.A2(n_721),
.B(n_732),
.C(n_734),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1170),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1129),
.A2(n_1014),
.B(n_734),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1195),
.A2(n_1130),
.B(n_1025),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1025),
.A2(n_734),
.B(n_732),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1176),
.A2(n_1145),
.B(n_1189),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1172),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1192),
.A2(n_1201),
.B(n_1043),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1204),
.B(n_773),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1042),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1111),
.B(n_683),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1208),
.B(n_773),
.Y(n_1284)
);

AOI211x1_ASAP7_75t_L g1285 ( 
.A1(n_1052),
.A2(n_407),
.B(n_439),
.C(n_392),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1201),
.A2(n_732),
.B(n_806),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1019),
.A2(n_839),
.B(n_806),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1165),
.B(n_319),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1027),
.B(n_773),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1117),
.B(n_773),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1019),
.A2(n_839),
.B(n_746),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1056),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1068),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1173),
.A2(n_746),
.A3(n_743),
.B(n_790),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1173),
.A2(n_1158),
.B(n_1156),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1157),
.A2(n_393),
.B(n_392),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1155),
.B(n_773),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1049),
.A2(n_1071),
.B(n_1116),
.C(n_1167),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1139),
.B(n_773),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1116),
.B(n_683),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1058),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1068),
.A2(n_788),
.B(n_743),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1062),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1101),
.B(n_319),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1062),
.B(n_1077),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1079),
.A2(n_790),
.B(n_788),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1025),
.A2(n_756),
.B(n_745),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1083),
.B(n_742),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1085),
.B(n_742),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1186),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1079),
.A2(n_1098),
.B(n_1094),
.Y(n_1311)
);

O2A1O1Ixp5_ASAP7_75t_L g1312 ( 
.A1(n_1034),
.A2(n_413),
.B(n_395),
.C(n_430),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1157),
.A2(n_756),
.B(n_745),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1032),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1157),
.A2(n_771),
.B(n_756),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1094),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1115),
.B(n_406),
.Y(n_1317)
);

AOI211x1_ASAP7_75t_L g1318 ( 
.A1(n_1059),
.A2(n_432),
.B(n_430),
.C(n_413),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1098),
.A2(n_432),
.B(n_406),
.Y(n_1319)
);

AND2x2_ASAP7_75t_SL g1320 ( 
.A(n_1134),
.B(n_307),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1149),
.B(n_742),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1158),
.A2(n_279),
.B(n_275),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1061),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1102),
.A2(n_742),
.A3(n_685),
.B(n_686),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1102),
.A2(n_1108),
.B(n_1104),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1211),
.B(n_685),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1104),
.A2(n_686),
.B(n_685),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1211),
.B(n_685),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1152),
.A2(n_453),
.B1(n_771),
.B2(n_787),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1184),
.B(n_742),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1023),
.B(n_686),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1096),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1180),
.A2(n_771),
.B(n_756),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_SL g1335 ( 
.A(n_1062),
.B(n_686),
.Y(n_1335)
);

BUFx5_ASAP7_75t_L g1336 ( 
.A(n_1026),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1062),
.B(n_771),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1124),
.B(n_426),
.C(n_775),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1191),
.B(n_742),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1191),
.B(n_775),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1152),
.B(n_775),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_SL g1342 ( 
.A1(n_1180),
.A2(n_787),
.B(n_775),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1152),
.B(n_787),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1186),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1108),
.A2(n_787),
.B(n_835),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1110),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1110),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1023),
.B(n_835),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1143),
.A2(n_426),
.B(n_333),
.C(n_612),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1180),
.A2(n_835),
.B(n_830),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1118),
.A2(n_835),
.B(n_830),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1211),
.B(n_830),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1209),
.A2(n_830),
.B(n_285),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1118),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_SL g1355 ( 
.A(n_1047),
.B(n_287),
.C(n_284),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1017),
.A2(n_426),
.B1(n_830),
.B2(n_396),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1023),
.B(n_366),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1016),
.B(n_1051),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1016),
.B(n_366),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1051),
.B(n_366),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1125),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1046),
.B(n_428),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1125),
.A2(n_588),
.B(n_600),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1121),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1209),
.A2(n_388),
.B(n_293),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1127),
.A2(n_588),
.B(n_600),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1057),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1128),
.Y(n_1368)
);

AOI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1164),
.A2(n_397),
.B(n_299),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1106),
.B(n_428),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1106),
.B(n_426),
.Y(n_1371)
);

AOI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1145),
.A2(n_612),
.B(n_593),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1127),
.A2(n_588),
.B(n_600),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1209),
.A2(n_399),
.B(n_301),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1211),
.A2(n_400),
.B(n_311),
.Y(n_1375)
);

AND3x4_ASAP7_75t_L g1376 ( 
.A(n_1093),
.B(n_20),
.C(n_22),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1132),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1162),
.B(n_24),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1131),
.A2(n_588),
.B(n_600),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1037),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1084),
.Y(n_1381)
);

INVx5_ASAP7_75t_L g1382 ( 
.A(n_1037),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1275),
.A2(n_1175),
.B(n_1131),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1275),
.A2(n_1178),
.B(n_1175),
.Y(n_1384)
);

AO32x2_ASAP7_75t_L g1385 ( 
.A1(n_1330),
.A2(n_1164),
.A3(n_1084),
.B1(n_1080),
.B2(n_1161),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1213),
.Y(n_1386)
);

CKINVDCx12_ASAP7_75t_R g1387 ( 
.A(n_1317),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1325),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1225),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1232),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1282),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1262),
.A2(n_1146),
.B1(n_1036),
.B2(n_1081),
.C(n_1109),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1292),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1325),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1305),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1367),
.B(n_1055),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1325),
.Y(n_1397)
);

BUFx2_ASAP7_75t_R g1398 ( 
.A(n_1367),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1271),
.A2(n_1221),
.B(n_1250),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1247),
.A2(n_1065),
.B1(n_1202),
.B2(n_1183),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1213),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1314),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1246),
.A2(n_1190),
.B(n_1202),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1303),
.B(n_1062),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1241),
.A2(n_1193),
.B1(n_1109),
.B2(n_1196),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1255),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1262),
.A2(n_1122),
.B1(n_1206),
.B2(n_1199),
.C(n_1166),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1280),
.A2(n_1188),
.B(n_1178),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1222),
.A2(n_1161),
.B1(n_1198),
.B2(n_1072),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1250),
.A2(n_1188),
.B(n_1044),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1219),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1372),
.A2(n_1145),
.B(n_1194),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1227),
.B(n_1072),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1301),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1248),
.A2(n_1044),
.B(n_1030),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1320),
.B(n_1135),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1311),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1287),
.A2(n_1044),
.B(n_1030),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1265),
.B(n_1137),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1272),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1241),
.A2(n_1057),
.B1(n_1075),
.B2(n_1169),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1303),
.B(n_1077),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1323),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1274),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1265),
.B(n_1140),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1287),
.A2(n_1144),
.B(n_1142),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1252),
.B(n_1065),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1278),
.A2(n_1145),
.B(n_1159),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1305),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1311),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1333),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1215),
.A2(n_1030),
.B(n_1147),
.C(n_1182),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1261),
.B(n_1075),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1226),
.A2(n_1122),
.B1(n_1093),
.B2(n_1095),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1316),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1242),
.A2(n_1057),
.B1(n_1053),
.B2(n_1026),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1320),
.B(n_1105),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1230),
.A2(n_1077),
.B1(n_1211),
.B2(n_1182),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1223),
.B(n_1105),
.Y(n_1441)
);

OAI211xp5_ASAP7_75t_L g1442 ( 
.A1(n_1298),
.A2(n_1357),
.B(n_1270),
.C(n_1288),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1382),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1346),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1291),
.A2(n_1159),
.B(n_1067),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1240),
.A2(n_1087),
.B(n_1078),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1291),
.A2(n_1067),
.B(n_1103),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1363),
.A2(n_1067),
.B(n_1171),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1231),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1363),
.A2(n_1373),
.B(n_1366),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1366),
.A2(n_1379),
.B(n_1373),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1364),
.B(n_1060),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1267),
.A2(n_1114),
.A3(n_1107),
.B(n_1171),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1276),
.A2(n_1041),
.B(n_1028),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1368),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1251),
.B(n_1060),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1237),
.B(n_1060),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1377),
.B(n_1147),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1223),
.B(n_1078),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1329),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1379),
.A2(n_1171),
.B(n_1087),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1345),
.A2(n_1171),
.B(n_1087),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1233),
.A2(n_1181),
.B(n_1133),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1254),
.A2(n_1041),
.B(n_1028),
.Y(n_1464)
);

AO31x2_ASAP7_75t_L g1465 ( 
.A1(n_1349),
.A2(n_1107),
.A3(n_1114),
.B(n_1090),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1233),
.A2(n_1181),
.B(n_1133),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1349),
.A2(n_1181),
.B(n_1080),
.Y(n_1467)
);

OAI222xp33_ASAP7_75t_L g1468 ( 
.A1(n_1359),
.A2(n_1095),
.B1(n_1133),
.B2(n_1100),
.C1(n_1107),
.C2(n_1114),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1263),
.B(n_1078),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1303),
.B(n_1077),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1272),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1347),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_SL g1473 ( 
.A(n_1237),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1229),
.A2(n_1077),
.B1(n_1119),
.B2(n_1120),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1347),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1230),
.A2(n_1100),
.B(n_1120),
.C(n_1119),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1314),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1270),
.A2(n_1100),
.B(n_1026),
.C(n_1207),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1274),
.B(n_1078),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1244),
.A2(n_1207),
.B1(n_1026),
.B2(n_1150),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1354),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1218),
.A2(n_1026),
.B(n_30),
.C(n_31),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1345),
.A2(n_1090),
.B(n_1092),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1361),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1361),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1279),
.B(n_1087),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1378),
.A2(n_1026),
.B(n_32),
.C(n_33),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1256),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1310),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1245),
.A2(n_1150),
.B(n_1179),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1236),
.A2(n_1092),
.B(n_1090),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1239),
.B(n_1090),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1327),
.A2(n_1092),
.B(n_1120),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1273),
.A2(n_401),
.B(n_314),
.Y(n_1495)
);

INVx8_ASAP7_75t_L g1496 ( 
.A(n_1382),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1237),
.B(n_1092),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1217),
.A2(n_1119),
.B(n_1120),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1256),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1279),
.B(n_1153),
.Y(n_1500)
);

AOI21xp33_ASAP7_75t_L g1501 ( 
.A1(n_1322),
.A2(n_1119),
.B(n_583),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1259),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1256),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1259),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1327),
.A2(n_1153),
.B(n_1099),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1382),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1319),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1269),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1344),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1382),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1269),
.A2(n_1099),
.B(n_1179),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1319),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1351),
.A2(n_588),
.B(n_600),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1370),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1338),
.A2(n_426),
.B(n_289),
.C(n_380),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1304),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1264),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1351),
.A2(n_600),
.B(n_612),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1214),
.A2(n_600),
.B(n_612),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1312),
.A2(n_426),
.B(n_320),
.C(n_370),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1300),
.B(n_323),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1214),
.A2(n_593),
.B(n_592),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1381),
.B(n_583),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1358),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1234),
.A2(n_593),
.B(n_592),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1300),
.B(n_328),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1302),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1289),
.A2(n_1299),
.B(n_1266),
.C(n_1281),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1251),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1302),
.Y(n_1530)
);

CKINVDCx14_ASAP7_75t_R g1531 ( 
.A(n_1371),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1251),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1306),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1235),
.A2(n_333),
.B(n_331),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1256),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1342),
.A2(n_24),
.B(n_36),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1326),
.B(n_583),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1306),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1243),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1340),
.B(n_592),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1294),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1284),
.A2(n_416),
.B(n_350),
.C(n_351),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1294),
.Y(n_1543)
);

INVx3_ASAP7_75t_SL g1544 ( 
.A(n_1380),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1253),
.A2(n_36),
.B(n_38),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1294),
.Y(n_1546)
);

AO31x2_ASAP7_75t_L g1547 ( 
.A1(n_1238),
.A2(n_593),
.A3(n_592),
.B(n_612),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1326),
.B(n_612),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1290),
.A2(n_418),
.B(n_352),
.C(n_454),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1234),
.A2(n_592),
.B(n_593),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1294),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1228),
.B(n_592),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1212),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1249),
.A2(n_593),
.B(n_447),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1220),
.A2(n_281),
.B(n_447),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1258),
.A2(n_281),
.B(n_447),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1224),
.B(n_450),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1245),
.A2(n_281),
.B(n_447),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1360),
.A2(n_1362),
.B1(n_1297),
.B2(n_1339),
.C(n_1369),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1283),
.A2(n_1286),
.B(n_1315),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1380),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1257),
.B(n_38),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1324),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1260),
.A2(n_333),
.B1(n_281),
.B2(n_447),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1324),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1376),
.A2(n_333),
.B1(n_447),
.B2(n_435),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1426),
.B(n_1295),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1389),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1562),
.A2(n_1308),
.B(n_1309),
.C(n_1331),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1390),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1391),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1539),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1402),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1414),
.A2(n_1376),
.B1(n_1348),
.B2(n_1283),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1566),
.A2(n_1332),
.B1(n_1318),
.B2(n_1285),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1497),
.B(n_1228),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1429),
.A2(n_1332),
.B1(n_1268),
.B2(n_1341),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1562),
.A2(n_1322),
.B1(n_1295),
.B2(n_1321),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1393),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1412),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1388),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1456),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1496),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1388),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1412),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1415),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1514),
.A2(n_1322),
.B1(n_1355),
.B2(n_1296),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1442),
.A2(n_1336),
.B1(n_1243),
.B2(n_1257),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1426),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1489),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1421),
.B(n_1343),
.Y(n_1591)
);

OR2x4_ASAP7_75t_L g1592 ( 
.A(n_1493),
.B(n_1380),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1524),
.A2(n_1243),
.B1(n_1336),
.B2(n_1374),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1427),
.B(n_1380),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1539),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1394),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1458),
.B(n_1257),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1460),
.B(n_1243),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1392),
.A2(n_1365),
.B1(n_1375),
.B2(n_1277),
.C(n_1353),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1531),
.A2(n_1418),
.B1(n_1400),
.B2(n_1473),
.Y(n_1600)
);

CKINVDCx8_ASAP7_75t_R g1601 ( 
.A(n_1422),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1535),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1529),
.B(n_1532),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_SL g1604 ( 
.A(n_1407),
.B(n_356),
.C(n_361),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1516),
.A2(n_1405),
.B1(n_1438),
.B2(n_1449),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1517),
.B(n_1243),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1456),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1418),
.A2(n_1336),
.B1(n_1216),
.B2(n_1356),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1425),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1394),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1473),
.A2(n_1336),
.B1(n_1257),
.B2(n_1335),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1449),
.A2(n_1328),
.B1(n_1313),
.B2(n_1334),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1559),
.A2(n_1336),
.B1(n_1216),
.B2(n_1328),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1535),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1496),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1397),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1399),
.A2(n_1410),
.B(n_1450),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1539),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1490),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1397),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1402),
.A2(n_368),
.B1(n_405),
.B2(n_414),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1458),
.B(n_1324),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1488),
.B(n_449),
.C(n_419),
.Y(n_1623)
);

AND2x2_ASAP7_75t_SL g1624 ( 
.A(n_1467),
.B(n_1336),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1490),
.Y(n_1625)
);

BUFx4f_ASAP7_75t_L g1626 ( 
.A(n_1496),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1509),
.B(n_40),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1496),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1443),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1546),
.A2(n_1352),
.B(n_1350),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1403),
.A2(n_1216),
.B1(n_1352),
.B2(n_333),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1457),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1434),
.A2(n_1307),
.B(n_1216),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1469),
.B(n_1324),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1440),
.B(n_333),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1443),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1473),
.B(n_1337),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1459),
.B(n_1441),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1482),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.C(n_50),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1409),
.A2(n_1216),
.B1(n_45),
.B2(n_50),
.Y(n_1640)
);

AOI222xp33_ASAP7_75t_L g1641 ( 
.A1(n_1433),
.A2(n_41),
.B1(n_51),
.B2(n_54),
.C1(n_55),
.C2(n_59),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1557),
.B(n_51),
.C(n_54),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1529),
.B(n_60),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1455),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1546),
.A2(n_447),
.B(n_104),
.Y(n_1645)
);

CKINVDCx9p33_ASAP7_75t_R g1646 ( 
.A(n_1500),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1456),
.A2(n_447),
.B1(n_63),
.B2(n_65),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1436),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.C(n_68),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1477),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1477),
.B(n_67),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1481),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1452),
.B(n_69),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1497),
.B(n_122),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1489),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1532),
.B(n_69),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1456),
.A2(n_447),
.B1(n_71),
.B2(n_72),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1476),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1457),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1544),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1463),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1484),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1469),
.B(n_75),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1457),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1452),
.B(n_76),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1520),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.C(n_80),
.Y(n_1665)
);

AOI222xp33_ASAP7_75t_L g1666 ( 
.A1(n_1564),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.C1(n_82),
.C2(n_85),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1485),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1443),
.B(n_86),
.Y(n_1668)
);

INVx4_ASAP7_75t_L g1669 ( 
.A(n_1544),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1446),
.A2(n_87),
.B(n_88),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1506),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1486),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1466),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1422),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1480),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1386),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1479),
.B(n_95),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1471),
.B(n_99),
.C(n_100),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1561),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1423),
.A2(n_102),
.B1(n_108),
.B2(n_114),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1386),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1439),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1487),
.B(n_133),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1549),
.A2(n_134),
.B1(n_140),
.B2(n_143),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1489),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1435),
.B(n_146),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1439),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1401),
.A2(n_154),
.B1(n_155),
.B2(n_158),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1489),
.Y(n_1689)
);

INVx4_ASAP7_75t_L g1690 ( 
.A(n_1506),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1545),
.A2(n_162),
.B1(n_164),
.B2(n_174),
.C(n_177),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1497),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1399),
.A2(n_178),
.B(n_179),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1556),
.A2(n_187),
.B(n_193),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1553),
.A2(n_196),
.B1(n_205),
.B2(n_212),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1444),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1556),
.A2(n_220),
.B(n_222),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1444),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1553),
.B(n_1401),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1471),
.Y(n_1700)
);

BUFx10_ASAP7_75t_L g1701 ( 
.A(n_1489),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1542),
.A2(n_1526),
.B1(n_1495),
.B2(n_1398),
.Y(n_1702)
);

CKINVDCx6p67_ASAP7_75t_R g1703 ( 
.A(n_1387),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1521),
.B(n_1396),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1406),
.A2(n_1437),
.B1(n_1417),
.B2(n_1411),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1478),
.A2(n_1534),
.B(n_1528),
.C(n_1501),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1396),
.B(n_1406),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1472),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1411),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1545),
.A2(n_1536),
.B1(n_1468),
.B2(n_1507),
.C(n_1512),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1472),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1417),
.A2(n_1437),
.B1(n_1396),
.B2(n_1475),
.Y(n_1712)
);

BUFx4f_ASAP7_75t_L g1713 ( 
.A(n_1404),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1387),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_R g1715 ( 
.A(n_1467),
.B(n_1408),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1555),
.A2(n_1410),
.B(n_1451),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1555),
.A2(n_1450),
.B(n_1451),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1565),
.A2(n_1563),
.B1(n_1523),
.B2(n_1467),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1541),
.B(n_1543),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1416),
.A2(n_1498),
.B(n_1454),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1523),
.B(n_1561),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1536),
.A2(n_1512),
.B1(n_1507),
.B2(n_1541),
.C(n_1551),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1499),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1522),
.A2(n_1550),
.B(n_1525),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1499),
.Y(n_1726)
);

AOI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1413),
.A2(n_1430),
.B(n_1538),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1474),
.A2(n_1515),
.B1(n_1537),
.B2(n_1548),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1543),
.A2(n_1551),
.B1(n_1540),
.B2(n_1523),
.C(n_1464),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1428),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1408),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1428),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1499),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1510),
.A2(n_1431),
.B1(n_1395),
.B2(n_1503),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1563),
.A2(n_1565),
.B1(n_1491),
.B2(n_1558),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1419),
.B(n_1432),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1385),
.B(n_1465),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1419),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1464),
.A2(n_1502),
.B1(n_1504),
.B2(n_1508),
.C(n_1558),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1432),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1465),
.B(n_1502),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1416),
.A2(n_1454),
.B(n_1461),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1499),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1537),
.A2(n_1548),
.B(n_1510),
.C(n_1504),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1503),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1503),
.B(n_1552),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1385),
.A2(n_1491),
.B1(n_1558),
.B2(n_1511),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1491),
.A2(n_1552),
.B(n_1560),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1430),
.B(n_1511),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1503),
.B(n_1552),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1503),
.B(n_1395),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_SL g1752 ( 
.A(n_1413),
.B(n_1508),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1554),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1465),
.B(n_1527),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1554),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1385),
.B(n_1465),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1383),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1395),
.B(n_1431),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1431),
.B(n_1465),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1383),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1384),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1384),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1453),
.B(n_1548),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1642),
.A2(n_1385),
.B1(n_1538),
.B2(n_1533),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_SL g1765 ( 
.A(n_1619),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1641),
.A2(n_1385),
.B1(n_1533),
.B2(n_1530),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1568),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1580),
.B(n_1453),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1588),
.A2(n_1530),
.B1(n_1527),
.B2(n_1560),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1639),
.A2(n_1505),
.B1(n_1537),
.B2(n_1445),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1660),
.A2(n_1505),
.B1(n_1445),
.B2(n_1424),
.Y(n_1771)
);

NAND4xp25_ASAP7_75t_L g1772 ( 
.A(n_1650),
.B(n_1547),
.C(n_1492),
.D(n_1453),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1635),
.A2(n_1462),
.B(n_1492),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1673),
.A2(n_1404),
.B1(n_1470),
.B2(n_1424),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1585),
.B(n_1453),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1647),
.A2(n_1404),
.B1(n_1470),
.B2(n_1424),
.C(n_1453),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1666),
.A2(n_1470),
.B1(n_1519),
.B2(n_1522),
.Y(n_1777)
);

NAND2x1_ASAP7_75t_L g1778 ( 
.A(n_1671),
.B(n_1690),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1678),
.A2(n_1519),
.B1(n_1462),
.B2(n_1420),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1662),
.B(n_1483),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1657),
.A2(n_1547),
.B1(n_1420),
.B2(n_1461),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1570),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1638),
.B(n_1483),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1643),
.A2(n_1655),
.B1(n_1640),
.B2(n_1665),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1589),
.B(n_1547),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1589),
.B(n_1494),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1635),
.A2(n_1448),
.B(n_1494),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1571),
.Y(n_1788)
);

AOI222xp33_ASAP7_75t_L g1789 ( 
.A1(n_1648),
.A2(n_1702),
.B1(n_1656),
.B2(n_1605),
.C1(n_1627),
.C2(n_1675),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1574),
.A2(n_1547),
.B1(n_1518),
.B2(n_1513),
.C(n_1448),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1668),
.A2(n_1447),
.B(n_1518),
.C(n_1513),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1631),
.A2(n_1447),
.B1(n_1547),
.B2(n_1680),
.Y(n_1792)
);

CKINVDCx11_ASAP7_75t_R g1793 ( 
.A(n_1649),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1604),
.A2(n_1600),
.B(n_1611),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1579),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1575),
.A2(n_1577),
.B1(n_1621),
.B2(n_1609),
.C(n_1586),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1668),
.A2(n_1703),
.B1(n_1643),
.B2(n_1655),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1703),
.A2(n_1597),
.B1(n_1645),
.B2(n_1623),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1591),
.B(n_1662),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1670),
.A2(n_1684),
.B(n_1691),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1652),
.A2(n_1714),
.B1(n_1567),
.B2(n_1582),
.Y(n_1801)
);

OAI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1714),
.A2(n_1567),
.B1(n_1582),
.B2(n_1677),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1597),
.A2(n_1645),
.B1(n_1578),
.B2(n_1756),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1645),
.A2(n_1737),
.B1(n_1756),
.B2(n_1664),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1725),
.A2(n_1717),
.B(n_1716),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1646),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1587),
.A2(n_1593),
.B1(n_1599),
.B2(n_1706),
.C(n_1710),
.Y(n_1807)
);

AOI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1693),
.A2(n_1727),
.B(n_1742),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1644),
.A2(n_1737),
.B1(n_1598),
.B2(n_1594),
.C(n_1606),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1664),
.B(n_1707),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_L g1811 ( 
.A1(n_1699),
.A2(n_1706),
.B(n_1730),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1723),
.A2(n_1695),
.B1(n_1748),
.B2(n_1699),
.C(n_1739),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1736),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1569),
.A2(n_1732),
.B1(n_1634),
.B2(n_1676),
.C(n_1681),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1651),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1633),
.A2(n_1721),
.B(n_1744),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1601),
.A2(n_1704),
.B(n_1755),
.C(n_1753),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1679),
.B(n_1634),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1582),
.A2(n_1624),
.B1(n_1622),
.B2(n_1653),
.Y(n_1819)
);

AOI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1693),
.A2(n_1612),
.B(n_1757),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1682),
.A2(n_1687),
.B(n_1613),
.C(n_1608),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1583),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1622),
.A2(n_1573),
.B1(n_1661),
.B2(n_1667),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1569),
.A2(n_1686),
.B1(n_1688),
.B2(n_1683),
.C(n_1722),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1672),
.A2(n_1747),
.B1(n_1653),
.B2(n_1709),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1603),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1718),
.A2(n_1729),
.B1(n_1712),
.B2(n_1705),
.C(n_1603),
.Y(n_1827)
);

OA21x2_ASAP7_75t_L g1828 ( 
.A1(n_1716),
.A2(n_1717),
.B(n_1731),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1653),
.A2(n_1658),
.B1(n_1632),
.B2(n_1663),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1718),
.A2(n_1759),
.B1(n_1619),
.B2(n_1625),
.C(n_1763),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1683),
.A2(n_1741),
.B1(n_1625),
.B2(n_1754),
.C(n_1734),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1632),
.A2(n_1663),
.B1(n_1658),
.B2(n_1692),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1758),
.A2(n_1728),
.B1(n_1741),
.B2(n_1735),
.C(n_1740),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1659),
.B(n_1576),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_SL g1835 ( 
.A(n_1602),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1637),
.A2(n_1624),
.B(n_1626),
.C(n_1697),
.Y(n_1836)
);

AOI33xp33_ASAP7_75t_L g1837 ( 
.A1(n_1743),
.A2(n_1745),
.A3(n_1762),
.B1(n_1590),
.B2(n_1576),
.B3(n_1719),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1601),
.A2(n_1626),
.B1(n_1649),
.B2(n_1700),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1583),
.Y(n_1839)
);

A2O1A1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1637),
.A2(n_1626),
.B(n_1694),
.C(n_1713),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1632),
.A2(n_1658),
.B1(n_1663),
.B2(n_1692),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1736),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1738),
.A2(n_1740),
.B1(n_1576),
.B2(n_1754),
.C(n_1746),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1738),
.A2(n_1750),
.B1(n_1751),
.B2(n_1731),
.C(n_1700),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1632),
.A2(n_1663),
.B1(n_1658),
.B2(n_1692),
.Y(n_1845)
);

AO21x2_ASAP7_75t_L g1846 ( 
.A1(n_1752),
.A2(n_1761),
.B(n_1760),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1733),
.B(n_1671),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1592),
.A2(n_1713),
.B1(n_1615),
.B2(n_1614),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1630),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1602),
.A2(n_1614),
.B1(n_1674),
.B2(n_1572),
.C(n_1618),
.Y(n_1850)
);

AO21x2_ASAP7_75t_L g1851 ( 
.A1(n_1760),
.A2(n_1761),
.B(n_1630),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1674),
.A2(n_1669),
.B1(n_1592),
.B2(n_1713),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1669),
.A2(n_1671),
.B(n_1690),
.C(n_1595),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1572),
.A2(n_1595),
.B1(n_1618),
.B2(n_1698),
.C(n_1696),
.Y(n_1854)
);

AOI222xp33_ASAP7_75t_L g1855 ( 
.A1(n_1708),
.A2(n_1711),
.B1(n_1581),
.B2(n_1584),
.C1(n_1620),
.C2(n_1616),
.Y(n_1855)
);

AOI222xp33_ASAP7_75t_L g1856 ( 
.A1(n_1711),
.A2(n_1616),
.B1(n_1581),
.B2(n_1620),
.C1(n_1584),
.C2(n_1610),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1572),
.A2(n_1618),
.B1(n_1595),
.B2(n_1610),
.C(n_1596),
.Y(n_1857)
);

NAND3xp33_ASAP7_75t_L g1858 ( 
.A(n_1690),
.B(n_1669),
.C(n_1590),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1628),
.B(n_1685),
.Y(n_1859)
);

AOI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1583),
.A2(n_1628),
.B(n_1726),
.C(n_1724),
.Y(n_1860)
);

OAI21xp33_ASAP7_75t_L g1861 ( 
.A1(n_1654),
.A2(n_1685),
.B(n_1726),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1630),
.A2(n_1583),
.B1(n_1749),
.B2(n_1615),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1749),
.A2(n_1715),
.B1(n_1615),
.B2(n_1726),
.C(n_1689),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1629),
.A2(n_1636),
.B1(n_1654),
.B2(n_1689),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1689),
.B(n_1724),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1720),
.A2(n_1724),
.B1(n_1629),
.B2(n_1636),
.C(n_1715),
.Y(n_1866)
);

OAI33xp33_ASAP7_75t_L g1867 ( 
.A1(n_1720),
.A2(n_1749),
.A3(n_1701),
.B1(n_1636),
.B2(n_1629),
.B3(n_1617),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1701),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1749),
.B(n_1617),
.Y(n_1869)
);

AOI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1701),
.A2(n_1488),
.B(n_1442),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1568),
.Y(n_1871)
);

OAI211xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1641),
.A2(n_1049),
.B(n_960),
.C(n_1036),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1660),
.A2(n_1215),
.B1(n_1009),
.B2(n_1222),
.Y(n_1873)
);

OAI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1641),
.A2(n_748),
.B(n_680),
.C(n_1648),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1574),
.A2(n_891),
.B1(n_661),
.B2(n_1016),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1877)
);

BUFx4f_ASAP7_75t_L g1878 ( 
.A(n_1583),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1642),
.A2(n_680),
.B1(n_801),
.B2(n_867),
.C(n_752),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1642),
.A2(n_680),
.B1(n_801),
.B2(n_867),
.C(n_752),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1568),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1635),
.A2(n_1440),
.B(n_1633),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1884)
);

OAI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1660),
.A2(n_1215),
.B1(n_1009),
.B2(n_1222),
.Y(n_1885)
);

INVxp67_ASAP7_75t_SL g1886 ( 
.A(n_1589),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1567),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1568),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1639),
.A2(n_1029),
.B1(n_1566),
.B2(n_1376),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1638),
.B(n_1426),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1619),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1619),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1574),
.A2(n_891),
.B1(n_661),
.B2(n_1016),
.Y(n_1897)
);

OAI211xp5_ASAP7_75t_L g1898 ( 
.A1(n_1641),
.A2(n_748),
.B(n_680),
.C(n_1648),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1638),
.B(n_1426),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1642),
.A2(n_1009),
.B(n_748),
.Y(n_1900)
);

OAI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1641),
.A2(n_748),
.B(n_680),
.C(n_1648),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1639),
.A2(n_1029),
.B1(n_1566),
.B2(n_1376),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1903)
);

NAND2xp33_ASAP7_75t_R g1904 ( 
.A(n_1607),
.B(n_1047),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1568),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1642),
.A2(n_680),
.B1(n_801),
.B2(n_867),
.C(n_752),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1568),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1714),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1638),
.B(n_1426),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1639),
.A2(n_1029),
.B1(n_1566),
.B2(n_1376),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1638),
.B(n_1426),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1574),
.A2(n_891),
.B1(n_661),
.B2(n_1016),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1641),
.A2(n_1029),
.B(n_1040),
.Y(n_1917)
);

AND2x6_ASAP7_75t_L g1918 ( 
.A(n_1653),
.B(n_1539),
.Y(n_1918)
);

AND2x4_ASAP7_75t_SL g1919 ( 
.A(n_1703),
.B(n_1402),
.Y(n_1919)
);

OAI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1639),
.A2(n_680),
.B1(n_1009),
.B2(n_869),
.C(n_854),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1568),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1635),
.A2(n_1440),
.B(n_1633),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1574),
.A2(n_891),
.B1(n_661),
.B2(n_1016),
.Y(n_1923)
);

O2A1O1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1642),
.A2(n_1029),
.B(n_853),
.C(n_1049),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1925)
);

AOI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1670),
.A2(n_1693),
.B(n_1562),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1642),
.A2(n_1016),
.B1(n_1191),
.B2(n_947),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1780),
.B(n_1869),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1828),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1828),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1818),
.B(n_1768),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1815),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1785),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1775),
.B(n_1846),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1846),
.B(n_1804),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1893),
.B(n_1899),
.Y(n_1936)
);

AO31x2_ASAP7_75t_L g1937 ( 
.A1(n_1816),
.A2(n_1883),
.A3(n_1922),
.B(n_1792),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1851),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1865),
.B(n_1847),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1888),
.B(n_1842),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1851),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1806),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1886),
.Y(n_1943)
);

AO21x2_ASAP7_75t_L g1944 ( 
.A1(n_1808),
.A2(n_1781),
.B(n_1820),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1804),
.B(n_1783),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1767),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1805),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1782),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1910),
.B(n_1914),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1847),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1888),
.B(n_1842),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1920),
.A2(n_1927),
.B1(n_1925),
.B2(n_1875),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1811),
.B(n_1786),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1788),
.B(n_1871),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1881),
.B(n_1889),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1879),
.A2(n_1880),
.B1(n_1907),
.B2(n_1901),
.C(n_1898),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1905),
.Y(n_1957)
);

OAI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1900),
.A2(n_1917),
.B1(n_1874),
.B2(n_1875),
.C(n_1925),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1877),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1908),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1921),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1882),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1814),
.B(n_1795),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1884),
.A2(n_1927),
.B1(n_1887),
.B2(n_1890),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1826),
.B(n_1813),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1896),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1906),
.B(n_1769),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1769),
.B(n_1862),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1862),
.B(n_1823),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1817),
.B(n_1772),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1863),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1830),
.B(n_1837),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1823),
.B(n_1926),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1790),
.B(n_1787),
.Y(n_1976)
);

INVxp67_ASAP7_75t_L g1977 ( 
.A(n_1867),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1918),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1773),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1855),
.Y(n_1980)
);

AOI21xp33_ASAP7_75t_L g1981 ( 
.A1(n_1873),
.A2(n_1885),
.B(n_1789),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1856),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1810),
.B(n_1819),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1799),
.B(n_1809),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1866),
.B(n_1825),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1825),
.B(n_1833),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_R g1987 ( 
.A(n_1904),
.B(n_1793),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1859),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1918),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1834),
.B(n_1802),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1857),
.Y(n_1991)
);

INVx5_ASAP7_75t_L g1992 ( 
.A(n_1918),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1812),
.B(n_1771),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1778),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1859),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1807),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1868),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1854),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1827),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1861),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1771),
.B(n_1770),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1836),
.B(n_1858),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1844),
.B(n_1802),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1864),
.Y(n_2004)
);

BUFx12f_ASAP7_75t_L g2005 ( 
.A(n_1822),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1843),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1884),
.A2(n_1911),
.B1(n_1892),
.B2(n_1890),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1781),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1770),
.B(n_1764),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1764),
.B(n_1766),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1801),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1766),
.B(n_1779),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1801),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1797),
.B(n_1831),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1822),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_SL g2016 ( 
.A1(n_1891),
.A2(n_1912),
.B1(n_1902),
.B2(n_1824),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1791),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1779),
.B(n_1797),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1796),
.B(n_1798),
.Y(n_2019)
);

AOI221xp5_ASAP7_75t_L g2020 ( 
.A1(n_1958),
.A2(n_1911),
.B1(n_1915),
.B2(n_1913),
.C(n_1903),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1928),
.B(n_1909),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1933),
.Y(n_2022)
);

OAI321xp33_ASAP7_75t_L g2023 ( 
.A1(n_1958),
.A2(n_1993),
.A3(n_2019),
.B1(n_1964),
.B2(n_2007),
.C(n_1977),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1987),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1999),
.A2(n_1916),
.B1(n_1876),
.B2(n_1923),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1977),
.A2(n_1887),
.B1(n_1903),
.B2(n_1915),
.C(n_1913),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1942),
.B(n_1850),
.Y(n_2027)
);

OA21x2_ASAP7_75t_L g2028 ( 
.A1(n_1929),
.A2(n_1798),
.B(n_1794),
.Y(n_2028)
);

NAND2x1_ASAP7_75t_L g2029 ( 
.A(n_2002),
.B(n_1895),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1999),
.A2(n_1897),
.B1(n_1885),
.B2(n_1873),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1959),
.B(n_1894),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1932),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1932),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1981),
.A2(n_1800),
.B(n_1840),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1928),
.B(n_1919),
.Y(n_2035)
);

OAI211xp5_ASAP7_75t_SL g2036 ( 
.A1(n_1956),
.A2(n_2016),
.B(n_2017),
.C(n_1981),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1936),
.B(n_1860),
.Y(n_2037)
);

AOI211xp5_ASAP7_75t_L g2038 ( 
.A1(n_1993),
.A2(n_1784),
.B(n_1924),
.C(n_1872),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_2010),
.A2(n_1892),
.B1(n_1784),
.B2(n_1870),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1946),
.Y(n_2040)
);

OAI33xp33_ASAP7_75t_L g2041 ( 
.A1(n_2019),
.A2(n_1838),
.A3(n_1848),
.B1(n_1852),
.B2(n_1774),
.B3(n_1765),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1928),
.B(n_1839),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1929),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1959),
.B(n_1839),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1987),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1936),
.B(n_1853),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_1952),
.A2(n_1821),
.B1(n_1829),
.B2(n_1904),
.C(n_1777),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_1988),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1940),
.B(n_1832),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1942),
.B(n_1996),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2016),
.A2(n_1777),
.B1(n_1878),
.B2(n_1835),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1952),
.A2(n_1878),
.B1(n_1835),
.B2(n_1776),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1959),
.B(n_1839),
.Y(n_2053)
);

AOI222xp33_ASAP7_75t_L g2054 ( 
.A1(n_1964),
.A2(n_1765),
.B1(n_1839),
.B2(n_1841),
.C1(n_1845),
.C2(n_2007),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1946),
.Y(n_2055)
);

AND2x2_ASAP7_75t_SL g2056 ( 
.A(n_2008),
.B(n_1845),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1933),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1956),
.A2(n_1996),
.B1(n_2014),
.B2(n_1993),
.Y(n_2058)
);

OAI211xp5_ASAP7_75t_L g2059 ( 
.A1(n_2008),
.A2(n_1972),
.B(n_2017),
.C(n_1976),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1996),
.A2(n_1972),
.B(n_2003),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2010),
.A2(n_1986),
.B1(n_2012),
.B2(n_2009),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1948),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_1996),
.A2(n_1974),
.B1(n_1986),
.B2(n_2012),
.C(n_1984),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1986),
.A2(n_2012),
.B1(n_2009),
.B2(n_1982),
.Y(n_2064)
);

NAND2xp33_ASAP7_75t_R g2065 ( 
.A(n_2002),
.B(n_1985),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1948),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_SL g2067 ( 
.A1(n_2009),
.A2(n_1985),
.B1(n_2001),
.B2(n_1974),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1957),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1949),
.B(n_1962),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_R g2070 ( 
.A(n_2002),
.B(n_1985),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1962),
.B(n_1967),
.Y(n_2071)
);

NOR2x1_ASAP7_75t_L g2072 ( 
.A(n_2002),
.B(n_1994),
.Y(n_2072)
);

OAI221xp5_ASAP7_75t_SL g2073 ( 
.A1(n_2014),
.A2(n_2003),
.B1(n_2018),
.B2(n_1976),
.C(n_2001),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1978),
.B(n_1989),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1949),
.B(n_1962),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1960),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1940),
.B(n_1951),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1967),
.B(n_1953),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1931),
.B(n_1969),
.Y(n_2079)
);

NAND4xp25_ASAP7_75t_SL g2080 ( 
.A(n_2018),
.B(n_2014),
.C(n_2001),
.D(n_1976),
.Y(n_2080)
);

AOI221xp5_ASAP7_75t_L g2081 ( 
.A1(n_1984),
.A2(n_1998),
.B1(n_1991),
.B2(n_1975),
.C(n_1945),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1940),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_1930),
.A2(n_1947),
.B(n_1938),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1960),
.Y(n_2084)
);

NOR2x1_ASAP7_75t_R g2085 ( 
.A(n_2002),
.B(n_2005),
.Y(n_2085)
);

NOR4xp25_ASAP7_75t_SL g2086 ( 
.A(n_1943),
.B(n_2011),
.C(n_2013),
.D(n_1991),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1988),
.Y(n_2087)
);

AO21x2_ASAP7_75t_L g2088 ( 
.A1(n_1944),
.A2(n_1941),
.B(n_1938),
.Y(n_2088)
);

OA21x2_ASAP7_75t_L g2089 ( 
.A1(n_1930),
.A2(n_1947),
.B(n_1941),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_1951),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2018),
.A2(n_1975),
.B(n_1979),
.C(n_2000),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_1988),
.Y(n_2092)
);

OAI21xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1975),
.A2(n_1969),
.B(n_1953),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1961),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1998),
.A2(n_2006),
.B1(n_1983),
.B2(n_1970),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_SL g2096 ( 
.A1(n_1970),
.A2(n_1968),
.B1(n_1966),
.B2(n_1935),
.Y(n_2096)
);

OAI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_1973),
.A2(n_1963),
.B1(n_2006),
.B2(n_1935),
.C(n_2013),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_1973),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2069),
.B(n_1945),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2079),
.B(n_1939),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_2072),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2082),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2026),
.A2(n_2020),
.B1(n_2080),
.B2(n_2063),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2022),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2079),
.B(n_1939),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2083),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2081),
.A2(n_1970),
.B1(n_1980),
.B2(n_1982),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2071),
.B(n_2048),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2058),
.A2(n_1980),
.B1(n_1968),
.B2(n_1966),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2057),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2083),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2092),
.B(n_2069),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2077),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2075),
.B(n_1939),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2074),
.B(n_1992),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2074),
.B(n_1992),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2083),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2075),
.B(n_1939),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2077),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2089),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2044),
.B(n_1931),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2065),
.Y(n_2122)
);

OAI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2059),
.A2(n_1935),
.B(n_1979),
.Y(n_2123)
);

NOR2x1_ASAP7_75t_L g2124 ( 
.A(n_2046),
.B(n_2029),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2074),
.B(n_1992),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2090),
.B(n_1945),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2044),
.B(n_1931),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2032),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2098),
.B(n_1954),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2033),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2050),
.B(n_1943),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2050),
.B(n_1943),
.Y(n_2132)
);

NAND2xp67_ASAP7_75t_L g2133 ( 
.A(n_2034),
.B(n_1954),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2053),
.B(n_1969),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2087),
.B(n_1992),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2024),
.B(n_1950),
.Y(n_2136)
);

NAND2xp67_ASAP7_75t_L g2137 ( 
.A(n_2021),
.B(n_1955),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2078),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2091),
.B(n_1955),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2049),
.B(n_1965),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2040),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2049),
.B(n_1965),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2093),
.B(n_1955),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2089),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2031),
.B(n_1937),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2042),
.B(n_2035),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2024),
.B(n_1950),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_2035),
.B(n_1992),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2055),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2037),
.B(n_2000),
.Y(n_2150)
);

INVxp67_ASAP7_75t_SL g2151 ( 
.A(n_2065),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2042),
.B(n_1992),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_2062),
.B(n_1937),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2045),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2096),
.B(n_1995),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_2060),
.B(n_2045),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2027),
.B(n_1950),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2061),
.B(n_2027),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_2066),
.B(n_1937),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_2043),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2068),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_2036),
.B(n_1997),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2076),
.B(n_2084),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2094),
.B(n_1934),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2023),
.B(n_1997),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2099),
.B(n_2095),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2150),
.B(n_2067),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2161),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2115),
.B(n_1978),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2128),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2100),
.B(n_1937),
.Y(n_2171)
);

OAI32xp33_ASAP7_75t_L g2172 ( 
.A1(n_2123),
.A2(n_2070),
.A3(n_2097),
.B1(n_2051),
.B2(n_2039),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2162),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2139),
.B(n_2123),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2126),
.B(n_1937),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_2165),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2106),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2128),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_2154),
.B(n_2156),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_2115),
.B(n_1978),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2130),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2130),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2103),
.A2(n_2070),
.B1(n_2030),
.B2(n_2038),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2141),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2141),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_2115),
.B(n_1978),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2139),
.B(n_1937),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2126),
.B(n_1937),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_2124),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2124),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2100),
.B(n_1937),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2149),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2149),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_2115),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_2116),
.Y(n_2195)
);

OAI21xp33_ASAP7_75t_L g2196 ( 
.A1(n_2133),
.A2(n_2073),
.B(n_1990),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2113),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_2108),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2140),
.B(n_1990),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2113),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2129),
.B(n_2112),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2104),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2119),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2119),
.Y(n_2204)
);

AOI311xp33_ASAP7_75t_L g2205 ( 
.A1(n_2104),
.A2(n_2047),
.A3(n_1961),
.B(n_2052),
.C(n_2011),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2154),
.B(n_2085),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_2116),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2105),
.B(n_2004),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2163),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2106),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2140),
.B(n_1990),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2106),
.Y(n_2212)
);

INVxp67_ASAP7_75t_SL g2213 ( 
.A(n_2122),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2111),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2111),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2105),
.B(n_2004),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2108),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2142),
.B(n_2028),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2134),
.B(n_2004),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2102),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2111),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2166),
.B(n_2133),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2170),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2177),
.Y(n_2224)
);

NAND2x1p5_ASAP7_75t_L g2225 ( 
.A(n_2189),
.B(n_1992),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2198),
.B(n_2114),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2176),
.A2(n_2028),
.B1(n_2158),
.B2(n_2151),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2170),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2178),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2177),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2198),
.B(n_2114),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2217),
.B(n_2118),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_2202),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2209),
.B(n_2143),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2178),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2210),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2169),
.B(n_2116),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_2169),
.B(n_2116),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2209),
.B(n_2143),
.Y(n_2239)
);

INVx3_ASAP7_75t_SL g2240 ( 
.A(n_2190),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_R g2241 ( 
.A(n_2206),
.B(n_2136),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2181),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2179),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2181),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_2169),
.Y(n_2245)
);

NOR2x1_ASAP7_75t_R g2246 ( 
.A(n_2189),
.B(n_2148),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2217),
.B(n_2118),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2199),
.B(n_2142),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2182),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2168),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2168),
.Y(n_2251)
);

NAND4xp25_ASAP7_75t_L g2252 ( 
.A(n_2205),
.B(n_2174),
.C(n_2183),
.D(n_2187),
.Y(n_2252)
);

NAND4xp25_ASAP7_75t_L g2253 ( 
.A(n_2172),
.B(n_2145),
.C(n_2025),
.D(n_2107),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2199),
.B(n_2153),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2211),
.B(n_2153),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2194),
.B(n_2112),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2194),
.B(n_2121),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2211),
.B(n_2159),
.Y(n_2258)
);

NAND4xp25_ASAP7_75t_L g2259 ( 
.A(n_2172),
.B(n_2145),
.C(n_2159),
.D(n_2109),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2197),
.B(n_2129),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2182),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2173),
.B(n_2110),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2194),
.B(n_2121),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2184),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2210),
.Y(n_2265)
);

INVx1_ASAP7_75t_SL g2266 ( 
.A(n_2167),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_2213),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2184),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2185),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2195),
.B(n_2127),
.Y(n_2270)
);

NAND2xp33_ASAP7_75t_SL g2271 ( 
.A(n_2190),
.B(n_2157),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_2169),
.B(n_2125),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2195),
.B(n_2127),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2212),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2185),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2195),
.B(n_2157),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2212),
.Y(n_2277)
);

OAI21xp33_ASAP7_75t_L g2278 ( 
.A1(n_2252),
.A2(n_2188),
.B(n_2175),
.Y(n_2278)
);

INVxp67_ASAP7_75t_SL g2279 ( 
.A(n_2267),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2267),
.B(n_2196),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2250),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2243),
.B(n_2101),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2251),
.Y(n_2283)
);

NAND2x1_ASAP7_75t_L g2284 ( 
.A(n_2237),
.B(n_2207),
.Y(n_2284)
);

AOI211xp5_ASAP7_75t_L g2285 ( 
.A1(n_2252),
.A2(n_2175),
.B(n_2171),
.C(n_2191),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2241),
.B(n_2101),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2233),
.B(n_2219),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2223),
.Y(n_2288)
);

AOI221xp5_ASAP7_75t_L g2289 ( 
.A1(n_2259),
.A2(n_2064),
.B1(n_2171),
.B2(n_2191),
.C(n_2218),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2223),
.Y(n_2290)
);

AOI221xp5_ASAP7_75t_L g2291 ( 
.A1(n_2259),
.A2(n_2218),
.B1(n_2214),
.B2(n_2215),
.C(n_2221),
.Y(n_2291)
);

OAI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_2253),
.A2(n_2028),
.B1(n_1963),
.B2(n_2131),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2248),
.B(n_2234),
.Y(n_2293)
);

XOR2x2_ASAP7_75t_L g2294 ( 
.A(n_2266),
.B(n_2155),
.Y(n_2294)
);

OAI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2253),
.A2(n_2221),
.B1(n_2214),
.B2(n_2215),
.C(n_2200),
.Y(n_2295)
);

OAI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2227),
.A2(n_2222),
.B1(n_2239),
.B2(n_2271),
.C(n_2254),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2262),
.A2(n_2041),
.B1(n_2054),
.B2(n_1971),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2248),
.B(n_2219),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2228),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_2240),
.Y(n_2300)
);

INVx1_ASAP7_75t_SL g2301 ( 
.A(n_2240),
.Y(n_2301)
);

XOR2x2_ASAP7_75t_L g2302 ( 
.A(n_2225),
.B(n_2155),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2226),
.B(n_2207),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2256),
.B(n_2208),
.Y(n_2304)
);

OAI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2240),
.A2(n_2132),
.B1(n_2254),
.B2(n_2255),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2224),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2224),
.A2(n_1968),
.B1(n_1966),
.B2(n_2056),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2256),
.B(n_2208),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2224),
.Y(n_2309)
);

AOI322xp5_ASAP7_75t_L g2310 ( 
.A1(n_2230),
.A2(n_2134),
.A3(n_2164),
.B1(n_2201),
.B2(n_1983),
.C1(n_2056),
.C2(n_1971),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2226),
.B(n_2216),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2228),
.Y(n_2312)
);

OAI211xp5_ASAP7_75t_L g2313 ( 
.A1(n_2245),
.A2(n_2207),
.B(n_2086),
.C(n_2220),
.Y(n_2313)
);

AOI222xp33_ASAP7_75t_L g2314 ( 
.A1(n_2230),
.A2(n_1971),
.B1(n_2144),
.B2(n_2120),
.C1(n_2117),
.C2(n_1983),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2245),
.A2(n_2180),
.B1(n_2186),
.B2(n_2216),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2229),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2260),
.B(n_2197),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_SL g2318 ( 
.A1(n_2245),
.A2(n_2147),
.B(n_2135),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2229),
.Y(n_2319)
);

NAND2x1_ASAP7_75t_L g2320 ( 
.A(n_2303),
.B(n_2245),
.Y(n_2320)
);

AOI222xp33_ASAP7_75t_L g2321 ( 
.A1(n_2292),
.A2(n_2277),
.B1(n_2274),
.B2(n_2265),
.C1(n_2236),
.C2(n_2230),
.Y(n_2321)
);

OAI21xp33_ASAP7_75t_L g2322 ( 
.A1(n_2278),
.A2(n_2276),
.B(n_2257),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2288),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2300),
.B(n_2276),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2293),
.B(n_2260),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2290),
.Y(n_2326)
);

AOI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2292),
.A2(n_2277),
.B(n_2236),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2279),
.B(n_2237),
.Y(n_2328)
);

INVxp67_ASAP7_75t_L g2329 ( 
.A(n_2286),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2306),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2299),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2312),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2316),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2319),
.Y(n_2334)
);

OAI322xp33_ASAP7_75t_L g2335 ( 
.A1(n_2280),
.A2(n_2255),
.A3(n_2258),
.B1(n_2264),
.B2(n_2269),
.C1(n_2268),
.C2(n_2242),
.Y(n_2335)
);

NAND2x1p5_ASAP7_75t_L g2336 ( 
.A(n_2301),
.B(n_2237),
.Y(n_2336)
);

AOI322xp5_ASAP7_75t_L g2337 ( 
.A1(n_2291),
.A2(n_2289),
.A3(n_2297),
.B1(n_2307),
.B2(n_2279),
.C1(n_2305),
.C2(n_2285),
.Y(n_2337)
);

O2A1O1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_2282),
.A2(n_2249),
.B(n_2275),
.C(n_2235),
.Y(n_2338)
);

INVx2_ASAP7_75t_SL g2339 ( 
.A(n_2284),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2306),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2311),
.B(n_2237),
.Y(n_2341)
);

INVxp67_ASAP7_75t_L g2342 ( 
.A(n_2286),
.Y(n_2342)
);

AOI221xp5_ASAP7_75t_L g2343 ( 
.A1(n_2295),
.A2(n_2277),
.B1(n_2265),
.B2(n_2236),
.C(n_2274),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2281),
.B(n_2231),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2297),
.A2(n_2265),
.B1(n_2274),
.B2(n_2258),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2294),
.A2(n_1944),
.B1(n_2117),
.B2(n_2120),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2304),
.B(n_2238),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2296),
.A2(n_2238),
.B1(n_2272),
.B2(n_2231),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2308),
.B(n_2238),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2282),
.B(n_2246),
.Y(n_2350)
);

INVx1_ASAP7_75t_SL g2351 ( 
.A(n_2328),
.Y(n_2351)
);

XNOR2x1_ASAP7_75t_L g2352 ( 
.A(n_2345),
.B(n_2302),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2325),
.Y(n_2353)
);

OAI21xp33_ASAP7_75t_L g2354 ( 
.A1(n_2337),
.A2(n_2287),
.B(n_2313),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2324),
.B(n_2283),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2324),
.B(n_2328),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2330),
.Y(n_2357)
);

NOR2x1_ASAP7_75t_L g2358 ( 
.A(n_2328),
.B(n_2305),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2336),
.B(n_2238),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2336),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2330),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2329),
.B(n_2310),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2340),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2340),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2347),
.B(n_2272),
.Y(n_2365)
);

XNOR2x2_ASAP7_75t_L g2366 ( 
.A(n_2350),
.B(n_2317),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2342),
.B(n_2350),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2341),
.B(n_2298),
.Y(n_2368)
);

INVx5_ASAP7_75t_L g2369 ( 
.A(n_2339),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2341),
.B(n_2347),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2323),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2326),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2331),
.Y(n_2373)
);

AOI221x1_ASAP7_75t_L g2374 ( 
.A1(n_2327),
.A2(n_2309),
.B1(n_2315),
.B2(n_2235),
.C(n_2242),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2367),
.B(n_2349),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2359),
.Y(n_2376)
);

AOI211xp5_ASAP7_75t_L g2377 ( 
.A1(n_2354),
.A2(n_2335),
.B(n_2348),
.C(n_2338),
.Y(n_2377)
);

NOR3xp33_ASAP7_75t_L g2378 ( 
.A(n_2360),
.B(n_2343),
.C(n_2322),
.Y(n_2378)
);

INVx1_ASAP7_75t_SL g2379 ( 
.A(n_2351),
.Y(n_2379)
);

AOI322xp5_ASAP7_75t_L g2380 ( 
.A1(n_2362),
.A2(n_2346),
.A3(n_2321),
.B1(n_2332),
.B2(n_2334),
.C1(n_2333),
.C2(n_2309),
.Y(n_2380)
);

O2A1O1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2366),
.A2(n_2346),
.B(n_2344),
.C(n_2339),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2353),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_SL g2383 ( 
.A(n_2366),
.Y(n_2383)
);

OAI221xp5_ASAP7_75t_L g2384 ( 
.A1(n_2352),
.A2(n_2358),
.B1(n_2361),
.B2(n_2364),
.C(n_2357),
.Y(n_2384)
);

XNOR2xp5_ASAP7_75t_L g2385 ( 
.A(n_2352),
.B(n_2349),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2374),
.B(n_2244),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2370),
.A2(n_2320),
.B(n_2246),
.Y(n_2387)
);

NOR4xp25_ASAP7_75t_SL g2388 ( 
.A(n_2363),
.B(n_2318),
.C(n_2275),
.D(n_2244),
.Y(n_2388)
);

NOR3xp33_ASAP7_75t_L g2389 ( 
.A(n_2356),
.B(n_2269),
.C(n_2249),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_SL g2390 ( 
.A(n_2381),
.B(n_2359),
.C(n_2355),
.Y(n_2390)
);

NAND4xp25_ASAP7_75t_L g2391 ( 
.A(n_2375),
.B(n_2368),
.C(n_2365),
.D(n_2371),
.Y(n_2391)
);

OAI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2383),
.A2(n_2377),
.B1(n_2384),
.B2(n_2385),
.Y(n_2392)
);

OAI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2380),
.A2(n_2365),
.B(n_2369),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2379),
.B(n_2372),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2378),
.A2(n_2386),
.B1(n_2376),
.B2(n_2382),
.Y(n_2395)
);

AOI322xp5_ASAP7_75t_L g2396 ( 
.A1(n_2386),
.A2(n_2389),
.A3(n_2373),
.B1(n_2388),
.B2(n_2314),
.C1(n_2369),
.C2(n_2120),
.Y(n_2396)
);

NOR2x1_ASAP7_75t_L g2397 ( 
.A(n_2387),
.B(n_2369),
.Y(n_2397)
);

AOI222xp33_ASAP7_75t_L g2398 ( 
.A1(n_2384),
.A2(n_2369),
.B1(n_2117),
.B2(n_2144),
.C1(n_2261),
.C2(n_2268),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2375),
.B(n_2369),
.Y(n_2399)
);

OAI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2384),
.A2(n_2225),
.B1(n_2261),
.B2(n_2264),
.Y(n_2400)
);

AOI211xp5_ASAP7_75t_SL g2401 ( 
.A1(n_2384),
.A2(n_2272),
.B(n_2270),
.C(n_2263),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2392),
.B(n_2232),
.Y(n_2402)
);

O2A1O1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_2390),
.A2(n_2225),
.B(n_2220),
.C(n_2270),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2394),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2396),
.B(n_2232),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2399),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2395),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2393),
.B(n_2272),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2407),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2406),
.B(n_2391),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_L g2411 ( 
.A(n_2404),
.B(n_2400),
.C(n_2397),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2405),
.A2(n_2401),
.B1(n_2204),
.B2(n_2203),
.Y(n_2412)
);

NAND4xp25_ASAP7_75t_L g2413 ( 
.A(n_2402),
.B(n_2398),
.C(n_2273),
.D(n_2263),
.Y(n_2413)
);

NOR4xp25_ASAP7_75t_L g2414 ( 
.A(n_2403),
.B(n_2273),
.C(n_2257),
.D(n_2204),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2408),
.B(n_2247),
.Y(n_2415)
);

NAND4xp25_ASAP7_75t_L g2416 ( 
.A(n_2406),
.B(n_2247),
.C(n_2180),
.D(n_2186),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2409),
.Y(n_2417)
);

NOR2x1_ASAP7_75t_L g2418 ( 
.A(n_2410),
.B(n_2413),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_SL g2419 ( 
.A(n_2411),
.B(n_2414),
.C(n_2412),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2415),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2416),
.Y(n_2421)
);

HB1xp67_ASAP7_75t_L g2422 ( 
.A(n_2415),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2417),
.A2(n_2144),
.B1(n_2088),
.B2(n_1944),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2422),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2420),
.B(n_2200),
.Y(n_2425)
);

NAND2x1p5_ASAP7_75t_L g2426 ( 
.A(n_2418),
.B(n_2180),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2424),
.Y(n_2427)
);

OAI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2427),
.A2(n_2424),
.B1(n_2426),
.B2(n_2421),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_2428),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2428),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2430),
.Y(n_2431)
);

AOI31xp33_ASAP7_75t_L g2432 ( 
.A1(n_2429),
.A2(n_2419),
.A3(n_2425),
.B(n_2423),
.Y(n_2432)
);

AOI222xp33_ASAP7_75t_L g2433 ( 
.A1(n_2431),
.A2(n_2203),
.B1(n_2193),
.B2(n_2192),
.C1(n_2110),
.C2(n_2180),
.Y(n_2433)
);

OAI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2432),
.A2(n_2193),
.B1(n_2192),
.B2(n_2102),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2434),
.A2(n_2186),
.B1(n_2088),
.B2(n_2160),
.Y(n_2435)
);

OAI221xp5_ASAP7_75t_R g2436 ( 
.A1(n_2435),
.A2(n_2433),
.B1(n_2138),
.B2(n_2137),
.C(n_2146),
.Y(n_2436)
);

AOI211xp5_ASAP7_75t_L g2437 ( 
.A1(n_2436),
.A2(n_2125),
.B(n_2015),
.C(n_2152),
.Y(n_2437)
);


endmodule