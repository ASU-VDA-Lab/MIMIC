module fake_netlist_6_755_n_182 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_182);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_182;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVxp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVxp33_ASAP7_75t_SL g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_4),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_32),
.B(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_45),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_53),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_44),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_32),
.B1(n_35),
.B2(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_51),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_39),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_75),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_72),
.B(n_73),
.Y(n_93)
);

AO31x2_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_71),
.A3(n_64),
.B(n_63),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_71),
.B(n_64),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_65),
.C(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx4_ASAP7_75t_SL g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_56),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_77),
.B(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_81),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_87),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_87),
.Y(n_107)
);

O2A1O1Ixp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_76),
.B(n_82),
.C(n_81),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_35),
.Y(n_110)
);

AOI222xp33_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_83),
.B1(n_69),
.B2(n_106),
.C1(n_38),
.C2(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_96),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OR2x6_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_99),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_121),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OAI31xp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_111),
.A3(n_103),
.B(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI33xp33_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_57),
.A3(n_54),
.B1(n_58),
.B2(n_80),
.B3(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AOI222xp33_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_98),
.B1(n_57),
.B2(n_56),
.C1(n_99),
.C2(n_58),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_115),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_99),
.B(n_115),
.Y(n_142)
);

AOI211xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_128),
.B(n_126),
.C(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_138),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_126),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_127),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_127),
.B(n_108),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_129),
.B(n_133),
.C(n_132),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_132),
.B(n_100),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_113),
.Y(n_150)
);

OAI221xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_80),
.B1(n_104),
.B2(n_113),
.C(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_110),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_142),
.B(n_151),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_98),
.B1(n_56),
.B2(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_8),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_9),
.B(n_10),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_10),
.Y(n_167)
);

OAI322xp33_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_155),
.A3(n_159),
.B1(n_157),
.B2(n_160),
.C1(n_11),
.C2(n_12),
.Y(n_168)
);

OAI211xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_159),
.B(n_11),
.C(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_158),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_158),
.B1(n_98),
.B2(n_99),
.C(n_82),
.Y(n_171)
);

OAI211xp5_ASAP7_75t_SL g172 ( 
.A1(n_162),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_166),
.B(n_167),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_166),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_95),
.B1(n_20),
.B2(n_26),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_19),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_95),
.B1(n_56),
.B2(n_94),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_174),
.B(n_176),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_178),
.B1(n_177),
.B2(n_179),
.Y(n_182)
);


endmodule