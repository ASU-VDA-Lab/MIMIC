module real_jpeg_19843_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_0),
.A2(n_7),
.B1(n_21),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_54),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_53),
.B(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_7),
.B(n_10),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_2),
.A2(n_18),
.B1(n_24),
.B2(n_81),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_35),
.B1(n_48),
.B2(n_90),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_18),
.B1(n_24),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_7),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_25),
.B1(n_52),
.B2(n_54),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_4),
.A2(n_7),
.B1(n_21),
.B2(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_7),
.B1(n_21),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_18),
.B1(n_24),
.B2(n_38),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_10),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_8),
.B1(n_21),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_18),
.Y(n_19)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_68),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_44),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_28),
.C(n_34),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_16),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_17),
.A2(n_20),
.B1(n_26),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_17),
.A2(n_20),
.B1(n_23),
.B2(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g51 ( 
.A1(n_18),
.A2(n_33),
.A3(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_94),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_24),
.B(n_81),
.C(n_82),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_24),
.B(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_31),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_32),
.B(n_54),
.C(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_54),
.Y(n_59)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B(n_39),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_35),
.A2(n_41),
.B1(n_75),
.B2(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_42),
.B(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_81),
.Y(n_94)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_97),
.B(n_102),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_86),
.B(n_96),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_95),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);


endmodule