module real_aes_2582_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_769;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_0), .B(n_112), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_1), .A2(n_125), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_2), .B(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_3), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g119 ( .A(n_4), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_5), .B(n_134), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_6), .B(n_121), .Y(n_494) );
INVx1_ASAP7_75t_L g470 ( .A(n_7), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_8), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_9), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_10), .B(n_132), .Y(n_197) );
INVx2_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
AOI221x1_ASAP7_75t_L g141 ( .A1(n_12), .A2(n_24), .B1(n_112), .B2(n_125), .C(n_142), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_13), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_14), .B(n_112), .Y(n_193) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_15), .A2(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g502 ( .A(n_16), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_17), .B(n_139), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_18), .B(n_134), .Y(n_185) );
AO21x1_ASAP7_75t_L g111 ( .A1(n_19), .A2(n_112), .B(n_120), .Y(n_111) );
INVx1_ASAP7_75t_L g435 ( .A(n_20), .Y(n_435) );
INVx1_ASAP7_75t_L g500 ( .A(n_21), .Y(n_500) );
INVx1_ASAP7_75t_SL g551 ( .A(n_22), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_23), .B(n_113), .Y(n_514) );
NAND2x1_ASAP7_75t_L g152 ( .A(n_25), .B(n_134), .Y(n_152) );
AOI33xp33_ASAP7_75t_L g538 ( .A1(n_26), .A2(n_52), .A3(n_451), .B1(n_458), .B2(n_539), .B3(n_540), .Y(n_538) );
NAND2x1_ASAP7_75t_L g211 ( .A(n_27), .B(n_132), .Y(n_211) );
INVx1_ASAP7_75t_L g478 ( .A(n_28), .Y(n_478) );
OR2x2_ASAP7_75t_L g122 ( .A(n_29), .B(n_85), .Y(n_122) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_29), .A2(n_85), .B(n_123), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_30), .B(n_449), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_31), .B(n_132), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_32), .B(n_134), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_33), .B(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_34), .A2(n_125), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g797 ( .A(n_35), .Y(n_797) );
AND2x2_ASAP7_75t_L g118 ( .A(n_36), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g126 ( .A(n_36), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g457 ( .A(n_36), .Y(n_457) );
OR2x6_ASAP7_75t_L g433 ( .A(n_37), .B(n_434), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_38), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_39), .B(n_112), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_40), .B(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_41), .A2(n_121), .B1(n_157), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_42), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_43), .B(n_113), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_44), .Y(n_189) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_45), .A2(n_100), .B1(n_787), .B2(n_788), .C1(n_794), .C2(n_797), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_45), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_46), .B(n_132), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_47), .B(n_191), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_48), .B(n_113), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_49), .A2(n_125), .B(n_210), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_50), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_51), .B(n_132), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_53), .B(n_113), .Y(n_463) );
INVx1_ASAP7_75t_L g115 ( .A(n_54), .Y(n_115) );
INVx1_ASAP7_75t_L g129 ( .A(n_54), .Y(n_129) );
AND2x2_ASAP7_75t_L g464 ( .A(n_55), .B(n_139), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_56), .A2(n_74), .B1(n_449), .B2(n_455), .C(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_57), .B(n_449), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_58), .B(n_134), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_59), .B(n_157), .Y(n_487) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_60), .A2(n_455), .B(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_61), .A2(n_125), .B(n_151), .Y(n_150) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_62), .A2(n_99), .B1(n_798), .B2(n_809), .C1(n_823), .C2(n_827), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_62), .A2(n_103), .B1(n_812), .B2(n_813), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_62), .Y(n_813) );
INVx1_ASAP7_75t_L g497 ( .A(n_63), .Y(n_497) );
AO21x1_ASAP7_75t_L g124 ( .A1(n_64), .A2(n_125), .B(n_130), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_65), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_66), .B(n_112), .Y(n_202) );
INVx1_ASAP7_75t_L g461 ( .A(n_67), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_68), .B(n_112), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_69), .A2(n_455), .B(n_460), .Y(n_454) );
AND2x2_ASAP7_75t_L g169 ( .A(n_70), .B(n_140), .Y(n_169) );
INVx1_ASAP7_75t_L g117 ( .A(n_71), .Y(n_117) );
INVx1_ASAP7_75t_L g127 ( .A(n_71), .Y(n_127) );
AND2x2_ASAP7_75t_L g215 ( .A(n_72), .B(n_156), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_73), .B(n_449), .Y(n_541) );
AND2x2_ASAP7_75t_L g553 ( .A(n_75), .B(n_156), .Y(n_553) );
INVx1_ASAP7_75t_L g498 ( .A(n_76), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_77), .A2(n_455), .B(n_550), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_78), .A2(n_455), .B(n_513), .C(n_517), .Y(n_512) );
INVx1_ASAP7_75t_L g436 ( .A(n_79), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_80), .B(n_112), .Y(n_187) );
AND2x2_ASAP7_75t_L g200 ( .A(n_81), .B(n_156), .Y(n_200) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_82), .B(n_156), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_83), .A2(n_455), .B1(n_536), .B2(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g120 ( .A(n_84), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g159 ( .A(n_86), .B(n_156), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_87), .B(n_132), .Y(n_186) );
INVx1_ASAP7_75t_L g524 ( .A(n_88), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_89), .B(n_134), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_90), .B(n_132), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_91), .A2(n_125), .B(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g542 ( .A(n_92), .B(n_156), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_93), .B(n_134), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_94), .A2(n_476), .B(n_477), .C(n_480), .Y(n_475) );
BUFx2_ASAP7_75t_L g806 ( .A(n_95), .Y(n_806) );
BUFx2_ASAP7_75t_SL g831 ( .A(n_95), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_96), .A2(n_125), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_97), .B(n_113), .Y(n_525) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_428), .B1(n_437), .B2(n_783), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_103), .A2(n_790), .B1(n_792), .B2(n_793), .Y(n_789) );
INVx1_ASAP7_75t_L g812 ( .A(n_103), .Y(n_812) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_327), .Y(n_103) );
NOR3xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_264), .C(n_287), .Y(n_104) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_216), .C(n_233), .Y(n_105) );
OAI31xp33_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_146), .A3(n_170), .B(n_177), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_107), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_138), .Y(n_108) );
AND2x4_ASAP7_75t_L g219 ( .A(n_109), .B(n_138), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_109), .B(n_161), .Y(n_248) );
AND2x4_ASAP7_75t_L g250 ( .A(n_109), .B(n_244), .Y(n_250) );
AND2x2_ASAP7_75t_L g381 ( .A(n_109), .B(n_174), .Y(n_381) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g226 ( .A(n_110), .Y(n_226) );
OAI21x1_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_124), .B(n_136), .Y(n_110) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_118), .Y(n_112) );
INVx1_ASAP7_75t_L g479 ( .A(n_113), .Y(n_479) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
AND2x6_ASAP7_75t_L g132 ( .A(n_114), .B(n_127), .Y(n_132) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g134 ( .A(n_116), .B(n_129), .Y(n_134) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx5_ASAP7_75t_L g135 ( .A(n_118), .Y(n_135) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_118), .Y(n_480) );
AND2x2_ASAP7_75t_L g128 ( .A(n_119), .B(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_119), .Y(n_452) );
INVx1_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_121), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_SL g181 ( .A(n_121), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_121), .A2(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_121), .B(n_135), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_121), .A2(n_522), .B(n_526), .Y(n_521) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_122), .B(n_123), .Y(n_140) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
BUFx3_ASAP7_75t_L g453 ( .A(n_126), .Y(n_453) );
INVx2_ASAP7_75t_L g459 ( .A(n_127), .Y(n_459) );
AND2x4_ASAP7_75t_L g455 ( .A(n_128), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g451 ( .A(n_129), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_135), .Y(n_130) );
INVxp67_ASAP7_75t_L g501 ( .A(n_132), .Y(n_501) );
INVxp67_ASAP7_75t_L g503 ( .A(n_134), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_135), .A2(n_143), .B(n_144), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_135), .A2(n_152), .B(n_153), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_135), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_135), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_135), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_135), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_135), .A2(n_211), .B(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_135), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g469 ( .A1(n_135), .A2(n_462), .B(n_470), .C(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_135), .A2(n_514), .B(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_135), .A2(n_462), .B(n_524), .C(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g536 ( .A(n_135), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_135), .A2(n_462), .B(n_551), .C(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g160 ( .A(n_138), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_138), .B(n_225), .Y(n_317) );
AND2x2_ASAP7_75t_L g323 ( .A(n_138), .B(n_162), .Y(n_323) );
AND2x2_ASAP7_75t_L g412 ( .A(n_138), .B(n_413), .Y(n_412) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_141), .B(n_145), .Y(n_138) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_139), .A2(n_141), .B(n_145), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_139), .A2(n_202), .B(n_203), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_139), .Y(n_214) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_SL g394 ( .A(n_146), .Y(n_394) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_160), .Y(n_146) );
BUFx2_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
AND2x2_ASAP7_75t_L g257 ( .A(n_147), .B(n_161), .Y(n_257) );
AND2x2_ASAP7_75t_L g306 ( .A(n_147), .B(n_162), .Y(n_306) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g263 ( .A(n_148), .B(n_162), .Y(n_263) );
INVxp67_ASAP7_75t_L g275 ( .A(n_148), .Y(n_275) );
BUFx3_ASAP7_75t_L g320 ( .A(n_148), .Y(n_320) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_155), .B(n_159), .Y(n_148) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_149), .A2(n_155), .B(n_159), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_155), .A2(n_163), .B(n_169), .Y(n_162) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_155), .A2(n_163), .B(n_169), .Y(n_176) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_155), .A2(n_447), .B(n_464), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_155), .A2(n_156), .B1(n_475), .B2(n_481), .Y(n_474) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_155), .A2(n_447), .B(n_464), .Y(n_603) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_157), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
OAI31xp33_ASAP7_75t_L g216 ( .A1(n_160), .A2(n_217), .A3(n_222), .B(n_227), .Y(n_216) );
AND2x2_ASAP7_75t_L g224 ( .A(n_161), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g243 ( .A(n_162), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_164), .B(n_168), .Y(n_163) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_170), .A2(n_292), .A3(n_321), .B1(n_326), .B2(n_418), .C1(n_421), .C2(n_422), .Y(n_417) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_171), .B(n_263), .Y(n_268) );
NAND2x1_ASAP7_75t_L g305 ( .A(n_171), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g349 ( .A(n_171), .B(n_253), .Y(n_349) );
INVx1_ASAP7_75t_SL g363 ( .A(n_171), .Y(n_363) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g244 ( .A(n_172), .Y(n_244) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_172), .Y(n_387) );
AND2x2_ASAP7_75t_L g316 ( .A(n_173), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_173), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_SL g173 ( .A(n_174), .B(n_175), .Y(n_173) );
BUFx2_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
INVx1_ASAP7_75t_L g413 ( .A(n_174), .Y(n_413) );
OR2x2_ASAP7_75t_L g280 ( .A(n_175), .B(n_225), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_175), .B(n_250), .Y(n_314) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x4_ASAP7_75t_L g253 ( .A(n_176), .B(n_225), .Y(n_253) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_198), .Y(n_177) );
INVxp67_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g309 ( .A(n_179), .Y(n_309) );
OR2x2_ASAP7_75t_L g336 ( .A(n_179), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_190), .Y(n_179) );
NOR2x1_ASAP7_75t_SL g230 ( .A(n_180), .B(n_199), .Y(n_230) );
AND2x2_ASAP7_75t_L g237 ( .A(n_180), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g409 ( .A(n_180), .B(n_271), .Y(n_409) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_181), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
OR2x2_ASAP7_75t_L g231 ( .A(n_190), .B(n_232), .Y(n_231) );
BUFx3_ASAP7_75t_L g240 ( .A(n_190), .Y(n_240) );
INVx2_ASAP7_75t_L g271 ( .A(n_190), .Y(n_271) );
INVx1_ASAP7_75t_L g312 ( .A(n_190), .Y(n_312) );
AND2x2_ASAP7_75t_L g343 ( .A(n_190), .B(n_199), .Y(n_343) );
AND2x2_ASAP7_75t_L g374 ( .A(n_190), .B(n_301), .Y(n_374) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_191), .A2(n_468), .B(n_472), .Y(n_467) );
INVx2_ASAP7_75t_SL g517 ( .A(n_191), .Y(n_517) );
AND2x2_ASAP7_75t_L g270 ( .A(n_198), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_198), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_198), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_198), .B(n_240), .Y(n_378) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_207), .Y(n_198) );
INVx5_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_199), .B(n_232), .Y(n_310) );
BUFx2_ASAP7_75t_L g370 ( .A(n_199), .Y(n_370) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx4_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
AND2x2_ASAP7_75t_L g355 ( .A(n_207), .B(n_238), .Y(n_355) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_215), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_213), .Y(n_208) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_214), .A2(n_547), .B(n_553), .Y(n_546) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_218), .A2(n_345), .B1(n_348), .B2(n_350), .C(n_351), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g366 ( .A(n_219), .B(n_257), .Y(n_366) );
INVx1_ASAP7_75t_SL g392 ( .A(n_219), .Y(n_392) );
AND2x2_ASAP7_75t_L g377 ( .A(n_220), .B(n_349), .Y(n_377) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_221), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AND2x2_ASAP7_75t_L g246 ( .A(n_223), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g252 ( .A(n_223), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
AND2x2_ASAP7_75t_L g334 ( .A(n_224), .B(n_262), .Y(n_334) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
OR2x2_ASAP7_75t_L g423 ( .A(n_231), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g239 ( .A(n_232), .Y(n_239) );
AND2x4_ASAP7_75t_L g295 ( .A(n_232), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_232), .B(n_300), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_232), .B(n_238), .Y(n_337) );
AND2x2_ASAP7_75t_L g397 ( .A(n_232), .B(n_300), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_241), .B1(n_254), .B2(n_256), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_234), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND3x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .C(n_240), .Y(n_236) );
AND2x4_ASAP7_75t_L g254 ( .A(n_237), .B(n_255), .Y(n_254) );
INVx4_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_238), .B(n_295), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_239), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
AOI322xp5_ASAP7_75t_L g404 ( .A1(n_240), .A2(n_369), .A3(n_405), .B1(n_407), .B2(n_410), .C1(n_414), .C2(n_415), .Y(n_404) );
NAND4xp25_ASAP7_75t_SL g241 ( .A(n_242), .B(n_245), .C(n_249), .D(n_251), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_243), .B(n_259), .Y(n_371) );
BUFx2_ASAP7_75t_L g262 ( .A(n_244), .Y(n_262) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g386 ( .A(n_247), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g400 ( .A(n_248), .B(n_275), .Y(n_400) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g266 ( .A(n_250), .B(n_267), .Y(n_266) );
OAI211xp5_ASAP7_75t_L g318 ( .A1(n_250), .A2(n_319), .B(n_321), .C(n_324), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_250), .B(n_257), .Y(n_376) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_252), .A2(n_334), .B1(n_335), .B2(n_338), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_253), .A2(n_289), .B1(n_293), .B2(n_297), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_253), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_253), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_253), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g420 ( .A(n_253), .Y(n_420) );
INVx1_ASAP7_75t_L g359 ( .A(n_254), .Y(n_359) );
OAI21xp33_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_258), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g267 ( .A(n_257), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_257), .B(n_262), .Y(n_416) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g352 ( .A(n_259), .B(n_263), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_261), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g419 ( .A(n_262), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g393 ( .A(n_263), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B(n_269), .C(n_272), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI22xp33_ASAP7_75t_SL g379 ( .A1(n_267), .A2(n_298), .B1(n_345), .B2(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_271), .B(n_294), .Y(n_302) );
OR2x2_ASAP7_75t_L g331 ( .A(n_271), .B(n_332), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_277), .B(n_281), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g292 ( .A(n_275), .Y(n_292) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI211xp5_ASAP7_75t_SL g330 ( .A1(n_278), .A2(n_331), .B(n_333), .C(n_341), .Y(n_330) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp67_ASAP7_75t_SL g364 ( .A(n_283), .B(n_310), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_283), .Y(n_367) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_285), .B(n_294), .Y(n_424) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
INVx2_ASAP7_75t_L g301 ( .A(n_286), .Y(n_301) );
NAND4xp25_ASAP7_75t_L g287 ( .A(n_288), .B(n_303), .C(n_315), .D(n_318), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_291), .A2(n_423), .B1(n_425), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x4_ASAP7_75t_L g390 ( .A(n_294), .B(n_320), .Y(n_390) );
AND2x2_ASAP7_75t_L g311 ( .A(n_295), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
AND2x2_ASAP7_75t_L g342 ( .A(n_295), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
INVx1_ASAP7_75t_L g346 ( .A(n_302), .Y(n_346) );
AOI32xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .A3(n_310), .B1(n_311), .B2(n_313), .Y(n_303) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_352), .B(n_353), .Y(n_351) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_307), .A2(n_384), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_383) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g368 ( .A(n_309), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g326 ( .A(n_310), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_311), .A2(n_349), .B1(n_399), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g325 ( .A(n_312), .Y(n_325) );
AND2x2_ASAP7_75t_L g403 ( .A(n_312), .B(n_356), .Y(n_403) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_319), .B(n_371), .Y(n_406) );
INVx1_ASAP7_75t_L g425 ( .A(n_319), .Y(n_425) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g327 ( .A(n_328), .B(n_382), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_372), .Y(n_328) );
NOR3xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_344), .C(n_357), .Y(n_329) );
INVx1_ASAP7_75t_L g347 ( .A(n_332), .Y(n_347) );
INVx1_ASAP7_75t_SL g358 ( .A(n_334), .Y(n_358) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g340 ( .A(n_337), .Y(n_340) );
INVx2_ASAP7_75t_L g350 ( .A(n_338), .Y(n_350) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x4_ASAP7_75t_L g396 ( .A(n_339), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g414 ( .A(n_343), .B(n_397), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_354), .A2(n_366), .A3(n_367), .B1(n_368), .B2(n_371), .Y(n_365) );
NOR2xp33_ASAP7_75t_SL g384 ( .A(n_354), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g385 ( .A(n_356), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_359), .B(n_360), .C(n_365), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g421 ( .A(n_369), .B(n_409), .Y(n_421) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_370), .B(n_409), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B1(n_377), .B2(n_378), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g380 ( .A(n_381), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_398), .C(n_404), .D(n_417), .Y(n_382) );
INVxp33_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_394), .C(n_395), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
CKINVDCx11_ASAP7_75t_R g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_SL g793 ( .A(n_429), .Y(n_793) );
INVx3_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
AND2x6_ASAP7_75t_SL g431 ( .A(n_432), .B(n_433), .Y(n_431) );
OR2x6_ASAP7_75t_SL g785 ( .A(n_432), .B(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g796 ( .A(n_432), .B(n_433), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_432), .B(n_786), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_433), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_L g792 ( .A(n_437), .Y(n_792) );
NAND4xp75_ASAP7_75t_L g437 ( .A(n_438), .B(n_655), .C(n_700), .D(n_769), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_615), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_571), .C(n_596), .Y(n_440) );
OAI222xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_489), .B1(n_527), .B2(n_543), .C1(n_558), .C2(n_565), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_465), .Y(n_443) );
AND2x2_ASAP7_75t_L g780 ( .A(n_444), .B(n_594), .Y(n_780) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_446), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_446), .B(n_473), .Y(n_570) );
INVx3_ASAP7_75t_L g585 ( .A(n_446), .Y(n_585) );
AND2x2_ASAP7_75t_L g718 ( .A(n_446), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_454), .Y(n_447) );
INVx1_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g509 ( .A(n_450), .Y(n_509) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
OR2x6_ASAP7_75t_L g462 ( .A(n_451), .B(n_459), .Y(n_462) );
INVxp33_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
INVx1_ASAP7_75t_L g510 ( .A(n_453), .Y(n_510) );
INVxp67_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
NOR2x1p5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g540 ( .A(n_458), .Y(n_540) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_462), .A2(n_479), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
AND2x2_ASAP7_75t_L g648 ( .A(n_465), .B(n_601), .Y(n_648) );
AND2x2_ASAP7_75t_L g650 ( .A(n_465), .B(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g685 ( .A(n_465), .Y(n_685) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_473), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g568 ( .A(n_467), .Y(n_568) );
INVx1_ASAP7_75t_L g587 ( .A(n_467), .Y(n_587) );
AND2x4_ASAP7_75t_L g594 ( .A(n_467), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_467), .B(n_533), .Y(n_610) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_467), .Y(n_719) );
INVx1_ASAP7_75t_L g729 ( .A(n_467), .Y(n_729) );
INVx1_ASAP7_75t_L g530 ( .A(n_473), .Y(n_530) );
INVx2_ASAP7_75t_L g582 ( .A(n_473), .Y(n_582) );
INVx1_ASAP7_75t_L g663 ( .A(n_473), .Y(n_663) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_491), .B(n_518), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_491), .B(n_545), .Y(n_638) );
INVx2_ASAP7_75t_L g659 ( .A(n_491), .Y(n_659) );
AND2x2_ASAP7_75t_L g667 ( .A(n_491), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_505), .Y(n_491) );
AND2x4_ASAP7_75t_L g557 ( .A(n_492), .B(n_506), .Y(n_557) );
INVx1_ASAP7_75t_L g564 ( .A(n_492), .Y(n_564) );
AND2x2_ASAP7_75t_L g740 ( .A(n_492), .B(n_546), .Y(n_740) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g578 ( .A(n_493), .B(n_506), .Y(n_578) );
INVx2_ASAP7_75t_L g614 ( .A(n_493), .Y(n_614) );
AND2x2_ASAP7_75t_L g693 ( .A(n_493), .B(n_546), .Y(n_693) );
NOR2x1_ASAP7_75t_SL g736 ( .A(n_493), .B(n_519), .Y(n_736) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_499), .B(n_504), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g590 ( .A(n_506), .B(n_519), .Y(n_590) );
INVx1_ASAP7_75t_L g606 ( .A(n_506), .Y(n_606) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_506), .Y(n_714) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_512), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .C(n_511), .Y(n_508) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_517), .A2(n_534), .B(n_542), .Y(n_533) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_517), .A2(n_534), .B(n_542), .Y(n_583) );
AND2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_578), .Y(n_577) );
OR2x6_ASAP7_75t_L g658 ( .A(n_518), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g696 ( .A(n_518), .B(n_693), .Y(n_696) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_519), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g625 ( .A(n_519), .Y(n_625) );
OR2x2_ASAP7_75t_L g631 ( .A(n_519), .B(n_546), .Y(n_631) );
AND2x4_ASAP7_75t_L g645 ( .A(n_519), .B(n_606), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_519), .B(n_614), .Y(n_646) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g690 ( .A(n_530), .B(n_609), .Y(n_690) );
BUFx2_ASAP7_75t_L g742 ( .A(n_530), .Y(n_742) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g773 ( .A(n_532), .B(n_685), .Y(n_773) );
INVx2_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_541), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_554), .Y(n_543) );
AND2x2_ASAP7_75t_L g589 ( .A(n_544), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_SL g574 ( .A(n_545), .B(n_564), .Y(n_574) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g562 ( .A(n_546), .Y(n_562) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_546), .Y(n_668) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_546), .Y(n_735) );
INVx1_ASAP7_75t_L g775 ( .A(n_546), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
BUFx2_ASAP7_75t_L g689 ( .A(n_554), .Y(n_689) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x4_ASAP7_75t_L g605 ( .A(n_555), .B(n_606), .Y(n_605) );
NOR2xp67_ASAP7_75t_SL g637 ( .A(n_555), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g710 ( .A(n_555), .B(n_693), .Y(n_710) );
AND2x4_ASAP7_75t_SL g713 ( .A(n_555), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g762 ( .A(n_555), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
INVx4_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g624 ( .A(n_557), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_557), .B(n_622), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_557), .B(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_557), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g707 ( .A(n_561), .B(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g623 ( .A(n_562), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
AND2x2_ASAP7_75t_L g741 ( .A(n_566), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g749 ( .A(n_566), .B(n_678), .Y(n_749) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g618 ( .A(n_567), .B(n_603), .Y(n_618) );
AND2x4_ASAP7_75t_L g651 ( .A(n_567), .B(n_585), .Y(n_651) );
INVx1_ASAP7_75t_L g768 ( .A(n_567), .Y(n_768) );
AND2x2_ASAP7_75t_L g654 ( .A(n_569), .B(n_594), .Y(n_654) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g675 ( .A(n_570), .B(n_610), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_579), .B1(n_588), .B2(n_591), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_577), .Y(n_572) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_573), .A2(n_642), .B1(n_750), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_574), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g643 ( .A(n_574), .B(n_575), .Y(n_643) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_574), .B(n_645), .Y(n_673) );
AOI211xp5_ASAP7_75t_SL g761 ( .A1(n_574), .A2(n_762), .B(n_764), .C(n_765), .Y(n_761) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_575), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_575), .B(n_621), .Y(n_747) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
INVx2_ASAP7_75t_L g708 ( .A(n_578), .Y(n_708) );
AND2x2_ASAP7_75t_L g782 ( .A(n_578), .B(n_775), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_579), .A2(n_731), .B(n_737), .Y(n_730) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g717 ( .A(n_581), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g727 ( .A(n_581), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g634 ( .A(n_582), .B(n_587), .Y(n_634) );
NOR2xp67_ASAP7_75t_L g636 ( .A(n_582), .B(n_603), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_582), .B(n_603), .Y(n_678) );
INVx2_ASAP7_75t_L g595 ( .A(n_583), .Y(n_595) );
AND2x4_ASAP7_75t_L g601 ( .A(n_583), .B(n_602), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx3_ASAP7_75t_L g593 ( .A(n_585), .Y(n_593) );
INVx3_ASAP7_75t_L g599 ( .A(n_586), .Y(n_599) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_590), .A2(n_696), .B(n_772), .Y(n_776) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g608 ( .A(n_593), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_593), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_593), .B(n_668), .Y(n_683) );
OR2x2_ASAP7_75t_L g698 ( .A(n_593), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g705 ( .A(n_593), .B(n_609), .Y(n_705) );
AND2x2_ASAP7_75t_L g661 ( .A(n_594), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g677 ( .A(n_594), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g694 ( .A(n_594), .B(n_663), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_604), .B1(n_607), .B2(n_611), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_599), .B(n_600), .Y(n_671) );
NOR2xp67_ASAP7_75t_SL g709 ( .A(n_599), .B(n_617), .Y(n_709) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_603), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g612 ( .A(n_605), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g676 ( .A(n_605), .B(n_622), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_605), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g779 ( .A(n_613), .B(n_645), .Y(n_779) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_614), .B(n_725), .Y(n_724) );
NOR2xp67_ASAP7_75t_SL g615 ( .A(n_616), .B(n_639), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B(n_626), .C(n_635), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_617), .A2(n_670), .B(n_680), .C(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g759 ( .A(n_618), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g670 ( .A(n_622), .B(n_646), .Y(n_670) );
AND2x2_ASAP7_75t_L g757 ( .A(n_622), .B(n_736), .Y(n_757) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g725 ( .A(n_625), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_632), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_629), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g699 ( .A(n_634), .Y(n_699) );
NAND2xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_647), .B1(n_649), .B2(n_652), .C(n_653), .Y(n_639) );
NOR4xp25_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .C(n_644), .D(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g758 ( .A(n_645), .B(n_721), .Y(n_758) );
INVx2_ASAP7_75t_L g764 ( .A(n_645), .Y(n_764) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_648), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g751 ( .A(n_651), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND4xp75_ASAP7_75t_L g656 ( .A(n_657), .B(n_679), .C(n_686), .D(n_695), .Y(n_656) );
OA211x2_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_664), .C(n_672), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_658), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g752 ( .A(n_662), .Y(n_752) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g760 ( .A(n_663), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_671), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx2_ASAP7_75t_L g721 ( .A(n_668), .Y(n_721) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_672) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_676), .A2(n_727), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g755 ( .A(n_677), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_678), .B(n_768), .Y(n_767) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVxp67_ASAP7_75t_L g753 ( .A(n_689), .Y(n_753) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_693), .B(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_694), .A2(n_757), .B1(n_779), .B2(n_780), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND3x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_743), .C(n_756), .Y(n_701) );
NOR3x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_715), .C(n_730), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_711), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_709), .B2(n_710), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_720), .B1(n_722), .B2(n_726), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g774 ( .A(n_724), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g763 ( .A(n_740), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g771 ( .A1(n_741), .A2(n_772), .B(n_774), .Y(n_771) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_754), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B1(n_750), .B2(n_753), .Y(n_744) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
O2A1O1Ixp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_759), .C(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR2x1_ASAP7_75t_SL g769 ( .A(n_770), .B(n_777), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_776), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_778), .B(n_781), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_784), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx4f_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_807), .Y(n_800) );
INVxp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_803), .B(n_806), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_SL g826 ( .A(n_804), .B(n_806), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_804), .A2(n_829), .B(n_832), .Y(n_828) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_R g816 ( .A(n_808), .Y(n_816) );
BUFx3_ASAP7_75t_L g821 ( .A(n_808), .Y(n_821) );
BUFx2_ASAP7_75t_L g833 ( .A(n_808), .Y(n_833) );
INVxp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_814), .B(n_817), .Y(n_810) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_SL g817 ( .A(n_818), .B(n_822), .Y(n_817) );
INVx1_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
BUFx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
CKINVDCx11_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
CKINVDCx8_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
endmodule