module fake_jpeg_15497_n_216 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_25),
.Y(n_65)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_52),
.B1(n_59),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_0),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.C(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_93),
.B1(n_58),
.B2(n_57),
.Y(n_109)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_18),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_21),
.B1(n_24),
.B2(n_20),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_17),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_21),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_50),
.C(n_32),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_27),
.B1(n_32),
.B2(n_4),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_35),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_111),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_61),
.B(n_31),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_48),
.C(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_58),
.B1(n_57),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_81),
.B1(n_75),
.B2(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_56),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_57),
.B1(n_48),
.B2(n_60),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_32),
.B1(n_27),
.B2(n_56),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_79),
.B(n_69),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_77),
.A3(n_71),
.B1(n_82),
.B2(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_126),
.B(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_85),
.B1(n_94),
.B2(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_74),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_92),
.C(n_96),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_130),
.C(n_106),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_133),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_91),
.C(n_68),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_8),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_106),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_115),
.B(n_107),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_152),
.B(n_156),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_100),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_158),
.C(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_159),
.B1(n_105),
.B2(n_56),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_97),
.B(n_108),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_119),
.A3(n_15),
.B1(n_16),
.B2(n_14),
.C1(n_11),
.C2(n_7),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_22),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_125),
.A3(n_128),
.B1(n_131),
.B2(n_127),
.C1(n_130),
.C2(n_121),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_138),
.B(n_140),
.C(n_132),
.D(n_56),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_111),
.Y(n_160)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_123),
.CI(n_137),
.CON(n_163),
.SN(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_173),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.C(n_175),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_3),
.B(n_5),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_5),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_158),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_6),
.C(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_161),
.C(n_146),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_143),
.B1(n_150),
.B2(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_143),
.C(n_148),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_172),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_196),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_169),
.B1(n_167),
.B2(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_146),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_165),
.B(n_179),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_203),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_189),
.B(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_177),
.B(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_171),
.B1(n_163),
.B2(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_194),
.B1(n_163),
.B2(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_145),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_145),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_186),
.C(n_198),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_210),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_148),
.B(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_209),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_214),
.Y(n_216)
);


endmodule