module fake_jpeg_293_n_446 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_446);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_10),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_56),
.B(n_73),
.Y(n_125)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_58),
.Y(n_169)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_61),
.B(n_62),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_66),
.B(n_68),
.Y(n_166)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_69),
.B(n_74),
.Y(n_170)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_13),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_76),
.B(n_81),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_78),
.Y(n_157)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_12),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_30),
.B(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_82),
.B(n_3),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_88),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_22),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_96),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_94),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_19),
.B(n_2),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_104),
.Y(n_156)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

CKINVDCx9p33_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_43),
.C(n_45),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_118),
.B(n_124),
.C(n_122),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_173),
.Y(n_200)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g216 ( 
.A(n_121),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_45),
.C(n_51),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_59),
.B(n_53),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_41),
.B1(n_53),
.B2(n_47),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_168),
.Y(n_211)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_71),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_143),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_47),
.B(n_49),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_109),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_67),
.A2(n_49),
.B1(n_28),
.B2(n_48),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_72),
.A2(n_51),
.B1(n_48),
.B2(n_101),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_75),
.A2(n_95),
.B1(n_93),
.B2(n_110),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_152),
.A2(n_154),
.B1(n_123),
.B2(n_186),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_135),
.C(n_134),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_28),
.B1(n_32),
.B2(n_5),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_167),
.A2(n_127),
.B1(n_141),
.B2(n_158),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_60),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_174),
.A2(n_189),
.B1(n_194),
.B2(n_175),
.Y(n_254)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_174),
.B1(n_194),
.B2(n_158),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_115),
.B(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_10),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_58),
.A2(n_9),
.B1(n_10),
.B2(n_77),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_85),
.B(n_9),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_139),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_90),
.A2(n_10),
.B1(n_108),
.B2(n_109),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_195),
.B(n_208),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_98),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_196),
.B(n_199),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_153),
.B(n_105),
.Y(n_199)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_203),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_209),
.Y(n_288)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_107),
.B1(n_79),
.B2(n_91),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_214),
.A2(n_255),
.B1(n_205),
.B2(n_238),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_215),
.B(n_226),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_125),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_131),
.B(n_83),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_132),
.B(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_221),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_147),
.A2(n_152),
.B1(n_189),
.B2(n_142),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_220),
.A2(n_223),
.B1(n_203),
.B2(n_204),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_133),
.Y(n_221)
);

HAxp5_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_146),
.CON(n_222),
.SN(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_222),
.A2(n_254),
.B(n_211),
.C(n_223),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_225),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_136),
.B(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_144),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_231),
.Y(n_280)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_145),
.B(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_138),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_126),
.B(n_151),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_236),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_234),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_119),
.A2(n_184),
.B(n_161),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_247),
.B(n_209),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_184),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_150),
.A2(n_191),
.B1(n_165),
.B2(n_163),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_123),
.B(n_119),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_251),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_141),
.A2(n_162),
.B1(n_169),
.B2(n_155),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_245),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_162),
.B(n_155),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_169),
.A2(n_155),
.B1(n_160),
.B2(n_122),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_259),
.B1(n_207),
.B2(n_235),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_160),
.B(n_163),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_154),
.B(n_191),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_165),
.B(n_140),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_204),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_180),
.A2(n_166),
.B(n_170),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_200),
.B(n_222),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_185),
.A2(n_187),
.B1(n_116),
.B2(n_94),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_182),
.B(n_166),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_208),
.A3(n_258),
.B1(n_218),
.B2(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_216),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_167),
.A2(n_71),
.B1(n_65),
.B2(n_78),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_269),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_195),
.A2(n_244),
.B(n_242),
.C(n_203),
.D(n_252),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_270),
.A2(n_290),
.B(n_295),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_272),
.A2(n_281),
.B1(n_298),
.B2(n_265),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_251),
.B1(n_214),
.B2(n_211),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_274),
.A2(n_307),
.B1(n_306),
.B2(n_301),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_301),
.B1(n_265),
.B2(n_295),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_215),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_297),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_227),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_211),
.A2(n_206),
.B(n_257),
.C(n_213),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_281),
.B(n_270),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_202),
.B(n_211),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_246),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_237),
.C(n_254),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_238),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_240),
.A2(n_254),
.B1(n_209),
.B2(n_230),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_216),
.B(n_210),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_302),
.A2(n_281),
.B(n_307),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_205),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_197),
.Y(n_324)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_328),
.B1(n_273),
.B2(n_267),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_317),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g348 ( 
.A1(n_315),
.A2(n_331),
.B(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_264),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_318),
.A2(n_333),
.B(n_342),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_320),
.C(n_326),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_201),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_227),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_334),
.Y(n_352)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_274),
.A2(n_197),
.B1(n_201),
.B2(n_279),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_325),
.A2(n_332),
.B1(n_288),
.B2(n_305),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_263),
.B(n_201),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_SL g327 ( 
.A(n_290),
.B(n_201),
.C(n_299),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_327),
.B(n_288),
.CI(n_303),
.CON(n_347),
.SN(n_347)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_336),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_286),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_302),
.B1(n_281),
.B2(n_268),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_294),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_280),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_300),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_341),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_285),
.B(n_260),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_266),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_313),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_260),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_296),
.A2(n_266),
.B(n_276),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_349),
.B1(n_357),
.B2(n_336),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_353),
.B(n_358),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_314),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_313),
.B(n_267),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_350),
.B(n_359),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_273),
.B1(n_292),
.B2(n_277),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_262),
.B1(n_278),
.B2(n_277),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_285),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_365),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_262),
.B(n_278),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_363),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_319),
.A2(n_308),
.A3(n_333),
.B1(n_309),
.B2(n_332),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_309),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_366),
.B(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_322),
.B(n_317),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_345),
.A2(n_318),
.B1(n_326),
.B2(n_339),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_373),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_352),
.B(n_362),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_377),
.Y(n_395)
);

AOI221x1_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_314),
.B1(n_327),
.B2(n_325),
.C(n_317),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_343),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_384),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_320),
.C(n_312),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_364),
.C(n_351),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_340),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_386),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_331),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_366),
.B(n_342),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_388),
.B(n_390),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_346),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_391),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_321),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_329),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_363),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_344),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_406),
.C(n_407),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_356),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_400),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_356),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_380),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_387),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_376),
.C(n_374),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_347),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_330),
.C(n_347),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_386),
.C(n_381),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_418),
.Y(n_425)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_406),
.A2(n_378),
.B(n_391),
.C(n_371),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_410),
.B(n_411),
.Y(n_427)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_385),
.C(n_377),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_400),
.C(n_399),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_403),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_372),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_420),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_387),
.B(n_370),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_396),
.A2(n_375),
.B1(n_392),
.B2(n_373),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_421),
.A2(n_349),
.B1(n_396),
.B2(n_358),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_421),
.A2(n_396),
.B1(n_405),
.B2(n_402),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_424),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_410),
.B1(n_415),
.B2(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_416),
.C(n_412),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_420),
.A2(n_365),
.B1(n_384),
.B2(n_353),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_425),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_432),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_425),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_435),
.B(n_436),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_427),
.A2(n_412),
.B1(n_347),
.B2(n_390),
.Y(n_436)
);

AOI322xp5_ASAP7_75t_L g437 ( 
.A1(n_427),
.A2(n_414),
.A3(n_408),
.B1(n_368),
.B2(n_355),
.C1(n_361),
.C2(n_360),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_422),
.C(n_430),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_436),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_416),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_442),
.C(n_443),
.Y(n_444)
);

NOR4xp25_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_422),
.C(n_434),
.D(n_433),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_435),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_424),
.Y(n_446)
);


endmodule