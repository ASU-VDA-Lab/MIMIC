module fake_jpeg_22235_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_28),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_19),
.B1(n_23),
.B2(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_12),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_25),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_21),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_46),
.CON(n_69),
.SN(n_69)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_64),
.B1(n_46),
.B2(n_42),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_20),
.B(n_2),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_39),
.B(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_56),
.B1(n_41),
.B2(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_54),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_49),
.C(n_41),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_52),
.Y(n_78)
);

NOR4xp25_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_74),
.C(n_66),
.D(n_65),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_81),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_56),
.B1(n_53),
.B2(n_50),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_84),
.B1(n_73),
.B2(n_76),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_73),
.B(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_62),
.B1(n_60),
.B2(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_78),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_77),
.Y(n_97)
);

AOI21x1_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_91),
.B(n_98),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_90),
.C(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule