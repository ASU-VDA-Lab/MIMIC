module fake_jpeg_10570_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_38),
.Y(n_40)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_22),
.B1(n_21),
.B2(n_29),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_46),
.B1(n_53),
.B2(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_14),
.B1(n_27),
.B2(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_55),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_38),
.B1(n_36),
.B2(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_24),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_0),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_64),
.B(n_66),
.Y(n_88)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_34),
.B1(n_28),
.B2(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_70),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_38),
.B1(n_14),
.B2(n_16),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_73),
.B1(n_45),
.B2(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_32),
.B1(n_30),
.B2(n_18),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_42),
.C(n_40),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_45),
.B(n_1),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_84),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_7),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_7),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_60),
.B1(n_49),
.B2(n_4),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_45),
.B1(n_30),
.B2(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_30),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_91),
.C(n_0),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_0),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_57),
.B(n_74),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_97),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_103),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_61),
.B(n_62),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_59),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_75),
.C(n_84),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_70),
.A3(n_68),
.B1(n_69),
.B2(n_59),
.C1(n_64),
.C2(n_13),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_59),
.B(n_68),
.C(n_60),
.D(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.C(n_102),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_91),
.B1(n_80),
.B2(n_81),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_123),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_81),
.B1(n_87),
.B2(n_82),
.Y(n_117)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_124),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_79),
.B1(n_3),
.B2(n_5),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_130),
.C(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_109),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_135),
.B(n_121),
.C(n_115),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_99),
.B(n_107),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_105),
.C(n_99),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_122),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_144),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_118),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_100),
.C(n_119),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_114),
.C(n_2),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_126),
.CI(n_134),
.CON(n_146),
.SN(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_144),
.C(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_147),
.B1(n_143),
.B2(n_151),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_137),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_6),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_156),
.C(n_6),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_155),
.A2(n_142),
.B(n_114),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_149),
.CI(n_147),
.CON(n_160),
.SN(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule