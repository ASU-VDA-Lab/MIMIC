module fake_ariane_1898_n_1868 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1868);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1868;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_29),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_67),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_80),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

BUFx8_ASAP7_75t_SL g181 ( 
.A(n_106),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_138),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_98),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_59),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_4),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_50),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_77),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_17),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_8),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_37),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_40),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_45),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_99),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_72),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_109),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_7),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_102),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_55),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_40),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_160),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_103),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_48),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_18),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_108),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_129),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_121),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_52),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_7),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_131),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_59),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_82),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_97),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_125),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_17),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_91),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_81),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_89),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_94),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_100),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_85),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_21),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_150),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_87),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_92),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_47),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_162),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_38),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_52),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_151),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_30),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_157),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_42),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_28),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_21),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_167),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_134),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_79),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_155),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_137),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_170),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_38),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_139),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_78),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_116),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_23),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_127),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_73),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_28),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_133),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_0),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_50),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_154),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_30),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_5),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_55),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_9),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_153),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_45),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_136),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_57),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_62),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_158),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_27),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_88),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_145),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_27),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_58),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_143),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_48),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_10),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_70),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_174),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_181),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_228),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_187),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_236),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_254),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_187),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_190),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_331),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_180),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_184),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_189),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_192),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_192),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_218),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_202),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_202),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_205),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_241),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_205),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_326),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_263),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_209),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_209),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_214),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_214),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_227),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_263),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_204),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_253),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_230),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_336),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_230),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_220),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_298),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_233),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_176),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_204),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_231),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_270),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_182),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_191),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_245),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_251),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_289),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_193),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_290),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_231),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_324),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_325),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_196),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_232),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_198),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_232),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_206),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_240),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_291),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_291),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_179),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_250),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_250),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_179),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_275),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_275),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_207),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_208),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_304),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_210),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_212),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_264),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_296),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_298),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_215),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_296),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_341),
.B(n_293),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_188),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_343),
.B(n_298),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_355),
.A2(n_262),
.B(n_255),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_255),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_388),
.B(n_259),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_360),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_352),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_374),
.B(n_385),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_374),
.B(n_262),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_361),
.A2(n_282),
.B(n_271),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_361),
.B(n_293),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_363),
.B(n_366),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_370),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_371),
.B(n_334),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_373),
.B(n_377),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_408),
.A2(n_269),
.B1(n_277),
.B2(n_337),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_388),
.B(n_296),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_365),
.B(n_172),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_353),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_411),
.A2(n_274),
.B1(n_261),
.B2(n_260),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_334),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_409),
.B(n_301),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_410),
.A2(n_282),
.B(n_271),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_SL g495 ( 
.A(n_412),
.B(n_334),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_285),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g498 ( 
.A1(n_364),
.A2(n_305),
.B(n_285),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_358),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_439),
.Y(n_500)
);

INVx11_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_439),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_447),
.B(n_416),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_439),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_439),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_446),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_447),
.A2(n_476),
.B1(n_346),
.B2(n_406),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_439),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_454),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_454),
.B(n_334),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_447),
.B(n_416),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_385),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_454),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_437),
.B(n_417),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_447),
.B(n_384),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_475),
.B(n_389),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_379),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_365),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_452),
.B(n_342),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_454),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_446),
.B(n_390),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_305),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_454),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_394),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

AND3x2_ASAP7_75t_L g537 ( 
.A(n_446),
.B(n_405),
.C(n_415),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_437),
.B(n_399),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_459),
.B(n_401),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_480),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_469),
.B(n_403),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_498),
.A2(n_413),
.B1(n_301),
.B2(n_307),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_469),
.B(n_414),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_458),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_430),
.B(n_418),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_469),
.B(n_422),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_496),
.B(n_431),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_458),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_476),
.A2(n_248),
.B1(n_224),
.B2(n_280),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_458),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_350),
.C(n_175),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_498),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_430),
.B(n_347),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_474),
.B(n_351),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_460),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_243),
.C(n_225),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_496),
.B(n_419),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_429),
.B(n_307),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_429),
.B(n_216),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_429),
.B(n_216),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_432),
.B(n_312),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_499),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_467),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_467),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_498),
.B(n_441),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_467),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_498),
.A2(n_246),
.B1(n_337),
.B2(n_335),
.Y(n_584)
);

BUFx10_ASAP7_75t_L g585 ( 
.A(n_455),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_497),
.A2(n_312),
.B(n_306),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_473),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_498),
.A2(n_456),
.B1(n_494),
.B2(n_441),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_476),
.A2(n_247),
.B1(n_335),
.B2(n_261),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_467),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_467),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_467),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_431),
.B(n_286),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_457),
.B(n_216),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_498),
.A2(n_495),
.B1(n_492),
.B2(n_457),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_431),
.B(n_300),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_425),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_368),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_431),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_478),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_457),
.B(n_172),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_425),
.A2(n_313),
.B1(n_249),
.B2(n_257),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_478),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_495),
.B(n_362),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_472),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_478),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_441),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_472),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_441),
.A2(n_175),
.B1(n_199),
.B2(n_211),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_472),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_478),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_478),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_472),
.B(n_247),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_493),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_497),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_171),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_436),
.Y(n_622)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_478),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_482),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_482),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_482),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_492),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_493),
.B(n_376),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_493),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_482),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_482),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_482),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_441),
.B(n_259),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_482),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_477),
.B(n_420),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_486),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_486),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_486),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_436),
.B(n_173),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_492),
.B(n_321),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_432),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_441),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_486),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_436),
.B(n_442),
.C(n_440),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_486),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_486),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_440),
.B(n_442),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_486),
.Y(n_651)
);

NOR2x1p5_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_445),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_620),
.B(n_440),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_L g655 ( 
.A1(n_548),
.A2(n_234),
.B1(n_199),
.B2(n_284),
.C(n_316),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_599),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_508),
.B(n_473),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_528),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_585),
.B(n_442),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_443),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_543),
.A2(n_470),
.B(n_444),
.C(n_490),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_540),
.B(n_443),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_607),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_520),
.B(n_443),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_585),
.B(n_444),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_444),
.Y(n_667)
);

AO22x2_ASAP7_75t_L g668 ( 
.A1(n_509),
.A2(n_234),
.B1(n_211),
.B2(n_244),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_615),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_630),
.B(n_451),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_557),
.A2(n_244),
.B1(n_274),
.B2(n_284),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_627),
.B(n_451),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_573),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_607),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_599),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_524),
.A2(n_445),
.B1(n_477),
.B2(n_490),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_573),
.B(n_451),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_611),
.A2(n_463),
.B(n_462),
.C(n_490),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_529),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_521),
.B(n_462),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_634),
.A2(n_494),
.B1(n_456),
.B2(n_466),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_574),
.B(n_462),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_503),
.B(n_463),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_599),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_650),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_574),
.B(n_463),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_622),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_517),
.B(n_464),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_531),
.A2(n_479),
.B1(n_464),
.B2(n_489),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_595),
.B(n_464),
.Y(n_692)
);

BUFx12f_ASAP7_75t_SL g693 ( 
.A(n_524),
.Y(n_693)
);

BUFx5_ASAP7_75t_L g694 ( 
.A(n_582),
.Y(n_694)
);

AND2x4_ASAP7_75t_SL g695 ( 
.A(n_595),
.B(n_378),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_644),
.A2(n_471),
.B(n_470),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_642),
.B(n_470),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_585),
.B(n_471),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_634),
.A2(n_494),
.B1(n_456),
.B2(n_438),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_642),
.B(n_471),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_531),
.B(n_486),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_536),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_644),
.A2(n_484),
.B(n_479),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_523),
.B(n_479),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_502),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_571),
.B(n_484),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_643),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_545),
.B(n_484),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_531),
.B(n_488),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_531),
.A2(n_488),
.B1(n_489),
.B2(n_434),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_542),
.B(n_381),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_611),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_643),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_523),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_563),
.B(n_488),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_502),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_550),
.A2(n_489),
.B(n_434),
.C(n_450),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_551),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_628),
.B(n_434),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_531),
.B(n_434),
.Y(n_723)
);

AO221x1_ASAP7_75t_L g724 ( 
.A1(n_590),
.A2(n_334),
.B1(n_319),
.B2(n_320),
.C(n_322),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_531),
.A2(n_461),
.B1(n_435),
.B2(n_487),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_569),
.B(n_435),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_569),
.B(n_435),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_584),
.A2(n_494),
.B1(n_456),
.B2(n_487),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_600),
.B(n_435),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_SL g730 ( 
.A(n_526),
.B(n_386),
.C(n_383),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_522),
.B(n_438),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_618),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_504),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_569),
.B(n_438),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_559),
.B(n_438),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_512),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_602),
.B(n_448),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_602),
.B(n_448),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_518),
.A2(n_449),
.B(n_448),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_524),
.B(n_423),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_512),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_501),
.B(n_448),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_512),
.B(n_449),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_608),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_504),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_602),
.B(n_449),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_501),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_619),
.B(n_449),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_507),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_619),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_619),
.B(n_450),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_572),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_572),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_594),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_604),
.B(n_572),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_604),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_605),
.B(n_450),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_507),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_604),
.B(n_450),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_608),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_575),
.A2(n_481),
.B1(n_466),
.B2(n_487),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_575),
.A2(n_481),
.B1(n_466),
.B2(n_487),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_516),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_516),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_604),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_575),
.A2(n_466),
.B1(n_461),
.B2(n_483),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_530),
.B(n_461),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_461),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_568),
.B(n_465),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_544),
.B(n_641),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_465),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_590),
.A2(n_465),
.B1(n_481),
.B2(n_483),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_590),
.A2(n_465),
.B1(n_481),
.B2(n_483),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_582),
.B(n_483),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_524),
.B(n_391),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_590),
.A2(n_494),
.B1(n_456),
.B2(n_468),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_575),
.B(n_432),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_527),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_575),
.B(n_432),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_527),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_538),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_614),
.B(n_553),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_575),
.B(n_432),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_538),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_512),
.B(n_267),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_512),
.Y(n_786)
);

AND2x2_ASAP7_75t_SL g787 ( 
.A(n_589),
.B(n_456),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_546),
.Y(n_788)
);

INVx8_ASAP7_75t_L g789 ( 
.A(n_513),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_558),
.B(n_432),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_546),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_558),
.A2(n_494),
.B1(n_491),
.B2(n_468),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_549),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_513),
.B(n_272),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_549),
.Y(n_795)
);

AND2x4_ASAP7_75t_SL g796 ( 
.A(n_537),
.B(n_392),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_637),
.B(n_468),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_513),
.B(n_491),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_586),
.B(n_468),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_554),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_510),
.B(n_468),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_586),
.B(n_468),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_554),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_586),
.A2(n_491),
.B1(n_288),
.B2(n_213),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_588),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_588),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_510),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_555),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_511),
.B(n_491),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_555),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_511),
.B(n_552),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_513),
.B(n_491),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_556),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_556),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_513),
.B(n_567),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_511),
.B(n_393),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_567),
.B(n_306),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_561),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_552),
.B(n_273),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_552),
.B(n_279),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_662),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_654),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_696),
.A2(n_505),
.B(n_500),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_665),
.B(n_631),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_673),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_705),
.A2(n_505),
.B(n_500),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_811),
.A2(n_660),
.B(n_726),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_727),
.A2(n_515),
.B(n_506),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_754),
.A2(n_515),
.B(n_506),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_734),
.A2(n_525),
.B(n_519),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_737),
.A2(n_525),
.B(n_519),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_755),
.B(n_631),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_695),
.B(n_395),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_695),
.B(n_397),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_746),
.A2(n_533),
.B(n_532),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_681),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_653),
.B(n_631),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_681),
.B(n_567),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_684),
.A2(n_649),
.B(n_565),
.C(n_648),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_751),
.A2(n_533),
.B(n_532),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_713),
.B(n_398),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_663),
.B(n_649),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_815),
.A2(n_774),
.B(n_768),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_708),
.B(n_649),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_789),
.Y(n_845)
);

OAI321xp33_ASAP7_75t_L g846 ( 
.A1(n_655),
.A2(n_246),
.A3(n_322),
.B1(n_319),
.B2(n_316),
.C(n_260),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_687),
.A2(n_587),
.B1(n_539),
.B2(n_646),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_815),
.A2(n_539),
.B(n_534),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_714),
.A2(n_587),
.B1(n_547),
.B2(n_646),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_708),
.B(n_561),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_771),
.A2(n_547),
.B(n_534),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_755),
.B(n_567),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_658),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_771),
.A2(n_564),
.B(n_562),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_677),
.B(n_565),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_678),
.A2(n_564),
.B(n_562),
.Y(n_856)
);

O2A1O1Ixp5_ASAP7_75t_L g857 ( 
.A1(n_769),
.A2(n_581),
.B(n_648),
.C(n_645),
.Y(n_857)
);

CKINVDCx16_ASAP7_75t_R g858 ( 
.A(n_730),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_738),
.A2(n_576),
.B(n_570),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_747),
.B(n_566),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_744),
.B(n_760),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_683),
.B(n_566),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_676),
.B(n_567),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_782),
.A2(n_320),
.B1(n_256),
.B2(n_321),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_570),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_756),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_688),
.B(n_581),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_765),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_709),
.B(n_591),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_817),
.A2(n_748),
.B(n_770),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_657),
.B(n_692),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_711),
.A2(n_577),
.B(n_576),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_693),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_674),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_L g875 ( 
.A1(n_731),
.A2(n_606),
.B(n_645),
.C(n_596),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_817),
.A2(n_739),
.B(n_799),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_669),
.A2(n_578),
.B(n_577),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_697),
.B(n_701),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_652),
.B(n_596),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_789),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_716),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_686),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_805),
.B(n_321),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_752),
.B(n_606),
.Y(n_884)
);

AOI21x1_ASAP7_75t_L g885 ( 
.A1(n_802),
.A2(n_580),
.B(n_578),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_684),
.A2(n_629),
.B(n_632),
.C(n_639),
.Y(n_886)
);

OR2x2_ASAP7_75t_SL g887 ( 
.A(n_740),
.B(n_256),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_671),
.A2(n_330),
.B1(n_427),
.B2(n_426),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_723),
.A2(n_583),
.B(n_580),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_671),
.A2(n_330),
.B1(n_427),
.B2(n_426),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_667),
.A2(n_592),
.B(n_583),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_789),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_670),
.A2(n_593),
.B(n_592),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_674),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_664),
.B(n_623),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_777),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_706),
.B(n_672),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_721),
.A2(n_626),
.B(n_640),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_593),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_690),
.A2(n_629),
.B(n_632),
.C(n_639),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_750),
.A2(n_610),
.B(n_640),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_806),
.B(n_601),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_690),
.A2(n_680),
.B(n_759),
.C(n_710),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_702),
.A2(n_610),
.B(n_638),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_718),
.A2(n_666),
.B(n_659),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_796),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_698),
.A2(n_613),
.B(n_638),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_809),
.A2(n_613),
.B(n_636),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_710),
.B(n_635),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_682),
.A2(n_601),
.B(n_636),
.Y(n_911)
);

AO21x1_ASAP7_75t_L g912 ( 
.A1(n_680),
.A2(n_616),
.B(n_617),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_SL g913 ( 
.A1(n_689),
.A2(n_617),
.B(n_603),
.C(n_633),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_732),
.A2(n_633),
.B(n_626),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_759),
.B(n_635),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_682),
.A2(n_603),
.B(n_616),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_735),
.B(n_591),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_707),
.A2(n_625),
.B(n_591),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_674),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_735),
.B(n_797),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_707),
.A2(n_625),
.B(n_591),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_797),
.B(n_591),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_719),
.A2(n_625),
.B(n_651),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_719),
.A2(n_625),
.B(n_651),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_715),
.B(n_625),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_733),
.A2(n_651),
.B(n_624),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_699),
.B(n_623),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_733),
.A2(n_651),
.B(n_624),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_720),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_700),
.A2(n_651),
.B(n_624),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_745),
.A2(n_758),
.B(n_749),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_745),
.A2(n_624),
.B(n_623),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_729),
.B(n_623),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_816),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_661),
.A2(n_514),
.B(n_427),
.C(n_426),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_767),
.A2(n_514),
.B(n_424),
.C(n_299),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_749),
.A2(n_624),
.B(n_623),
.Y(n_937)
);

CKINVDCx6p67_ASAP7_75t_R g938 ( 
.A(n_775),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_722),
.A2(n_314),
.B(n_287),
.C(n_340),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_L g940 ( 
.A1(n_819),
.A2(n_283),
.B(n_303),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_656),
.B(n_308),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_758),
.A2(n_183),
.B(n_177),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_SL g943 ( 
.A1(n_691),
.A2(n_757),
.B(n_712),
.C(n_801),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_781),
.A2(n_791),
.B(n_784),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_722),
.A2(n_338),
.B(n_328),
.C(n_311),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_675),
.B(n_178),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_790),
.B(n_424),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_753),
.B(n_424),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_700),
.A2(n_424),
.B(n_266),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_801),
.A2(n_790),
.B(n_819),
.C(n_820),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_812),
.A2(n_2),
.B(n_3),
.C(n_6),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_763),
.A2(n_265),
.B(n_339),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_664),
.A2(n_258),
.B1(n_186),
.B2(n_332),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_674),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_820),
.A2(n_428),
.B(n_268),
.C(n_329),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_793),
.A2(n_252),
.B(n_194),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_792),
.A2(n_276),
.B1(n_195),
.B2(n_327),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_792),
.A2(n_242),
.B1(n_197),
.B2(n_323),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_694),
.B(n_2),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_685),
.B(n_185),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_763),
.A2(n_278),
.B(n_201),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_777),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_668),
.B(n_428),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_694),
.B(n_200),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_764),
.A2(n_292),
.B(n_217),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_694),
.B(n_6),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_812),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_761),
.B(n_203),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_728),
.A2(n_818),
.B(n_778),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_800),
.A2(n_428),
.B(n_333),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_668),
.B(n_679),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_668),
.B(n_219),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_764),
.A2(n_295),
.B(n_222),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_679),
.B(n_221),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_787),
.A2(n_297),
.B1(n_229),
.B2(n_318),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_778),
.A2(n_302),
.B(n_237),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_762),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_798),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_803),
.A2(n_309),
.B(n_239),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_772),
.A2(n_15),
.B(n_16),
.C(n_19),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_813),
.A2(n_310),
.B(n_281),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_766),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_814),
.A2(n_317),
.B(n_315),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_773),
.A2(n_16),
.B(n_20),
.C(n_22),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_694),
.A2(n_294),
.B1(n_428),
.B2(n_333),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_796),
.B(n_23),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_787),
.A2(n_428),
.B1(n_333),
.B2(n_238),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_694),
.B(n_783),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_780),
.A2(n_818),
.B(n_788),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_785),
.B(n_24),
.C(n_25),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_671),
.B(n_428),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_779),
.B(n_428),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_780),
.A2(n_333),
.B(n_238),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_786),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_704),
.B(n_24),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_333),
.B(n_238),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_736),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_807),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_786),
.B(n_428),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_694),
.A2(n_428),
.B1(n_238),
.B2(n_223),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_807),
.B(n_31),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_804),
.B(n_32),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_795),
.A2(n_238),
.B(n_223),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_736),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_736),
.A2(n_223),
.B1(n_34),
.B2(n_36),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_L g1006 ( 
.A(n_794),
.B(n_33),
.C(n_41),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_725),
.A2(n_223),
.B(n_43),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_795),
.A2(n_808),
.B(n_743),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_962),
.B(n_741),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_987),
.A2(n_808),
.B(n_810),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_871),
.B(n_703),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_950),
.A2(n_741),
.B(n_736),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_962),
.B(n_741),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_871),
.B(n_741),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_897),
.B(n_776),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_827),
.A2(n_728),
.B(n_776),
.Y(n_1016)
);

BUFx2_ASAP7_75t_SL g1017 ( 
.A(n_906),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_883),
.B(n_724),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_850),
.A2(n_223),
.B(n_104),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_873),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_832),
.B(n_41),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_880),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_1002),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_903),
.A2(n_44),
.B1(n_46),
.B2(n_49),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_959),
.A2(n_49),
.B(n_51),
.C(n_53),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_960),
.B(n_53),
.C(n_56),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_938),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_907),
.B(n_56),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_846),
.A2(n_60),
.B1(n_66),
.B2(n_68),
.C(n_71),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_907),
.B(n_76),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_944),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_880),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_994),
.B(n_93),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_SL g1034 ( 
.A1(n_959),
.A2(n_105),
.B(n_112),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_841),
.B(n_118),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_878),
.A2(n_123),
.B1(n_130),
.B2(n_140),
.Y(n_1036)
);

CKINVDCx6p67_ASAP7_75t_R g1037 ( 
.A(n_833),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_966),
.A2(n_146),
.B1(n_152),
.B2(n_159),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_845),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_844),
.A2(n_161),
.B(n_163),
.C(n_168),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_861),
.A2(n_169),
.B1(n_966),
.B2(n_825),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_880),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_920),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_882),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_970),
.A2(n_876),
.B(n_885),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_899),
.A2(n_943),
.B(n_842),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_825),
.A2(n_941),
.B1(n_822),
.B2(n_902),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_896),
.B(n_866),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_880),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_SL g1050 ( 
.A1(n_1005),
.A2(n_863),
.B(n_925),
.C(n_869),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_939),
.A2(n_945),
.B(n_940),
.C(n_984),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_1007),
.B(n_845),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_980),
.A2(n_822),
.B(n_998),
.C(n_951),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_832),
.B(n_852),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_858),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_834),
.B(n_934),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_899),
.A2(n_854),
.B(n_851),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_1004),
.B(n_836),
.Y(n_1058)
);

OAI21xp33_ASAP7_75t_SL g1059 ( 
.A1(n_1001),
.A2(n_865),
.B(n_981),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_977),
.B(n_982),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_967),
.B(n_865),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_892),
.B(n_836),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_892),
.B(n_860),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_881),
.B(n_887),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_855),
.B(n_862),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_829),
.A2(n_912),
.B(n_989),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_919),
.B(n_874),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_881),
.B(n_946),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_824),
.A2(n_843),
.B(n_826),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_823),
.A2(n_917),
.B(n_889),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_919),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_971),
.B(n_866),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_884),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_867),
.A2(n_872),
.B(n_918),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_921),
.A2(n_898),
.B(n_830),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_868),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_868),
.B(n_879),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_955),
.A2(n_838),
.B(n_857),
.C(n_979),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_864),
.B(n_888),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_954),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_828),
.A2(n_831),
.B(n_835),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_915),
.B(n_910),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_990),
.B1(n_1006),
.B2(n_890),
.C(n_888),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_986),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_978),
.A2(n_1006),
.B(n_990),
.C(n_839),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_954),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_SL g1087 ( 
.A(n_905),
.B(n_956),
.C(n_983),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_860),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_837),
.B(n_929),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_964),
.A2(n_922),
.B(n_914),
.C(n_995),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_968),
.A2(n_927),
.B(n_985),
.C(n_847),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_988),
.B(n_992),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_954),
.B(n_953),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_954),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_840),
.A2(n_877),
.B(n_891),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_963),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_874),
.B(n_894),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_890),
.A2(n_849),
.B1(n_947),
.B2(n_911),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_972),
.B(n_948),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_930),
.A2(n_916),
.B(n_870),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_895),
.B(n_991),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_913),
.A2(n_900),
.B(n_886),
.C(n_975),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_969),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_992),
.B(n_894),
.Y(n_1104)
);

OAI21xp33_ASAP7_75t_SL g1105 ( 
.A1(n_856),
.A2(n_997),
.B(n_933),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_857),
.A2(n_875),
.B(n_932),
.C(n_937),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_957),
.B(n_958),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_997),
.B(n_999),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_931),
.B(n_999),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_908),
.A2(n_893),
.B(n_848),
.C(n_909),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_974),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1000),
.A2(n_904),
.B1(n_895),
.B2(n_949),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_SL g1113 ( 
.A(n_901),
.B(n_859),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_926),
.A2(n_928),
.B(n_923),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_924),
.B(n_1008),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_875),
.A2(n_935),
.B(n_936),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_942),
.B(n_952),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_961),
.A2(n_965),
.B(n_973),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_976),
.B(n_993),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_996),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_SL g1121 ( 
.A1(n_1003),
.A2(n_950),
.B(n_903),
.C(n_878),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1002),
.A2(n_588),
.B1(n_657),
.B2(n_755),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_871),
.B(n_620),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_903),
.A2(n_878),
.B1(n_897),
.B2(n_663),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_903),
.A2(n_1002),
.B(n_966),
.C(n_959),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_903),
.A2(n_548),
.B(n_665),
.C(n_542),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_871),
.B(n_620),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_987),
.A2(n_773),
.A3(n_772),
.B1(n_1005),
.B2(n_849),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_871),
.B(n_508),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_871),
.B(n_352),
.Y(n_1131)
);

AND2x4_ASAP7_75t_SL g1132 ( 
.A(n_906),
.B(n_962),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_871),
.A2(n_542),
.B1(n_1002),
.B2(n_548),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_822),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_903),
.A2(n_1002),
.B(n_966),
.C(n_959),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_871),
.B(n_620),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_903),
.A2(n_1002),
.B(n_966),
.C(n_959),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_873),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_903),
.A2(n_1002),
.B(n_966),
.C(n_959),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_L g1140 ( 
.A(n_878),
.B(n_903),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_903),
.A2(n_548),
.B(n_665),
.C(n_542),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_906),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_903),
.A2(n_548),
.B(n_665),
.C(n_542),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_871),
.B(n_805),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_871),
.B(n_878),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_871),
.B(n_878),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_871),
.B(n_620),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_903),
.A2(n_1002),
.B(n_966),
.C(n_959),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_853),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_833),
.B(n_755),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_821),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_821),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_871),
.B(n_508),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_871),
.B(n_805),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_950),
.A2(n_705),
.B(n_696),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_871),
.B(n_508),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1058),
.Y(n_1162)
);

BUFx4_ASAP7_75t_SL g1163 ( 
.A(n_1143),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1031),
.A2(n_1103),
.A3(n_1090),
.B(n_1137),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1044),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_1014),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1133),
.A2(n_1131),
.B1(n_1041),
.B2(n_1047),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_SL g1168 ( 
.A(n_1020),
.Y(n_1168)
);

AOI221x1_ASAP7_75t_L g1169 ( 
.A1(n_1125),
.A2(n_1151),
.B1(n_1139),
.B2(n_1135),
.C(n_1024),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_1095),
.A2(n_1081),
.B(n_1070),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1055),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1134),
.B(n_1153),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1009),
.Y(n_1175)
);

INVx3_ASAP7_75t_R g1176 ( 
.A(n_1021),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_1132),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1148),
.A2(n_1149),
.B1(n_1107),
.B2(n_1124),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1024),
.A2(n_1023),
.B(n_1126),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1010),
.A2(n_1066),
.B(n_1113),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1149),
.A2(n_1124),
.B1(n_1083),
.B2(n_1061),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1046),
.A2(n_1140),
.B(n_1159),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1153),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1153),
.B(n_1123),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_1048),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1128),
.A2(n_1145),
.B(n_1157),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1141),
.A2(n_1146),
.B(n_1059),
.C(n_1051),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_SL g1188 ( 
.A(n_1026),
.B(n_1087),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1130),
.A2(n_1160),
.B(n_1156),
.C(n_1025),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1127),
.B(n_1136),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1142),
.A2(n_1144),
.B(n_1057),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1069),
.A2(n_1106),
.B(n_1116),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1098),
.A2(n_1016),
.B(n_1050),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1076),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1027),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1150),
.B(n_1060),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1114),
.A2(n_1012),
.B(n_1116),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1028),
.A2(n_1068),
.B(n_1085),
.C(n_1121),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1065),
.A2(n_1082),
.B(n_1112),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1138),
.B(n_1122),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1152),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1065),
.A2(n_1082),
.B(n_1112),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1009),
.Y(n_1203)
);

AOI221xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1053),
.A2(n_1098),
.B1(n_1061),
.B2(n_1034),
.C(n_1089),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1089),
.A2(n_1079),
.B1(n_1060),
.B2(n_1015),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1088),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1102),
.A2(n_1109),
.B(n_1019),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1011),
.B(n_1052),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1035),
.A2(n_1038),
.B(n_1091),
.C(n_1036),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1027),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1022),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1029),
.A2(n_1077),
.B(n_1018),
.C(n_1111),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1037),
.Y(n_1213)
);

CKINVDCx6p67_ASAP7_75t_R g1214 ( 
.A(n_1017),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1021),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1064),
.B(n_1084),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1078),
.A2(n_1105),
.B(n_1030),
.C(n_1052),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1056),
.B(n_1054),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1154),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1100),
.A2(n_1109),
.B(n_1118),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1155),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1108),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_SL g1223 ( 
.A1(n_1093),
.A2(n_1033),
.B(n_1062),
.C(n_1110),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1115),
.A2(n_1120),
.B(n_1119),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1022),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1104),
.B(n_1073),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1096),
.B(n_1099),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1022),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1117),
.A2(n_1115),
.B(n_1100),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1092),
.A2(n_1038),
.B(n_1067),
.Y(n_1230)
);

AOI21xp33_ASAP7_75t_L g1231 ( 
.A1(n_1072),
.A2(n_1092),
.B(n_1036),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1072),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1063),
.A2(n_1013),
.B(n_1129),
.C(n_1071),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1072),
.B(n_1013),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1101),
.A2(n_1097),
.B1(n_1032),
.B2(n_1049),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1032),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_SL g1237 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1101),
.A2(n_1129),
.B1(n_1039),
.B2(n_1071),
.Y(n_1238)
);

INVx3_ASAP7_75t_SL g1239 ( 
.A(n_1042),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1101),
.A2(n_1129),
.B(n_1040),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1067),
.A2(n_1086),
.B(n_1080),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1042),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1049),
.A2(n_1094),
.B(n_1080),
.C(n_1086),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1080),
.B(n_1094),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1094),
.A2(n_1046),
.B(n_1140),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1049),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_1138),
.B(n_1047),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1125),
.A2(n_1135),
.B1(n_1139),
.B2(n_1137),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1044),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1044),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1131),
.A2(n_588),
.B1(n_524),
.B2(n_557),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_1132),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1044),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1134),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1027),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1146),
.C(n_1126),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1014),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1027),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1125),
.A2(n_1137),
.B(n_1135),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1133),
.A2(n_1131),
.B1(n_871),
.B2(n_1147),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1101),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1133),
.A2(n_1131),
.B1(n_871),
.B2(n_1147),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1020),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1134),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1125),
.A2(n_1137),
.B(n_1135),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1046),
.A2(n_1140),
.B(n_1135),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1020),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1134),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1014),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1058),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1044),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1046),
.A2(n_1140),
.B(n_1135),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1146),
.C(n_1126),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1146),
.C(n_1126),
.Y(n_1285)
);

AOI211x1_ASAP7_75t_L g1286 ( 
.A1(n_1024),
.A2(n_676),
.B(n_1130),
.C(n_1156),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1020),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1146),
.C(n_1126),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_1132),
.Y(n_1289)
);

AOI221x1_ASAP7_75t_L g1290 ( 
.A1(n_1125),
.A2(n_1135),
.B1(n_1151),
.B2(n_1139),
.C(n_1137),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1058),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1294)
);

AND2x6_ASAP7_75t_L g1295 ( 
.A(n_1021),
.B(n_755),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1046),
.A2(n_1140),
.B(n_1135),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1043),
.B(n_1148),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1045),
.A2(n_1074),
.B(n_1075),
.Y(n_1298)
);

AO21x1_ASAP7_75t_L g1299 ( 
.A1(n_1107),
.A2(n_1002),
.B(n_1124),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1146),
.C(n_1126),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_L g1301 ( 
.A(n_1133),
.B(n_1135),
.C(n_1125),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1125),
.A2(n_1137),
.B(n_1135),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1044),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1044),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1024),
.A2(n_1124),
.A3(n_1098),
.B1(n_1112),
.B2(n_485),
.Y(n_1305)
);

AOI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1010),
.A2(n_1066),
.B(n_1113),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1009),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1009),
.B(n_1013),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1031),
.A2(n_829),
.A3(n_912),
.B(n_1103),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1054),
.B(n_962),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1046),
.A2(n_1140),
.B(n_1135),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1044),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1301),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1165),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1287),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1252),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1162),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1249),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1168),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1161),
.B(n_1262),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1225),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1299),
.A2(n_1167),
.B1(n_1301),
.B2(n_1253),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1210),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1228),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1263),
.A2(n_1265),
.B1(n_1169),
.B2(n_1290),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1279),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1178),
.A2(n_1181),
.B1(n_1261),
.B2(n_1270),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1178),
.A2(n_1181),
.B1(n_1261),
.B2(n_1270),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1255),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1280),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1211),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1303),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1266),
.B(n_1271),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1177),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1302),
.A2(n_1248),
.B1(n_1307),
.B2(n_1205),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1172),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1304),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1315),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1201),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1275),
.B(n_1297),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1302),
.A2(n_1248),
.B1(n_1205),
.B2(n_1251),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1251),
.B(n_1281),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1295),
.A2(n_1305),
.B1(n_1196),
.B2(n_1193),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1254),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1314),
.A2(n_1281),
.B1(n_1188),
.B2(n_1295),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1258),
.A2(n_1285),
.B1(n_1284),
.B2(n_1288),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1256),
.B(n_1276),
.Y(n_1352)
);

BUFx8_ASAP7_75t_L g1353 ( 
.A(n_1168),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1179),
.A2(n_1314),
.B1(n_1190),
.B2(n_1247),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1295),
.A2(n_1200),
.B1(n_1208),
.B2(n_1227),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1185),
.B(n_1166),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1254),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1219),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1289),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1221),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1226),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1257),
.Y(n_1362)
);

INVx8_ASAP7_75t_L g1363 ( 
.A(n_1295),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1179),
.A2(n_1305),
.B1(n_1215),
.B2(n_1202),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1273),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1273),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1195),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1305),
.A2(n_1199),
.B1(n_1296),
.B2(n_1283),
.Y(n_1368)
);

CKINVDCx6p67_ASAP7_75t_R g1369 ( 
.A(n_1260),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1226),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1214),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1209),
.A2(n_1198),
.B(n_1300),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1272),
.A2(n_1313),
.B1(n_1276),
.B2(n_1256),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1163),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1195),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1269),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1268),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1264),
.B(n_1237),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1213),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1164),
.Y(n_1380)
);

BUFx2_ASAP7_75t_SL g1381 ( 
.A(n_1206),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1194),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1239),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1187),
.A2(n_1286),
.B1(n_1189),
.B2(n_1212),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1211),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1184),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1216),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1222),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1259),
.A2(n_1278),
.B1(n_1182),
.B2(n_1217),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1193),
.A2(n_1231),
.B1(n_1218),
.B2(n_1183),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1309),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1231),
.A2(n_1183),
.B1(n_1222),
.B2(n_1311),
.Y(n_1392)
);

INVxp33_ASAP7_75t_L g1393 ( 
.A(n_1234),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1311),
.B(n_1203),
.Y(n_1394)
);

BUFx4_ASAP7_75t_SL g1395 ( 
.A(n_1176),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1175),
.B(n_1308),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1238),
.A2(n_1264),
.B1(n_1204),
.B2(n_1191),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1238),
.A2(n_1264),
.B1(n_1204),
.B2(n_1191),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1242),
.Y(n_1399)
);

INVx6_ASAP7_75t_L g1400 ( 
.A(n_1175),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1234),
.A2(n_1232),
.B1(n_1308),
.B2(n_1203),
.Y(n_1401)
);

BUFx2_ASAP7_75t_SL g1402 ( 
.A(n_1246),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1246),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1235),
.A2(n_1186),
.B1(n_1220),
.B2(n_1207),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1233),
.B(n_1236),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1240),
.A2(n_1244),
.B1(n_1245),
.B2(n_1229),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1230),
.A2(n_1223),
.B1(n_1244),
.B2(n_1243),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1164),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1220),
.A2(n_1192),
.B1(n_1170),
.B2(n_1197),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1192),
.A2(n_1170),
.B1(n_1241),
.B2(n_1171),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1164),
.A2(n_1298),
.B1(n_1291),
.B2(n_1267),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1224),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1310),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1180),
.A2(n_1306),
.B1(n_1310),
.B2(n_1282),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1274),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1277),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1294),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1133),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1162),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1211),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1165),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1307),
.B(n_1147),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1195),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1263),
.A2(n_1265),
.B1(n_1293),
.B2(n_1250),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1168),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1133),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1165),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1133),
.Y(n_1428)
);

OAI22x1_ASAP7_75t_SL g1429 ( 
.A1(n_1172),
.A2(n_480),
.B1(n_499),
.B2(n_452),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1161),
.B(n_1262),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1299),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1312),
.B2(n_1299),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1161),
.B(n_1262),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1177),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1177),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1210),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1250),
.A2(n_1312),
.B1(n_1293),
.B2(n_1133),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1228),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1250),
.A2(n_1312),
.B(n_1293),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1166),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1162),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1210),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1168),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1415),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1362),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1351),
.B(n_1389),
.Y(n_1446)
);

INVxp33_ASAP7_75t_L g1447 ( 
.A(n_1422),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1409),
.A2(n_1410),
.B(n_1404),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1418),
.A2(n_1426),
.B1(n_1428),
.B2(n_1348),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1441),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1382),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1416),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1343),
.B(n_1330),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1362),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1408),
.B(n_1380),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1356),
.B(n_1440),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1330),
.B(n_1331),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1409),
.A2(n_1410),
.B(n_1404),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1407),
.A2(n_1413),
.B(n_1331),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1398),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1397),
.B(n_1398),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1437),
.A2(n_1432),
.B1(n_1431),
.B2(n_1439),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1352),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1317),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1321),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1381),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1332),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1333),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1415),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1335),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1347),
.B(n_1316),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1417),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1358),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1340),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1342),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1348),
.A2(n_1328),
.B1(n_1354),
.B2(n_1325),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1341),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1436),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1403),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1360),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1365),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1424),
.A2(n_1345),
.B1(n_1325),
.B2(n_1372),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1363),
.B(n_1412),
.Y(n_1484)
);

BUFx8_ASAP7_75t_SL g1485 ( 
.A(n_1318),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1436),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1421),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1427),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1338),
.B(n_1345),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1424),
.B(n_1323),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1414),
.A2(n_1406),
.B(n_1364),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1441),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1384),
.A2(n_1390),
.B(n_1405),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1406),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1338),
.B(n_1386),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1419),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1361),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1429),
.B(n_1326),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1370),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1319),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1393),
.B(n_1388),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1376),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1364),
.Y(n_1503)
);

AOI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1396),
.A2(n_1433),
.B(n_1430),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1390),
.A2(n_1378),
.B(n_1392),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1378),
.A2(n_1392),
.B(n_1350),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1322),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1320),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1387),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1368),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1368),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1373),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1350),
.A2(n_1401),
.B(n_1355),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1336),
.A2(n_1344),
.B(n_1394),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1393),
.B(n_1411),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1373),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1414),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1355),
.A2(n_1334),
.B(n_1420),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1354),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1377),
.B(n_1339),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1328),
.A2(n_1438),
.B(n_1327),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1329),
.B(n_1402),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1400),
.B(n_1366),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1324),
.B(n_1385),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1442),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1391),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1367),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1324),
.B(n_1383),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1324),
.B(n_1423),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1470),
.B(n_1324),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1500),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1456),
.B(n_1383),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1470),
.B(n_1399),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1485),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1515),
.B(n_1322),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1374),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1491),
.A2(n_1395),
.B(n_1435),
.Y(n_1538)
);

AO21x1_ASAP7_75t_L g1539 ( 
.A1(n_1462),
.A2(n_1395),
.B(n_1425),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1482),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1470),
.B(n_1371),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1450),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1446),
.A2(n_1379),
.B(n_1425),
.C(n_1443),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1446),
.A2(n_1443),
.B(n_1353),
.C(n_1375),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1460),
.A2(n_1353),
.B1(n_1369),
.B2(n_1442),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_L g1546 ( 
.A(n_1449),
.B(n_1375),
.C(n_1435),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1346),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_SL g1548 ( 
.A(n_1454),
.B(n_1357),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1491),
.B(n_1337),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1491),
.B(n_1337),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1454),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1450),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_L g1553 ( 
.A(n_1483),
.B(n_1349),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1509),
.B(n_1359),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1502),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1477),
.A2(n_1434),
.B(n_1435),
.C(n_1472),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1458),
.A2(n_1434),
.B(n_1494),
.Y(n_1557)
);

AOI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1463),
.A2(n_1503),
.B1(n_1511),
.B2(n_1510),
.C(n_1461),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1493),
.A2(n_1490),
.B(n_1457),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1484),
.B(n_1480),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1517),
.B(n_1453),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1460),
.A2(n_1461),
.B(n_1493),
.C(n_1494),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1489),
.A2(n_1457),
.B(n_1519),
.C(n_1503),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1489),
.A2(n_1519),
.B(n_1512),
.C(n_1516),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1513),
.A2(n_1444),
.B1(n_1495),
.B2(n_1521),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1448),
.B(n_1512),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1464),
.B(n_1451),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1516),
.A2(n_1521),
.B(n_1459),
.Y(n_1570)
);

AO21x2_ASAP7_75t_L g1571 ( 
.A1(n_1514),
.A2(n_1504),
.B(n_1505),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1459),
.A2(n_1505),
.B(n_1506),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1464),
.B(n_1451),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1448),
.B(n_1465),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1474),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1521),
.A2(n_1504),
.B(n_1506),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1521),
.A2(n_1518),
.B(n_1467),
.Y(n_1577)
);

CKINVDCx8_ASAP7_75t_R g1578 ( 
.A(n_1445),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1496),
.A2(n_1508),
.B1(n_1527),
.B2(n_1513),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1507),
.A2(n_1523),
.B(n_1527),
.C(n_1528),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1448),
.B(n_1465),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1513),
.A2(n_1447),
.B1(n_1522),
.B2(n_1492),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1466),
.B(n_1468),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1513),
.A2(n_1495),
.B1(n_1526),
.B2(n_1444),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1480),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1474),
.B(n_1481),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1466),
.B(n_1468),
.Y(n_1587)
);

AND2x2_ASAP7_75t_SL g1588 ( 
.A(n_1444),
.B(n_1452),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1444),
.A2(n_1498),
.B(n_1452),
.C(n_1518),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1497),
.B(n_1499),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1469),
.B(n_1471),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1469),
.B(n_1478),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1471),
.B(n_1478),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1497),
.B(n_1499),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1574),
.B(n_1487),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1564),
.B(n_1473),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1581),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1564),
.B(n_1568),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1583),
.B(n_1455),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1488),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1538),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1587),
.B(n_1455),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1587),
.B(n_1455),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1591),
.B(n_1455),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1522),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1592),
.B(n_1475),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1532),
.Y(n_1610)
);

BUFx5_ASAP7_75t_L g1611 ( 
.A(n_1549),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1563),
.A2(n_1529),
.B1(n_1525),
.B2(n_1530),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1577),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1585),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1593),
.B(n_1562),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1590),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1555),
.Y(n_1618)
);

BUFx3_ASAP7_75t_R g1619 ( 
.A(n_1542),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1560),
.B(n_1501),
.Y(n_1620)
);

BUFx4f_ASAP7_75t_SL g1621 ( 
.A(n_1541),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1594),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1559),
.B(n_1585),
.Y(n_1623)
);

AND2x2_ASAP7_75t_SL g1624 ( 
.A(n_1603),
.B(n_1549),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1616),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1613),
.A2(n_1539),
.B1(n_1558),
.B2(n_1553),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1598),
.B(n_1615),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1613),
.A2(n_1539),
.B1(n_1553),
.B2(n_1579),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1612),
.A2(n_1567),
.B1(n_1546),
.B2(n_1570),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1599),
.A2(n_1565),
.B1(n_1566),
.B2(n_1612),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1599),
.B(n_1569),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1608),
.A2(n_1584),
.B1(n_1550),
.B2(n_1582),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1615),
.B(n_1550),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1611),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1622),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1557),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1608),
.A2(n_1556),
.B1(n_1544),
.B2(n_1543),
.C(n_1576),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1604),
.B(n_1605),
.Y(n_1640)
);

AOI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1619),
.A2(n_1535),
.B(n_1551),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1618),
.B(n_1533),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1603),
.A2(n_1571),
.B(n_1572),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1601),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1571),
.B(n_1589),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1601),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1552),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1597),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1618),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1606),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1606),
.Y(n_1651)
);

AOI211x1_ASAP7_75t_SL g1652 ( 
.A1(n_1620),
.A2(n_1578),
.B(n_1486),
.C(n_1573),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1627),
.B(n_1605),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1650),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1648),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1650),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1641),
.B(n_1621),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1637),
.B(n_1602),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1650),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1605),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1642),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1637),
.B(n_1602),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1637),
.B(n_1617),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1651),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1648),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1617),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1651),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1635),
.B(n_1595),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1648),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1595),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_1607),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1596),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1636),
.B(n_1603),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1636),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1625),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1651),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1634),
.B(n_1614),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1625),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1625),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1644),
.B(n_1646),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1674),
.B(n_1640),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1631),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1649),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1686),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1654),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1657),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1662),
.A2(n_1628),
.B1(n_1626),
.B2(n_1629),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1663),
.B(n_1631),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1663),
.B(n_1631),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1660),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1665),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1662),
.B(n_1486),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1664),
.B(n_1649),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1664),
.B(n_1631),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1658),
.B(n_1551),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1669),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1669),
.Y(n_1707)
);

NOR3xp33_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1639),
.C(n_1630),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1683),
.B(n_1642),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1628),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1658),
.B(n_1479),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1667),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1680),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1683),
.B(n_1647),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1667),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1655),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_1653),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1636),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1668),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1684),
.A2(n_1630),
.B1(n_1626),
.B2(n_1632),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1670),
.B(n_1647),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1655),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1674),
.B(n_1640),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1684),
.B(n_1647),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1680),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1728)
);

OR2x6_ASAP7_75t_L g1729 ( 
.A(n_1676),
.B(n_1603),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1708),
.B(n_1684),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1695),
.A2(n_1630),
.B(n_1677),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1704),
.B(n_1670),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1720),
.B(n_1661),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1661),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1688),
.B(n_1661),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1721),
.B(n_1666),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1689),
.B(n_1670),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1724),
.B(n_1666),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1710),
.B(n_1666),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1691),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1535),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1691),
.B(n_1671),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1696),
.B(n_1671),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1701),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1701),
.B(n_1548),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1687),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1729),
.A2(n_1639),
.B1(n_1632),
.B2(n_1629),
.C(n_1676),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1724),
.B(n_1671),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1692),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1718),
.B(n_1675),
.Y(n_1753)
);

NOR4xp25_ASAP7_75t_L g1754 ( 
.A(n_1690),
.B(n_1639),
.C(n_1540),
.D(n_1682),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1705),
.B(n_1524),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1719),
.B(n_1641),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_L g1758 ( 
.A(n_1729),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1718),
.B(n_1675),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1638),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1693),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1694),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1697),
.Y(n_1763)
);

OAI31xp33_ASAP7_75t_L g1764 ( 
.A1(n_1705),
.A2(n_1547),
.A3(n_1536),
.B(n_1545),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1727),
.B(n_1675),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1753),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1747),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1754),
.A2(n_1729),
.B(n_1711),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1732),
.A2(n_1624),
.B1(n_1547),
.B2(n_1538),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1748),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1748),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1751),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1754),
.A2(n_1703),
.B(n_1729),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1737),
.A2(n_1624),
.B1(n_1611),
.B2(n_1536),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1751),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1741),
.B(n_1727),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1746),
.B(n_1728),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1749),
.A2(n_1703),
.B(n_1723),
.C(n_1712),
.Y(n_1778)
);

INVxp33_ASAP7_75t_L g1779 ( 
.A(n_1747),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1755),
.B(n_1728),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1730),
.B(n_1722),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1761),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1747),
.A2(n_1624),
.B1(n_1538),
.B2(n_1611),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1761),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1762),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1755),
.B(n_1711),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1740),
.B(n_1726),
.Y(n_1787)
);

OAI322xp33_ASAP7_75t_L g1788 ( 
.A1(n_1731),
.A2(n_1725),
.A3(n_1715),
.B1(n_1678),
.B2(n_1706),
.C1(n_1714),
.C2(n_1699),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1744),
.A2(n_1624),
.B1(n_1611),
.B2(n_1645),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1756),
.A2(n_1719),
.B(n_1624),
.Y(n_1790)
);

AOI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1762),
.A2(n_1713),
.B(n_1712),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1770),
.Y(n_1792)
);

O2A1O1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1778),
.A2(n_1752),
.B(n_1744),
.C(n_1764),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1777),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1777),
.B(n_1735),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1784),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_SL g1797 ( 
.A1(n_1768),
.A2(n_1734),
.B(n_1743),
.C(n_1731),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1781),
.B(n_1738),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1766),
.B(n_1735),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1771),
.Y(n_1800)
);

OAI31xp33_ASAP7_75t_L g1801 ( 
.A1(n_1779),
.A2(n_1764),
.A3(n_1752),
.B(n_1744),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_L g1802 ( 
.A1(n_1776),
.A2(n_1745),
.B(n_1733),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1772),
.B(n_1763),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1773),
.A2(n_1752),
.B(n_1763),
.C(n_1742),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1788),
.A2(n_1790),
.B(n_1791),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1775),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1769),
.A2(n_1758),
.B1(n_1645),
.B2(n_1760),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1782),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1785),
.Y(n_1809)
);

XOR2x2_ASAP7_75t_L g1810 ( 
.A(n_1769),
.B(n_1524),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1783),
.A2(n_1643),
.B(n_1719),
.C(n_1636),
.Y(n_1811)
);

OAI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1802),
.A2(n_1786),
.B(n_1787),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1798),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1793),
.B(n_1767),
.C(n_1783),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1796),
.B(n_1780),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1796),
.B(n_1780),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1794),
.A2(n_1767),
.B1(n_1578),
.B2(n_1554),
.Y(n_1817)
);

AOI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1797),
.A2(n_1789),
.B1(n_1723),
.B2(n_1713),
.C(n_1716),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1803),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1803),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1795),
.B(n_1736),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1799),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1792),
.B(n_1738),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1805),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1817),
.B(n_1804),
.Y(n_1825)
);

NAND5xp2_ASAP7_75t_L g1826 ( 
.A(n_1813),
.B(n_1801),
.C(n_1807),
.D(n_1811),
.E(n_1808),
.Y(n_1826)
);

AND3x2_ASAP7_75t_L g1827 ( 
.A(n_1819),
.B(n_1520),
.C(n_1800),
.Y(n_1827)
);

NAND4xp25_ASAP7_75t_L g1828 ( 
.A(n_1815),
.B(n_1812),
.C(n_1822),
.D(n_1821),
.Y(n_1828)
);

NAND4xp25_ASAP7_75t_L g1829 ( 
.A(n_1823),
.B(n_1820),
.C(n_1814),
.D(n_1809),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1818),
.A2(n_1806),
.B1(n_1774),
.B2(n_1758),
.C(n_1676),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1823),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1813),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1816),
.B(n_1736),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1816),
.B(n_1739),
.Y(n_1834)
);

NOR2xp67_ASAP7_75t_SL g1835 ( 
.A(n_1815),
.B(n_1757),
.Y(n_1835)
);

OAI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1831),
.A2(n_1810),
.B1(n_1716),
.B2(n_1733),
.C(n_1676),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1833),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1835),
.A2(n_1676),
.B1(n_1541),
.B2(n_1678),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1826),
.A2(n_1829),
.B1(n_1824),
.B2(n_1825),
.C(n_1830),
.Y(n_1839)
);

AOI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1828),
.A2(n_1757),
.B(n_1541),
.C(n_1750),
.Y(n_1840)
);

AOI211xp5_ASAP7_75t_L g1841 ( 
.A1(n_1832),
.A2(n_1750),
.B(n_1739),
.C(n_1534),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1837),
.Y(n_1842)
);

NAND4xp25_ASAP7_75t_L g1843 ( 
.A(n_1839),
.B(n_1834),
.C(n_1827),
.D(n_1652),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1836),
.A2(n_1676),
.B(n_1679),
.C(n_1682),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1840),
.Y(n_1845)
);

AOI21xp33_ASAP7_75t_L g1846 ( 
.A1(n_1838),
.A2(n_1682),
.B(n_1679),
.Y(n_1846)
);

NAND4xp25_ASAP7_75t_SL g1847 ( 
.A(n_1841),
.B(n_1759),
.C(n_1753),
.D(n_1765),
.Y(n_1847)
);

XNOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1845),
.B(n_1534),
.Y(n_1848)
);

NAND4xp75_ASAP7_75t_L g1849 ( 
.A(n_1842),
.B(n_1759),
.C(n_1765),
.D(n_1588),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1847),
.Y(n_1850)
);

NOR2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1843),
.B(n_1534),
.Y(n_1851)
);

INVxp33_ASAP7_75t_L g1852 ( 
.A(n_1844),
.Y(n_1852)
);

NOR3xp33_ASAP7_75t_L g1853 ( 
.A(n_1850),
.B(n_1846),
.C(n_1682),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1852),
.B(n_1676),
.C(n_1700),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1848),
.A2(n_1707),
.B(n_1702),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1854),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1849),
.B1(n_1851),
.B2(n_1855),
.Y(n_1857)
);

NAND2x1p5_ASAP7_75t_L g1858 ( 
.A(n_1857),
.B(n_1530),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1857),
.B(n_1853),
.Y(n_1859)
);

NAND4xp75_ASAP7_75t_L g1860 ( 
.A(n_1859),
.B(n_1588),
.C(n_1685),
.D(n_1679),
.Y(n_1860)
);

OA21x2_ASAP7_75t_L g1861 ( 
.A1(n_1858),
.A2(n_1655),
.B(n_1656),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1861),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1860),
.B(n_1679),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1862),
.A2(n_1672),
.B1(n_1655),
.B2(n_1656),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1864),
.A2(n_1863),
.B(n_1685),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_R g1867 ( 
.A1(n_1866),
.A2(n_1652),
.B1(n_1621),
.B2(n_1681),
.C(n_1686),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1530),
.B(n_1537),
.C(n_1531),
.Y(n_1868)
);


endmodule