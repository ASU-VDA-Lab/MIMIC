module fake_jpeg_3194_n_419 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_419);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_419;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_57),
.Y(n_81)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_16),
.B1(n_19),
.B2(n_32),
.Y(n_88)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_0),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_31),
.B(n_13),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_38),
.Y(n_115)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_31),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_26),
.B1(n_33),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_107),
.B1(n_27),
.B2(n_30),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_64),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_88),
.A2(n_100),
.B1(n_107),
.B2(n_114),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_25),
.B1(n_33),
.B2(n_23),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_95),
.B1(n_98),
.B2(n_105),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_41),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_39),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_50),
.A2(n_36),
.B1(n_33),
.B2(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_25),
.B1(n_22),
.B2(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_17),
.B1(n_47),
.B2(n_65),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_43),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_17),
.B1(n_61),
.B2(n_63),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_52),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_38),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_17),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_123),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_149),
.B1(n_78),
.B2(n_91),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_133),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_58),
.B(n_60),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_98),
.B(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_128),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_64),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_138),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_132),
.A2(n_154),
.B1(n_125),
.B2(n_134),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_70),
.C(n_45),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_106),
.C(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_137),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_142),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_54),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_68),
.B1(n_28),
.B2(n_2),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_111),
.B(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_153),
.Y(n_161)
);

BUFx8_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_75),
.B(n_13),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_87),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_159),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_77),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_162),
.A2(n_174),
.B(n_181),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_169),
.B1(n_175),
.B2(n_142),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_133),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_101),
.B(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_113),
.B1(n_96),
.B2(n_91),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_77),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_191),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_118),
.A2(n_113),
.B(n_96),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_103),
.C(n_104),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_194),
.C(n_198),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_126),
.A2(n_103),
.B(n_104),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_145),
.B(n_152),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_1),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_28),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_124),
.A2(n_28),
.B1(n_12),
.B2(n_4),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_28),
.C(n_3),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_201),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_202),
.A2(n_208),
.B1(n_213),
.B2(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_204),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_152),
.B(n_147),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_205),
.A2(n_230),
.B(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_165),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_143),
.B1(n_150),
.B2(n_130),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_186),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_143),
.B1(n_136),
.B2(n_144),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_143),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_129),
.Y(n_219)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_143),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_161),
.A2(n_158),
.B(n_146),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_222),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_137),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_225),
.Y(n_261)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_121),
.B1(n_148),
.B2(n_120),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_173),
.A2(n_139),
.B1(n_122),
.B2(n_5),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_168),
.B1(n_173),
.B2(n_160),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_2),
.B(n_4),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_4),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_198),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_168),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_194),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_172),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_178),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_179),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_252),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_170),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_250),
.C(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_269),
.B1(n_213),
.B2(n_208),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_187),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_161),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_173),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_172),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_266),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_174),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_220),
.Y(n_266)
);

OAI22x1_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_181),
.B1(n_197),
.B2(n_195),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_227),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_202),
.A2(n_164),
.B1(n_178),
.B2(n_180),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_205),
.B(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_223),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_273),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_278),
.B1(n_279),
.B2(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_215),
.B1(n_214),
.B2(n_230),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_249),
.A2(n_214),
.B1(n_231),
.B2(n_215),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_282),
.A2(n_286),
.B1(n_296),
.B2(n_299),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_225),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_288),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_231),
.B1(n_227),
.B2(n_228),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_290),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_246),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_229),
.B1(n_227),
.B2(n_200),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_246),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_240),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_238),
.A2(n_206),
.B1(n_201),
.B2(n_177),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_300),
.C(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_184),
.C(n_193),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_271),
.B1(n_261),
.B2(n_265),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_307),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_238),
.B1(n_255),
.B2(n_259),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_308),
.B1(n_320),
.B2(n_326),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_247),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_299),
.A2(n_255),
.B1(n_254),
.B2(n_244),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_260),
.C(n_248),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_314),
.C(n_317),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_242),
.C(n_252),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_254),
.C(n_270),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_257),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_327),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_279),
.A2(n_257),
.B1(n_268),
.B2(n_265),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_241),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_322),
.C(n_180),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_271),
.C(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_292),
.A2(n_265),
.B1(n_261),
.B2(n_218),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_193),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_276),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_329),
.B(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_280),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_274),
.B(n_273),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_340),
.B(n_317),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_286),
.B1(n_282),
.B2(n_289),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_338),
.B1(n_347),
.B2(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_294),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_335),
.B(n_336),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_323),
.A2(n_301),
.B1(n_291),
.B2(n_280),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_283),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_8),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_296),
.B1(n_281),
.B2(n_277),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_293),
.B(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_284),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_343),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_183),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_183),
.B1(n_6),
.B2(n_7),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_340),
.B1(n_349),
.B2(n_319),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_320),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_5),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_313),
.C(n_304),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_351),
.B(n_365),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_355),
.A2(n_333),
.B(n_338),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_318),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_358),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_305),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_334),
.A2(n_324),
.B1(n_311),
.B2(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_331),
.A2(n_326),
.B1(n_325),
.B2(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_349),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_346),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_366),
.B(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_372),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_369),
.A2(n_361),
.B1(n_352),
.B2(n_365),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_345),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_376),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_375),
.A2(n_355),
.B(n_367),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_353),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_342),
.C(n_330),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_378),
.B(n_379),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_342),
.C(n_330),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_385),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_380),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_358),
.C(n_357),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_386),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_360),
.C(n_354),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_388),
.C(n_375),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_354),
.C(n_352),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_377),
.B1(n_8),
.B2(n_11),
.Y(n_402)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_397),
.Y(n_407)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_396),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_387),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_370),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_401),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_369),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_402),
.Y(n_409)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_391),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_SL g404 ( 
.A(n_394),
.B(n_384),
.C(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_383),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_408),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_386),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_395),
.B(n_396),
.Y(n_410)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_400),
.C(n_385),
.Y(n_413)
);

O2A1O1Ixp33_ASAP7_75t_SL g414 ( 
.A1(n_413),
.A2(n_406),
.B(n_404),
.C(n_409),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_416),
.A2(n_412),
.B(n_415),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_417),
.A2(n_411),
.B(n_11),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_11),
.Y(n_419)
);


endmodule