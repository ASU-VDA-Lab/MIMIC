module real_jpeg_6555_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_32;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_5),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_24),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_3),
.A2(n_4),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g12 ( 
.A1(n_4),
.A2(n_13),
.B(n_14),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OR2x2_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_31),
.Y(n_7)
);

OAI22xp33_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_10),
.A2(n_27),
.B1(n_32),
.B2(n_34),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_12),
.B(n_15),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_19),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OR2x4_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);


endmodule