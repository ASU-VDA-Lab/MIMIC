module real_aes_7136_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1170;
wire n_1175;
wire n_1106;
wire n_778;
wire n_522;
wire n_800;
wire n_838;
wire n_933;
wire n_1092;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_448;
wire n_556;
wire n_545;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_958;
wire n_677;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_1140;
wire n_510;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_976;
wire n_1182;
wire n_636;
wire n_1053;
wire n_1049;
wire n_559;
wire n_477;
wire n_872;
wire n_515;
wire n_906;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1168;
wire n_1025;
wire n_755;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_725;
wire n_504;
wire n_973;
wire n_671;
wire n_1084;
wire n_960;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1135;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_1167;
wire n_1174;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1037;
wire n_1103;
wire n_1131;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_1179;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_810;
wire n_1079;
wire n_843;
wire n_1136;
wire n_579;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_1033;
wire n_1187;
wire n_727;
wire n_1014;
wire n_649;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_922;
wire n_926;
wire n_679;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1114;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_1156;
wire n_474;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_597;
wire n_1176;
wire n_483;
wire n_611;
wire n_640;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1101;
wire n_1076;
wire n_661;
wire n_463;
wire n_396;
wire n_1102;
wire n_804;
wire n_447;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_0), .A2(n_56), .B1(n_633), .B2(n_989), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g1060 ( .A1(n_1), .A2(n_295), .B1(n_482), .B2(n_649), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_2), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_3), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_4), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_5), .A2(n_51), .B1(n_571), .B2(n_574), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_6), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_7), .A2(n_14), .B1(n_423), .B2(n_528), .C(n_530), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_8), .A2(n_278), .B1(n_460), .B2(n_505), .C(n_506), .Y(n_504) );
AOI22x1_ASAP7_75t_L g695 ( .A1(n_9), .A2(n_696), .B1(n_731), .B2(n_732), .Y(n_695) );
INVx1_ASAP7_75t_L g731 ( .A(n_9), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_10), .A2(n_139), .B1(n_680), .B2(n_907), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_11), .Y(n_792) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_12), .A2(n_226), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g1148 ( .A(n_12), .Y(n_1148) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_13), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_15), .A2(n_300), .B1(n_607), .B2(n_964), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_16), .A2(n_95), .B1(n_495), .B2(n_651), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_17), .Y(n_973) );
AOI222xp33_ASAP7_75t_L g990 ( .A1(n_18), .A2(n_52), .B1(n_153), .B2(n_401), .C1(n_574), .C2(n_639), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_19), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_20), .A2(n_251), .B1(n_760), .B2(n_761), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_21), .A2(n_161), .B1(n_573), .B2(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_22), .B(n_726), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_23), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_24), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_25), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_26), .A2(n_365), .B1(n_597), .B2(n_746), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_27), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_28), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_29), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_30), .A2(n_124), .B1(n_807), .B2(n_808), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_31), .Y(n_1006) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_32), .A2(n_106), .B1(n_404), .B2(n_408), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_33), .A2(n_503), .B1(n_546), .B2(n_547), .Y(n_502) );
INVx1_ASAP7_75t_L g546 ( .A(n_33), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_34), .A2(n_376), .B1(n_603), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_35), .A2(n_213), .B1(n_476), .B2(n_604), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_36), .A2(n_855), .B1(n_885), .B2(n_886), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_36), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_37), .A2(n_111), .B1(n_462), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_38), .A2(n_53), .B1(n_484), .B2(n_761), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_39), .A2(n_166), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_40), .A2(n_285), .B1(n_810), .B2(n_907), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g1102 ( .A(n_41), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_42), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_43), .B(n_528), .Y(n_637) );
AOI22xp5_ASAP7_75t_SL g1063 ( .A1(n_44), .A2(n_1064), .B1(n_1065), .B2(n_1084), .Y(n_1063) );
INVx1_ASAP7_75t_L g1084 ( .A(n_44), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_45), .A2(n_196), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_46), .A2(n_304), .B1(n_454), .B2(n_592), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g1134 ( .A1(n_47), .A2(n_221), .B1(n_445), .B2(n_454), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_48), .A2(n_249), .B1(n_556), .B2(n_1079), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_49), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_50), .B(n_424), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g1168 ( .A(n_54), .Y(n_1168) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_55), .A2(n_381), .B1(n_683), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_57), .A2(n_296), .B1(n_518), .B2(n_1114), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_58), .A2(n_1152), .B1(n_1176), .B2(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_58), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_59), .A2(n_131), .B1(n_709), .B2(n_711), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_60), .B(n_726), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_61), .A2(n_328), .B1(n_512), .B2(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_62), .A2(n_1095), .B1(n_1116), .B2(n_1117), .Y(n_1094) );
INVx1_ASAP7_75t_L g1116 ( .A(n_62), .Y(n_1116) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_63), .A2(n_281), .B1(n_472), .B2(n_785), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_64), .Y(n_925) );
INVx1_ASAP7_75t_L g671 ( .A(n_65), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_66), .A2(n_191), .B1(n_680), .B2(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_67), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_68), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_69), .A2(n_100), .B1(n_631), .B2(n_808), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_70), .A2(n_345), .B1(n_558), .B2(n_683), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_71), .Y(n_415) );
INVx1_ASAP7_75t_L g986 ( .A(n_72), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_73), .A2(n_96), .B1(n_470), .B2(n_1011), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_74), .A2(n_255), .B1(n_430), .B2(n_435), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_75), .A2(n_264), .B1(n_454), .B2(n_592), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_76), .A2(n_323), .B1(n_591), .B2(n_639), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_77), .A2(n_217), .B1(n_591), .B2(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_78), .Y(n_877) );
INVx1_ASAP7_75t_L g1120 ( .A(n_79), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_80), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_81), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_82), .A2(n_134), .B1(n_581), .B2(n_582), .Y(n_580) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_83), .A2(n_256), .B1(n_404), .B2(n_405), .Y(n_413) );
INVx1_ASAP7_75t_L g1145 ( .A(n_83), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_84), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_85), .A2(n_86), .B1(n_607), .B2(n_681), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_87), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_88), .A2(n_104), .B1(n_613), .B2(n_931), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_89), .A2(n_232), .B1(n_455), .B2(n_592), .Y(n_1050) );
OA22x2_ASAP7_75t_L g944 ( .A1(n_90), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_90), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_91), .A2(n_152), .B1(n_470), .B2(n_476), .Y(n_469) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_92), .A2(n_101), .B1(n_138), .B2(n_444), .C1(n_543), .C2(n_545), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_93), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g1174 ( .A(n_94), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_97), .A2(n_145), .B1(n_435), .B2(n_452), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_98), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_99), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_102), .A2(n_219), .B1(n_760), .B2(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g1075 ( .A1(n_103), .A2(n_363), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_105), .A2(n_155), .B1(n_492), .B2(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g1149 ( .A(n_106), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_107), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_108), .A2(n_172), .B1(n_600), .B2(n_958), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_109), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_110), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_112), .A2(n_223), .B1(n_785), .B2(n_814), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g1049 ( .A(n_113), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_114), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_115), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_116), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_117), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_118), .A2(n_299), .B1(n_496), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_119), .A2(n_279), .B1(n_680), .B2(n_1076), .Y(n_1159) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_120), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_121), .A2(n_320), .B1(n_460), .B2(n_465), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_122), .A2(n_229), .B1(n_558), .B2(n_711), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_123), .A2(n_136), .B1(n_505), .B2(n_611), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_125), .A2(n_239), .B1(n_424), .B2(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_126), .A2(n_316), .B1(n_468), .B2(n_808), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_127), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_128), .B(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_129), .A2(n_183), .B1(n_573), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_130), .A2(n_311), .B1(n_607), .B2(n_608), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_132), .A2(n_179), .B1(n_555), .B2(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_133), .A2(n_340), .B1(n_455), .B2(n_600), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_135), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_137), .A2(n_336), .B1(n_592), .B2(n_775), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_140), .A2(n_200), .B1(n_430), .B2(n_633), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_141), .A2(n_319), .B1(n_643), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_142), .A2(n_321), .B1(n_760), .B2(n_761), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_143), .A2(n_210), .B1(n_651), .B2(n_652), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g1129 ( .A(n_144), .Y(n_1129) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_146), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_147), .B(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_148), .A2(n_208), .B1(n_810), .B2(n_811), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_149), .A2(n_244), .B1(n_646), .B2(n_980), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_150), .Y(n_397) );
AND2x6_ASAP7_75t_L g388 ( .A(n_151), .B(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_151), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g749 ( .A1(n_154), .A2(n_175), .B1(n_681), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_156), .A2(n_241), .B1(n_680), .B2(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_157), .A2(n_286), .B1(n_435), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_158), .A2(n_181), .B1(n_710), .B2(n_780), .Y(n_933) );
INVx1_ASAP7_75t_L g837 ( .A(n_159), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_160), .A2(n_268), .B1(n_670), .B2(n_931), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_162), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_163), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_164), .A2(n_266), .B1(n_484), .B2(n_863), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_165), .A2(n_189), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp5_ASAP7_75t_SL g654 ( .A1(n_167), .A2(n_655), .B1(n_692), .B2(n_693), .Y(n_654) );
INVx1_ASAP7_75t_L g693 ( .A(n_167), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_168), .A2(n_290), .B1(n_454), .B2(n_639), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g1124 ( .A1(n_169), .A2(n_315), .B1(n_652), .B2(n_710), .Y(n_1124) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_170), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g658 ( .A(n_171), .Y(n_658) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_173), .A2(n_245), .B1(n_404), .B2(n_408), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_173), .B(n_1147), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_174), .B(n_1170), .Y(n_1169) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_176), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_177), .A2(n_263), .B1(n_556), .B2(n_616), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_178), .Y(n_493) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_180), .A2(n_400), .B(n_414), .C(n_441), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_182), .A2(n_274), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_184), .A2(n_190), .B1(n_686), .B2(n_908), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_185), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_186), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_187), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_188), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_192), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_193), .A2(n_228), .B1(n_466), .B2(n_613), .Y(n_778) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_194), .A2(n_207), .B1(n_611), .B2(n_613), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g1127 ( .A1(n_195), .A2(n_234), .B1(n_607), .B2(n_910), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_197), .A2(n_230), .B1(n_581), .B2(n_582), .Y(n_1072) );
AOI22xp33_ASAP7_75t_SL g1081 ( .A1(n_198), .A2(n_366), .B1(n_863), .B2(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1068 ( .A(n_199), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_201), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_202), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_203), .A2(n_382), .B1(n_466), .B2(n_492), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_204), .B(n_880), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_205), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_206), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_209), .A2(n_303), .B1(n_687), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_211), .A2(n_310), .B1(n_472), .B2(n_484), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_212), .A2(n_360), .B1(n_603), .B2(n_604), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_214), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_215), .A2(n_260), .B1(n_780), .B2(n_808), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_216), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_218), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_220), .A2(n_225), .B1(n_591), .B2(n_1002), .Y(n_1001) );
XNOR2x2_ASAP7_75t_L g975 ( .A(n_222), .B(n_976), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_224), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_227), .A2(n_350), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_231), .A2(n_334), .B1(n_607), .B2(n_964), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_233), .A2(n_280), .B1(n_689), .B2(n_690), .Y(n_688) );
OA22x2_ASAP7_75t_L g912 ( .A1(n_235), .A2(n_913), .B1(n_914), .B2(n_935), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_235), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_236), .A2(n_375), .B1(n_512), .B2(n_754), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_237), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_238), .B(n_595), .Y(n_594) );
XNOR2x2_ASAP7_75t_L g550 ( .A(n_240), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_242), .A2(n_369), .B1(n_460), .B2(n_910), .Y(n_1032) );
INVx2_ASAP7_75t_L g392 ( .A(n_243), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_246), .A2(n_258), .B1(n_518), .B2(n_807), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_247), .B(n_582), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g1167 ( .A(n_248), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_250), .A2(n_282), .B1(n_430), .B2(n_438), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_252), .A2(n_378), .B1(n_492), .B2(n_910), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_253), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_254), .A2(n_373), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_257), .A2(n_352), .B1(n_431), .B2(n_639), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_259), .A2(n_384), .B(n_393), .C(n_1150), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_261), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_262), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_265), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_267), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_269), .A2(n_314), .B1(n_484), .B2(n_761), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_270), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_271), .A2(n_370), .B1(n_604), .B2(n_683), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_272), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_273), .A2(n_374), .B1(n_616), .B2(n_811), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_275), .A2(n_357), .B1(n_512), .B2(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_276), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_277), .Y(n_917) );
OA22x2_ASAP7_75t_L g736 ( .A1(n_283), .A2(n_737), .B1(n_738), .B2(n_762), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_283), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_284), .B(n_598), .Y(n_987) );
OA22x2_ASAP7_75t_L g1018 ( .A1(n_287), .A2(n_1019), .B1(n_1020), .B2(n_1037), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_287), .Y(n_1019) );
INVx1_ASAP7_75t_L g668 ( .A(n_288), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_289), .A2(n_312), .B1(n_608), .B2(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g674 ( .A(n_291), .Y(n_674) );
INVx1_ASAP7_75t_L g404 ( .A(n_292), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_292), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_293), .A2(n_372), .B1(n_808), .B2(n_931), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_294), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_297), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g1052 ( .A(n_298), .Y(n_1052) );
CKINVDCx20_ASAP7_75t_R g1164 ( .A(n_301), .Y(n_1164) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_302), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_305), .A2(n_322), .B1(n_515), .B2(n_518), .C(n_521), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_306), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_307), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_308), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_309), .Y(n_1023) );
INVx1_ASAP7_75t_L g1163 ( .A(n_313), .Y(n_1163) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_317), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_318), .A2(n_367), .B1(n_482), .B2(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_324), .A2(n_359), .B1(n_780), .B2(n_910), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_325), .A2(n_344), .B1(n_431), .B2(n_437), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g1151 ( .A1(n_326), .A2(n_1152), .B1(n_1175), .B2(n_1176), .Y(n_1151) );
CKINVDCx20_ASAP7_75t_R g1175 ( .A(n_326), .Y(n_1175) );
INVx1_ASAP7_75t_L g391 ( .A(n_327), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_329), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_330), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_331), .Y(n_617) );
INVx1_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_333), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_335), .Y(n_522) );
OA22x2_ASAP7_75t_L g888 ( .A1(n_337), .A2(n_889), .B1(n_890), .B2(n_911), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_337), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_338), .A2(n_364), .B1(n_680), .B2(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_339), .B(n_598), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_341), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_342), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_343), .B(n_574), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_346), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_347), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_348), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_349), .Y(n_833) );
INVx1_ASAP7_75t_L g1015 ( .A(n_351), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g1098 ( .A(n_353), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_354), .B(n_435), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g1173 ( .A(n_355), .Y(n_1173) );
INVx1_ASAP7_75t_L g663 ( .A(n_356), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_358), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_361), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_362), .Y(n_707) );
INVx1_ASAP7_75t_L g1062 ( .A(n_368), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_371), .Y(n_653) );
OA22x2_ASAP7_75t_SL g822 ( .A1(n_377), .A2(n_823), .B1(n_824), .B2(n_847), .Y(n_822) );
INVx1_ASAP7_75t_L g847 ( .A(n_377), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_379), .Y(n_1105) );
INVx1_ASAP7_75t_L g675 ( .A(n_380), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_389), .Y(n_1141) );
OAI21xp5_ASAP7_75t_L g1187 ( .A1(n_390), .A2(n_1140), .B(n_1188), .Y(n_1187) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_851), .B1(n_1135), .B2(n_1136), .C(n_1137), .Y(n_393) );
INVx1_ASAP7_75t_L g1135 ( .A(n_394), .Y(n_1135) );
XOR2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_499), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
XNOR2x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_457), .Y(n_398) );
INVx3_ASAP7_75t_L g893 ( .A(n_400), .Y(n_893) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx4_ASAP7_75t_L g544 ( .A(n_401), .Y(n_544) );
INVx2_ASAP7_75t_L g568 ( .A(n_401), .Y(n_568) );
INVx2_ASAP7_75t_L g588 ( .A(n_401), .Y(n_588) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_401), .Y(n_631) );
INVx2_ASAP7_75t_SL g1166 ( .A(n_401), .Y(n_1166) );
AND2x6_ASAP7_75t_L g401 ( .A(n_402), .B(n_409), .Y(n_401) );
AND2x4_ASAP7_75t_L g438 ( .A(n_402), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g540 ( .A(n_402), .Y(n_540) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .Y(n_402) );
INVx2_ASAP7_75t_L g420 ( .A(n_403), .Y(n_420) );
AND2x2_ASAP7_75t_L g434 ( .A(n_403), .B(n_411), .Y(n_434) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_406), .Y(n_408) );
AND2x2_ASAP7_75t_L g419 ( .A(n_407), .B(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g428 ( .A(n_407), .B(n_420), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVx2_ASAP7_75t_L g449 ( .A(n_407), .Y(n_449) );
AND2x2_ASAP7_75t_L g463 ( .A(n_409), .B(n_464), .Y(n_463) );
AND2x6_ASAP7_75t_L g468 ( .A(n_409), .B(n_427), .Y(n_468) );
AND2x4_ASAP7_75t_L g484 ( .A(n_409), .B(n_419), .Y(n_484) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
AND2x2_ASAP7_75t_L g421 ( .A(n_410), .B(n_413), .Y(n_421) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g475 ( .A(n_411), .B(n_440), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_411), .B(n_413), .Y(n_478) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
INVx1_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_422), .C(n_429), .Y(n_414) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g720 ( .A(n_417), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_417), .A2(n_661), .B1(n_1129), .B2(n_1130), .C(n_1131), .Y(n_1128) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g665 ( .A(n_418), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x2_ASAP7_75t_L g474 ( .A(n_419), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_419), .B(n_475), .Y(n_509) );
AND2x6_ASAP7_75t_L g529 ( .A(n_419), .B(n_421), .Y(n_529) );
AND2x2_ASAP7_75t_L g464 ( .A(n_420), .B(n_449), .Y(n_464) );
AND2x4_ASAP7_75t_L g426 ( .A(n_421), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g492 ( .A(n_421), .B(n_464), .Y(n_492) );
INVx1_ASAP7_75t_L g662 ( .A(n_421), .Y(n_662) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g581 ( .A(n_425), .Y(n_581) );
INVx5_ASAP7_75t_L g598 ( .A(n_425), .Y(n_598) );
INVx2_ASAP7_75t_L g636 ( .A(n_425), .Y(n_636) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g661 ( .A(n_428), .B(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g579 ( .A(n_431), .Y(n_579) );
BUFx2_ASAP7_75t_L g600 ( .A(n_431), .Y(n_600) );
BUFx3_ASAP7_75t_L g775 ( .A(n_431), .Y(n_775) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g477 ( .A(n_433), .B(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g446 ( .A(n_434), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g455 ( .A(n_434), .B(n_456), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_434), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_SL g592 ( .A(n_438), .Y(n_592) );
BUFx2_ASAP7_75t_SL g633 ( .A(n_438), .Y(n_633) );
INVx1_ASAP7_75t_L g541 ( .A(n_439), .Y(n_541) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_450), .B2(n_451), .Y(n_441) );
OAI222xp33_ASAP7_75t_L g721 ( .A1(n_443), .A2(n_722), .B1(n_723), .B2(n_724), .C1(n_725), .C2(n_727), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_443), .A2(n_667), .B1(n_877), .B2(n_878), .C(n_879), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_443), .A2(n_1166), .B1(n_1167), .B2(n_1168), .C(n_1169), .Y(n_1165) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g1053 ( .A(n_444), .Y(n_1053) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g801 ( .A(n_445), .Y(n_801) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_446), .Y(n_573) );
BUFx4f_ASAP7_75t_SL g639 ( .A(n_446), .Y(n_639) );
BUFx2_ASAP7_75t_L g670 ( .A(n_446), .Y(n_670) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_446), .Y(n_958) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g456 ( .A(n_448), .Y(n_456) );
INVx1_ASAP7_75t_L g535 ( .A(n_449), .Y(n_535) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx4f_ASAP7_75t_SL g545 ( .A(n_454), .Y(n_545) );
BUFx12f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_455), .Y(n_575) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_455), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_479), .C(n_489), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .Y(n_458) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_461), .A2(n_699), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_698) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_462), .Y(n_555) );
BUFx3_ASAP7_75t_L g680 ( .A(n_462), .Y(n_680) );
BUFx3_ASAP7_75t_L g859 ( .A(n_462), .Y(n_859) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_463), .Y(n_616) );
INVx2_ASAP7_75t_L g781 ( .A(n_463), .Y(n_781) );
BUFx2_ASAP7_75t_SL g1079 ( .A(n_463), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_464), .B(n_475), .Y(n_488) );
AND2x4_ASAP7_75t_L g497 ( .A(n_464), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g614 ( .A(n_464), .B(n_475), .Y(n_614) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g561 ( .A(n_466), .Y(n_561) );
INVx5_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g517 ( .A(n_467), .Y(n_517) );
INVx4_ASAP7_75t_L g643 ( .A(n_467), .Y(n_643) );
INVx2_ASAP7_75t_L g686 ( .A(n_467), .Y(n_686) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_467), .Y(n_751) );
INVx1_ASAP7_75t_L g860 ( .A(n_467), .Y(n_860) );
INVx11_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx11_ASAP7_75t_L g612 ( .A(n_468), .Y(n_612) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_472), .Y(n_558) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g605 ( .A(n_473), .Y(n_605) );
INVx3_ASAP7_75t_L g649 ( .A(n_473), .Y(n_649) );
INVx5_ASAP7_75t_L g710 ( .A(n_473), .Y(n_710) );
INVx2_ASAP7_75t_L g754 ( .A(n_473), .Y(n_754) );
INVx1_ASAP7_75t_L g863 ( .A(n_473), .Y(n_863) );
INVx8_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx6_ASAP7_75t_SL g513 ( .A(n_477), .Y(n_513) );
INVx1_ASAP7_75t_SL g785 ( .A(n_477), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_477), .A2(n_539), .B1(n_925), .B2(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g1011 ( .A(n_477), .Y(n_1011) );
INVx1_ASAP7_75t_L g498 ( .A(n_478), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_485), .B2(n_486), .Y(n_479) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_483), .A2(n_526), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g603 ( .A(n_483), .Y(n_603) );
INVx3_ASAP7_75t_L g908 ( .A(n_483), .Y(n_908) );
INVx2_ASAP7_75t_L g1082 ( .A(n_483), .Y(n_1082) );
INVx6_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g524 ( .A(n_484), .Y(n_524) );
BUFx3_ASAP7_75t_L g760 ( .A(n_484), .Y(n_760) );
BUFx3_ASAP7_75t_L g931 ( .A(n_484), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_486), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g526 ( .A(n_487), .Y(n_526) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_493), .B2(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g651 ( .A(n_491), .Y(n_651) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_492), .Y(n_520) );
BUFx3_ASAP7_75t_L g607 ( .A(n_492), .Y(n_607) );
BUFx3_ASAP7_75t_L g687 ( .A(n_492), .Y(n_687) );
BUFx3_ASAP7_75t_L g816 ( .A(n_492), .Y(n_816) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx3_ASAP7_75t_L g505 ( .A(n_497), .Y(n_505) );
BUFx2_ASAP7_75t_SL g556 ( .A(n_497), .Y(n_556) );
BUFx3_ASAP7_75t_L g646 ( .A(n_497), .Y(n_646) );
BUFx3_ASAP7_75t_L g681 ( .A(n_497), .Y(n_681) );
BUFx2_ASAP7_75t_SL g811 ( .A(n_497), .Y(n_811) );
BUFx2_ASAP7_75t_L g910 ( .A(n_497), .Y(n_910) );
AND2x2_ASAP7_75t_L g652 ( .A(n_498), .B(n_535), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_619), .B1(n_849), .B2(n_850), .Y(n_499) );
INVx1_ASAP7_75t_L g849 ( .A(n_500), .Y(n_849) );
OAI22xp5_ASAP7_75t_SL g500 ( .A1(n_501), .A2(n_502), .B1(n_548), .B2(n_618), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g547 ( .A(n_503), .Y(n_547) );
AND4x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .C(n_527), .D(n_542), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_510), .B2(n_511), .Y(n_506) );
BUFx2_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g608 ( .A(n_513), .Y(n_608) );
BUFx2_ASAP7_75t_L g683 ( .A(n_513), .Y(n_683) );
BUFx4f_ASAP7_75t_SL g711 ( .A(n_513), .Y(n_711) );
BUFx2_ASAP7_75t_L g964 ( .A(n_513), .Y(n_964) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_519), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_559) );
INVx3_ASAP7_75t_L g980 ( .A(n_519), .Y(n_980) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_525), .B2(n_526), .Y(n_521) );
INVx2_ASAP7_75t_L g689 ( .A(n_523), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_523), .A2(n_526), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_526), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
BUFx4f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g582 ( .A(n_529), .Y(n_582) );
BUFx2_ASAP7_75t_L g595 ( .A(n_529), .Y(n_595) );
INVx1_ASAP7_75t_SL g747 ( .A(n_529), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_536), .B2(n_537), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_532), .A2(n_537), .B1(n_729), .B2(n_730), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_532), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_532), .A2(n_537), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_SL g1005 ( .A(n_533), .Y(n_1005) );
INVx4_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_534), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
BUFx3_ASAP7_75t_L g803 ( .A(n_534), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_534), .A2(n_676), .B1(n_874), .B2(n_875), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_534), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_537), .A2(n_1005), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g676 ( .A(n_538), .Y(n_676) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g838 ( .A(n_539), .Y(n_838) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g667 ( .A(n_543), .Y(n_667) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_544), .Y(n_1000) );
OAI21xp5_ASAP7_75t_SL g1048 ( .A1(n_544), .A2(n_1049), .B(n_1050), .Y(n_1048) );
INVx2_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_583), .B2(n_584), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_552), .B(n_566), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_559), .C(n_563), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_576), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_569), .B(n_570), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_568), .A2(n_741), .B(n_742), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g768 ( .A1(n_568), .A2(n_769), .B(n_770), .Y(n_768) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx4_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g832 ( .A(n_573), .Y(n_832) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_573), .Y(n_1002) );
INVx1_ASAP7_75t_L g1025 ( .A(n_574), .Y(n_1025) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g793 ( .A(n_575), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g989 ( .A(n_579), .Y(n_989) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
XOR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_617), .Y(n_584) );
NAND3x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_601), .C(n_609), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_593), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_590), .Y(n_587) );
BUFx3_ASAP7_75t_L g726 ( .A(n_591), .Y(n_726) );
BUFx2_ASAP7_75t_L g880 ( .A(n_591), .Y(n_880) );
INVx2_ASAP7_75t_L g1171 ( .A(n_591), .Y(n_1171) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .C(n_599), .Y(n_593) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_606), .Y(n_601) );
INVx2_ASAP7_75t_L g866 ( .A(n_603), .Y(n_866) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_607), .Y(n_701) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
INVx4_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g807 ( .A(n_612), .Y(n_807) );
INVx4_ASAP7_75t_L g907 ( .A(n_612), .Y(n_907) );
OAI21xp33_ASAP7_75t_SL g921 ( .A1(n_612), .A2(n_922), .B(n_923), .Y(n_921) );
INVx3_ASAP7_75t_L g1076 ( .A(n_612), .Y(n_1076) );
BUFx3_ASAP7_75t_L g761 ( .A(n_613), .Y(n_761) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx3_ASAP7_75t_L g644 ( .A(n_614), .Y(n_644) );
BUFx3_ASAP7_75t_L g808 ( .A(n_614), .Y(n_808) );
BUFx3_ASAP7_75t_L g983 ( .A(n_614), .Y(n_983) );
INVx1_ASAP7_75t_L g967 ( .A(n_616), .Y(n_967) );
INVx1_ASAP7_75t_L g850 ( .A(n_619), .Y(n_850) );
XOR2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_733), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_694), .B2(n_695), .Y(n_620) );
INVx4_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_654), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI22x1_ASAP7_75t_L g821 ( .A1(n_624), .A2(n_625), .B1(n_765), .B2(n_818), .Y(n_821) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
XOR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_653), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_627), .B(n_640), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_634), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_632), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_630), .A2(n_792), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_791) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g723 ( .A(n_631), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .C(n_638), .Y(n_634) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_647), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g691 ( .A(n_644), .Y(n_691) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_646), .Y(n_704) );
INVx2_ASAP7_75t_L g1115 ( .A(n_646), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_SL g692 ( .A(n_655), .Y(n_692) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_656), .B(n_677), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_666), .C(n_673), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_663), .B2(n_664), .Y(n_657) );
OAI22xp5_ASAP7_75t_SL g949 ( .A1(n_659), .A2(n_719), .B1(n_950), .B2(n_951), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_659), .A2(n_719), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g828 ( .A(n_660), .Y(n_828) );
INVx1_ASAP7_75t_SL g996 ( .A(n_660), .Y(n_996) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_661), .Y(n_717) );
BUFx3_ASAP7_75t_L g918 ( .A(n_661), .Y(n_918) );
OA211x2_ASAP7_75t_L g985 ( .A1(n_664), .A2(n_986), .B(n_987), .C(n_988), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_664), .A2(n_918), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g884 ( .A(n_665), .Y(n_884) );
INVx1_ASAP7_75t_SL g920 ( .A(n_665), .Y(n_920) );
OAI221xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_671), .C(n_672), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g830 ( .A1(n_667), .A2(n_831), .B1(n_832), .B2(n_833), .C(n_834), .Y(n_830) );
OAI21xp5_ASAP7_75t_SL g1067 ( .A1(n_667), .A2(n_1068), .B(n_1069), .Y(n_1067) );
OAI221xp5_ASAP7_75t_SL g1100 ( .A1(n_667), .A2(n_957), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_676), .A2(n_1004), .B1(n_1005), .B2(n_1006), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_684), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_682), .Y(n_678) );
INVxp67_ASAP7_75t_L g871 ( .A(n_681), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g758 ( .A(n_687), .Y(n_758) );
BUFx2_ASAP7_75t_L g842 ( .A(n_687), .Y(n_842) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g732 ( .A(n_696), .Y(n_732) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_697), .B(n_712), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_710), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_721), .C(n_728), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_718), .B2(n_719), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_715), .A2(n_719), .B1(n_797), .B2(n_798), .Y(n_796) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_717), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_719), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_719), .A2(n_995), .B1(n_996), .B2(n_997), .Y(n_994) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI222xp33_ASAP7_75t_L g1022 ( .A1(n_723), .A2(n_832), .B1(n_1023), .B2(n_1024), .C1(n_1025), .C2(n_1026), .Y(n_1022) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_819), .B1(n_820), .B2(n_848), .Y(n_733) );
INVx1_ASAP7_75t_L g848 ( .A(n_734), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_763), .B2(n_764), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g762 ( .A(n_738), .Y(n_762) );
NAND3x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_748), .C(n_755), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g898 ( .A(n_747), .Y(n_898) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_758), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_868) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
AO22x2_ASAP7_75t_SL g764 ( .A1(n_765), .A2(n_787), .B1(n_788), .B2(n_818), .Y(n_764) );
INVx3_ASAP7_75t_L g818 ( .A(n_765), .Y(n_818) );
XOR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_786), .Y(n_765) );
NAND2x1_ASAP7_75t_SL g766 ( .A(n_767), .B(n_776), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .C(n_774), .Y(n_771) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_782), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx3_ASAP7_75t_L g810 ( .A(n_781), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
XOR2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_817), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_804), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_796), .C(n_799), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_803), .A2(n_956), .B1(n_957), .B2(n_959), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_812), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_808), .Y(n_1156) );
INVx1_ASAP7_75t_SL g969 ( .A(n_811), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
INVx2_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
XNOR2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_SL g824 ( .A(n_825), .B(n_839), .Y(n_824) );
NOR3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_830), .C(n_835), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g1162 ( .A1(n_828), .A2(n_920), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_841), .B(n_843), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g1136 ( .A(n_851), .Y(n_1136) );
XOR2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_1091), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_938), .B1(n_1089), .B2(n_1090), .Y(n_852) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_853), .Y(n_1089) );
OA22x2_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_887), .B1(n_936), .B2(n_937), .Y(n_853) );
INVx1_ASAP7_75t_L g936 ( .A(n_854), .Y(n_936) );
INVx1_ASAP7_75t_L g886 ( .A(n_855), .Y(n_886) );
AND2x2_ASAP7_75t_SL g855 ( .A(n_856), .B(n_872), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_864), .C(n_868), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_861), .Y(n_857) );
INVx2_ASAP7_75t_L g971 ( .A(n_860), .Y(n_971) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NOR3xp33_ASAP7_75t_SL g872 ( .A(n_873), .B(n_876), .C(n_881), .Y(n_872) );
INVx1_ASAP7_75t_L g937 ( .A(n_887), .Y(n_937) );
XOR2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_912), .Y(n_887) );
INVx1_ASAP7_75t_L g911 ( .A(n_890), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_901), .Y(n_890) );
NOR2xp67_ASAP7_75t_L g891 ( .A(n_892), .B(n_896), .Y(n_891) );
OAI21xp5_ASAP7_75t_SL g892 ( .A1(n_893), .A2(n_894), .B(n_895), .Y(n_892) );
OAI21xp33_ASAP7_75t_L g952 ( .A1(n_893), .A2(n_953), .B(n_954), .Y(n_952) );
OAI21xp5_ASAP7_75t_SL g1132 ( .A1(n_893), .A2(n_1133), .B(n_1134), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .C(n_900), .Y(n_896) );
NOR2x1_ASAP7_75t_L g901 ( .A(n_902), .B(n_905), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_909), .Y(n_905) );
INVx2_ASAP7_75t_L g935 ( .A(n_914), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_927), .Y(n_914) );
NOR3xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_921), .C(n_924), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g1090 ( .A(n_938), .Y(n_1090) );
XOR2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_1017), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B1(n_991), .B2(n_1016), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B1(n_974), .B2(n_975), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_944), .A2(n_1039), .B1(n_1040), .B2(n_1086), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_944), .Y(n_1039) );
INVx2_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_948), .B(n_960), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .C(n_955), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_958), .Y(n_957) );
NOR3xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_965), .C(n_970), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
NAND4xp75_ASAP7_75t_L g976 ( .A(n_977), .B(n_981), .C(n_985), .D(n_990), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
AND2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
BUFx4f_ASAP7_75t_SL g1077 ( .A(n_983), .Y(n_1077) );
INVx1_ASAP7_75t_L g1016 ( .A(n_991), .Y(n_1016) );
XOR2x2_ASAP7_75t_L g991 ( .A(n_992), .B(n_1015), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_1007), .Y(n_992) );
NOR3xp33_ASAP7_75t_L g993 ( .A(n_994), .B(n_998), .C(n_1003), .Y(n_993) );
OAI21xp33_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1000), .B(n_1001), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1014), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1038), .B1(n_1087), .B2(n_1088), .Y(n_1017) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1018), .Y(n_1087) );
INVx1_ASAP7_75t_SL g1037 ( .A(n_1020), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1030), .Y(n_1020) );
NOR2x1_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1027), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1034), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1038), .Y(n_1088) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1040), .Y(n_1086) );
OA22x2_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B1(n_1063), .B2(n_1085), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
XOR2x2_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1062), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1055), .Y(n_1043) );
NOR3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1048), .C(n_1051), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1059), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1063), .Y(n_1085) );
INVx1_ASAP7_75t_SL g1064 ( .A(n_1065), .Y(n_1064) );
NAND2xp5_ASAP7_75t_SL g1065 ( .A(n_1066), .B(n_1073), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1070), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .Y(n_1070) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1080), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1078), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1083), .Y(n_1080) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_SL g1092 ( .A1(n_1093), .A2(n_1094), .B1(n_1118), .B2(n_1119), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1095), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1107), .Y(n_1095) );
NOR3xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1100), .C(n_1104), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1111), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
XNOR2x2_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
NOR4xp75_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1125), .C(n_1128), .D(n_1132), .Y(n_1121) );
NAND2xp5_ASAP7_75t_SL g1122 ( .A(n_1123), .B(n_1124), .Y(n_1122) );
NAND2xp5_ASAP7_75t_SL g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
INVx1_ASAP7_75t_SL g1137 ( .A(n_1138), .Y(n_1137) );
NOR2x1_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1143), .Y(n_1138) );
OR2x2_ASAP7_75t_SL g1185 ( .A(n_1139), .B(n_1144), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1142), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1140), .B(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1141), .B(n_1178), .Y(n_1188) );
CKINVDCx16_ASAP7_75t_R g1178 ( .A(n_1142), .Y(n_1178) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_1144), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1146), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
OAI222xp33_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1177), .B1(n_1179), .B2(n_1182), .C1(n_1183), .C2(n_1186), .Y(n_1150) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1152), .Y(n_1176) );
AND2x2_ASAP7_75t_SL g1152 ( .A(n_1153), .B(n_1161), .Y(n_1152) );
NOR2xp33_ASAP7_75t_SL g1153 ( .A(n_1154), .B(n_1158), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1157), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
NOR3xp33_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1165), .C(n_1172), .Y(n_1161) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
CKINVDCx20_ASAP7_75t_R g1183 ( .A(n_1184), .Y(n_1183) );
CKINVDCx20_ASAP7_75t_R g1184 ( .A(n_1185), .Y(n_1184) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_1187), .Y(n_1186) );
endmodule