module fake_jpeg_28884_n_148 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_46),
.B1(n_49),
.B2(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_20),
.B1(n_15),
.B2(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_15),
.B1(n_28),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_24),
.B1(n_26),
.B2(n_22),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_22),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_30),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_42),
.B1(n_33),
.B2(n_3),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_7),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_79),
.B1(n_52),
.B2(n_51),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_42),
.C(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_14),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_8),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_44),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_52),
.B1(n_57),
.B2(n_51),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_85),
.B(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_33),
.B1(n_59),
.B2(n_1),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_104),
.B(n_67),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_68),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

AO21x2_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_75),
.B(n_77),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_90),
.A3(n_98),
.B1(n_75),
.B2(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_63),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_85),
.C(n_90),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_122),
.C(n_66),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_112),
.B(n_92),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_86),
.B(n_95),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_108),
.B(n_111),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_108),
.B1(n_106),
.B2(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_76),
.C(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_130),
.B1(n_129),
.B2(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_128),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_99),
.C(n_87),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_106),
.B1(n_94),
.B2(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_93),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_116),
.B(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_106),
.B1(n_134),
.B2(n_93),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_134),
.B(n_94),
.C(n_59),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_138),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_141),
.B(n_142),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_9),
.C(n_3),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_3),
.Y(n_148)
);


endmodule