module fake_jpeg_29079_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_15),
.B(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_0),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_48),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_55),
.B(n_46),
.C(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_56),
.Y(n_89)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_54),
.B1(n_57),
.B2(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_84),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_61),
.B1(n_54),
.B2(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_52),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_61),
.B1(n_49),
.B2(n_60),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_103),
.B1(n_88),
.B2(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_13),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_101),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_26),
.B1(n_41),
.B2(n_40),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_103),
.B1(n_19),
.B2(n_36),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_20),
.B1(n_39),
.B2(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_112),
.B(n_113),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_33),
.B(n_35),
.C(n_42),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_116),
.C(n_124),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

AOI31xp67_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_118),
.A3(n_120),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_115),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_107),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_104),
.Y(n_133)
);


endmodule