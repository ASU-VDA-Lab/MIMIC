module real_jpeg_22563_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_322, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_322;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_30),
.B1(n_59),
.B2(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_0),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_68),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_118),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_118),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_118),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_3),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_111),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_111),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_111),
.Y(n_191)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_5),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_6),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_10),
.B(n_59),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_8),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_107),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_107),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_107),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_9),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_113),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_113),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_113),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_34),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_116),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_96),
.B1(n_97),
.B2(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_42),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_36),
.B(n_206),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_12),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_13),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_81),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_81),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_14),
.A2(n_36),
.A3(n_45),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_16),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_16),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_22),
.B(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_27),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g115 ( 
.A(n_29),
.B(n_116),
.CON(n_115),
.SN(n_115)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_34),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_31),
.A2(n_34),
.B1(n_80),
.B2(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_32),
.B(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_33),
.A2(n_35),
.B1(n_115),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_35),
.B(n_116),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_50),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_47),
.B1(n_63),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_42),
.A2(n_47),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_42),
.A2(n_47),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_43),
.A2(n_48),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_48),
.B1(n_112),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_43),
.A2(n_48),
.B1(n_143),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_43),
.A2(n_48),
.B1(n_126),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_43),
.A2(n_48),
.B1(n_85),
.B2(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_44),
.B(n_46),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_45),
.A2(n_57),
.B(n_116),
.C(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_62),
.C(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_62),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_54),
.A2(n_77),
.B1(n_83),
.B2(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_61),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_58),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_58),
.B1(n_101),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_55),
.A2(n_58),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_55),
.A2(n_58),
.B1(n_170),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_55),
.A2(n_58),
.B1(n_191),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_55),
.A2(n_58),
.B1(n_106),
.B2(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_55),
.A2(n_58),
.B1(n_102),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_55),
.A2(n_58),
.B1(n_245),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_58),
.B(n_116),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_60),
.B(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_65),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_69),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_66),
.A2(n_69),
.B1(n_124),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_66),
.A2(n_69),
.B1(n_252),
.B2(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_82),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_308),
.Y(n_312)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.C(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_78),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_78),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_82),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_83),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_301),
.A3(n_313),
.B1(n_319),
.B2(n_320),
.C(n_322),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_282),
.B(n_300),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_258),
.B(n_281),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_149),
.B(n_234),
.C(n_257),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_134),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_92),
.B(n_134),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_119),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_94),
.B(n_103),
.C(n_119),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_95),
.B(n_100),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_98),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_97),
.B1(n_132),
.B2(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_96),
.A2(n_159),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_96),
.A2(n_133),
.B1(n_162),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_96),
.A2(n_97),
.B1(n_148),
.B2(n_193),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_96),
.A2(n_99),
.B1(n_133),
.B2(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_96),
.A2(n_97),
.B(n_243),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_116),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_114),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_128),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_121),
.B(n_127),
.C(n_128),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_131),
.Y(n_138)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_139),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_146),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_141),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_233),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_228),
.B(n_232),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_214),
.B(n_227),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_195),
.B(n_213),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_183),
.B(n_194),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_171),
.B(n_182),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_181),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_185),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_203),
.B1(n_211),
.B2(n_212),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_224),
.C(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_223),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_256),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_247),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_250),
.C(n_255),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_280),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_273),
.B2(n_274),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_274),
.C(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_276),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_293),
.B(n_296),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_284),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_298),
.B2(n_299),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_292),
.C(n_299),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_303),
.C(n_309),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_303),
.B1(n_304),
.B2(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_291),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_311),
.Y(n_320)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_310),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);


endmodule