module fake_ariane_1774_n_754 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_754);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_754;

wire n_295;
wire n_556;
wire n_356;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_552;
wire n_348;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_140;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_365;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_34),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_23),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_55),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_9),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_90),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_8),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_98),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_41),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_47),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_54),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_30),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_35),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_43),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_22),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_33),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_86),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_62),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_109),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_27),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

BUFx2_ASAP7_75t_SL g169 ( 
.A(n_70),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_46),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_78),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_1),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_63),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_50),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_53),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_44),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_0),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_1),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_2),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_2),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_4),
.Y(n_207)
);

BUFx8_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_159),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_4),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_5),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_5),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_6),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_6),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_182),
.B1(n_167),
.B2(n_162),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_175),
.B1(n_147),
.B2(n_190),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_192),
.B1(n_166),
.B2(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_191),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_166),
.B1(n_183),
.B2(n_184),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_228),
.B1(n_231),
.B2(n_222),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_192),
.B1(n_184),
.B2(n_183),
.Y(n_245)
);

AO22x2_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_169),
.B1(n_191),
.B2(n_10),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_181),
.B1(n_180),
.B2(n_174),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_171),
.B1(n_170),
.B2(n_164),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_158),
.B1(n_157),
.B2(n_155),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_154),
.B1(n_153),
.B2(n_152),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_139),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_150),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_254)
);

OR2x6_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_11),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_12),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_13),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_15),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_201),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_31),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_205),
.A2(n_206),
.B1(n_232),
.B2(n_220),
.Y(n_263)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_205),
.A2(n_201),
.B1(n_218),
.B2(n_214),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_205),
.B(n_16),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_205),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_32),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_224),
.A2(n_193),
.B1(n_195),
.B2(n_207),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_20),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_202),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_199),
.B(n_24),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_197),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_202),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

NOR2x1p5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_216),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_225),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_226),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_212),
.B(n_204),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_243),
.B(n_226),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_200),
.B(n_223),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_226),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_226),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_226),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_208),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_208),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_208),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_229),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_219),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_219),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_208),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_233),
.B(n_234),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_R g325 ( 
.A(n_255),
.B(n_229),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_255),
.B(n_229),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_200),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_254),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_255),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_200),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_219),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_251),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_251),
.B(n_230),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_219),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_276),
.B(n_200),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_240),
.B(n_219),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_240),
.B(n_200),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_240),
.B(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_243),
.B(n_200),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_238),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_230),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_230),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_194),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_196),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_196),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_332),
.A2(n_223),
.B(n_194),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_306),
.B(n_196),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_286),
.B(n_210),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_210),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g361 ( 
.A(n_299),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_318),
.B(n_210),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_213),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_213),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_213),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_213),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_213),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_217),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_217),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_217),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_217),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_217),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_307),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_217),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_316),
.B(n_198),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_302),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_340),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_223),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_283),
.B(n_223),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_223),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_315),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_283),
.B(n_223),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_337),
.B(n_28),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_28),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_304),
.B(n_36),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_291),
.B(n_37),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_38),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_293),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_290),
.B(n_138),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_332),
.A2(n_288),
.B(n_319),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_336),
.B(n_40),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_333),
.Y(n_405)
);

AND2x4_ASAP7_75t_SL g406 ( 
.A(n_329),
.B(n_137),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_303),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_311),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_280),
.B(n_42),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_304),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_346),
.B(n_284),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_321),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_361),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_282),
.Y(n_417)
);

AO21x2_ASAP7_75t_L g418 ( 
.A1(n_351),
.A2(n_369),
.B(n_353),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

CKINVDCx6p67_ASAP7_75t_R g421 ( 
.A(n_361),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_330),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_289),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_321),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_324),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_331),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_342),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_295),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

CKINVDCx10_ASAP7_75t_R g432 ( 
.A(n_391),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_354),
.B(n_403),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_325),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_371),
.B(n_407),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_387),
.B(n_45),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

NAND2x1_ASAP7_75t_L g439 ( 
.A(n_350),
.B(n_49),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_51),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_56),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_57),
.Y(n_442)
);

NOR2x1_ASAP7_75t_SL g443 ( 
.A(n_412),
.B(n_58),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_344),
.B(n_59),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_60),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_354),
.B(n_61),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_407),
.B(n_64),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_69),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_344),
.B(n_71),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_74),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_358),
.B(n_75),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_397),
.B(n_76),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_410),
.B(n_77),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_80),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_347),
.B(n_81),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_82),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_350),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_397),
.B(n_406),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_359),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_398),
.B(n_83),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_359),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_358),
.B(n_84),
.Y(n_467)
);

BUFx8_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_397),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_432),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_410),
.Y(n_476)
);

CKINVDCx6p67_ASAP7_75t_R g477 ( 
.A(n_432),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_400),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_363),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

BUFx6f_ASAP7_75t_SL g481 ( 
.A(n_422),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_347),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_374),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_453),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_453),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_453),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_416),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_426),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_441),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_406),
.B1(n_373),
.B2(n_370),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_436),
.B(n_393),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_419),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_417),
.Y(n_501)
);

INVx3_ASAP7_75t_SL g502 ( 
.A(n_417),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_449),
.A2(n_383),
.B1(n_404),
.B2(n_365),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_414),
.B(n_347),
.Y(n_506)
);

CKINVDCx6p67_ASAP7_75t_R g507 ( 
.A(n_437),
.Y(n_507)
);

BUFx4_ASAP7_75t_SL g508 ( 
.A(n_457),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_424),
.Y(n_509)
);

BUFx12f_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_463),
.A2(n_406),
.B1(n_373),
.B2(n_370),
.Y(n_511)
);

INVx2_ASAP7_75t_R g512 ( 
.A(n_444),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_469),
.A2(n_413),
.B1(n_456),
.B2(n_449),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_506),
.A2(n_413),
.B1(n_434),
.B2(n_442),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_468),
.B1(n_435),
.B2(n_415),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_475),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_497),
.A2(n_415),
.B1(n_458),
.B2(n_424),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_479),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_495),
.Y(n_522)
);

INVx8_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_497),
.A2(n_415),
.B1(n_458),
.B2(n_429),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_415),
.B1(n_373),
.B2(n_364),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_511),
.A2(n_370),
.B1(n_364),
.B2(n_442),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_470),
.A2(n_434),
.B1(n_383),
.B2(n_447),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_490),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_485),
.A2(n_364),
.B1(n_447),
.B2(n_408),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_485),
.A2(n_408),
.B1(n_390),
.B2(n_349),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_474),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_485),
.A2(n_390),
.B1(n_349),
.B2(n_352),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_485),
.A2(n_451),
.B1(n_395),
.B2(n_430),
.Y(n_538)
);

BUFx8_ASAP7_75t_SL g539 ( 
.A(n_500),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_477),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_484),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_496),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_485),
.A2(n_349),
.B1(n_352),
.B2(n_451),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_476),
.A2(n_352),
.B1(n_428),
.B2(n_420),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_481),
.A2(n_362),
.B1(n_365),
.B2(n_360),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_481),
.A2(n_480),
.B1(n_505),
.B2(n_478),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_503),
.A2(n_452),
.B1(n_430),
.B2(n_360),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_479),
.B(n_374),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_490),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_512),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_514),
.A2(n_473),
.B(n_504),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_543),
.A2(n_478),
.B1(n_507),
.B2(n_495),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_518),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_525),
.B(n_507),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_548),
.A2(n_495),
.B1(n_505),
.B2(n_443),
.Y(n_558)
);

AOI22x1_ASAP7_75t_SL g559 ( 
.A1(n_540),
.A2(n_500),
.B1(n_477),
.B2(n_509),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_524),
.A2(n_478),
.B1(n_512),
.B2(n_402),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_533),
.A2(n_412),
.B1(n_368),
.B2(n_378),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_520),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_539),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_529),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_526),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_529),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_552),
.Y(n_567)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_515),
.A2(n_452),
.B(n_351),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_498),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_519),
.A2(n_368),
.B1(n_378),
.B2(n_501),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_538),
.A2(n_498),
.B1(n_471),
.B2(n_502),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_539),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_528),
.A2(n_446),
.B1(n_437),
.B2(n_450),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_531),
.A2(n_510),
.B1(n_482),
.B2(n_502),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_532),
.A2(n_471),
.B1(n_366),
.B2(n_438),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_537),
.A2(n_366),
.B1(n_362),
.B2(n_437),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_542),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_516),
.A2(n_450),
.B1(n_446),
.B2(n_510),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_535),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_552),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_545),
.A2(n_450),
.B1(n_446),
.B2(n_357),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_520),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_527),
.A2(n_450),
.B1(n_446),
.B2(n_357),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_552),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_549),
.A2(n_398),
.B1(n_379),
.B2(n_367),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_551),
.A2(n_508),
.B(n_471),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_523),
.A2(n_482),
.B1(n_467),
.B2(n_454),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_547),
.A2(n_367),
.B1(n_379),
.B2(n_363),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_552),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_523),
.A2(n_353),
.B1(n_440),
.B2(n_369),
.Y(n_591)
);

OAI21xp33_ASAP7_75t_L g592 ( 
.A1(n_544),
.A2(n_348),
.B(n_376),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_536),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_540),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_L g595 ( 
.A1(n_517),
.A2(n_348),
.B(n_376),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_552),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_517),
.A2(n_461),
.B1(n_513),
.B2(n_494),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_536),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_558),
.B(n_522),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_557),
.A2(n_523),
.B1(n_522),
.B2(n_541),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_546),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_554),
.A2(n_520),
.B1(n_541),
.B2(n_530),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_557),
.A2(n_523),
.B1(n_522),
.B2(n_541),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_557),
.A2(n_379),
.B1(n_367),
.B2(n_418),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_584),
.A2(n_573),
.B1(n_579),
.B2(n_570),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_555),
.A2(n_559),
.B1(n_571),
.B2(n_553),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_556),
.A2(n_418),
.B1(n_401),
.B2(n_472),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_553),
.B(n_535),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_559),
.A2(n_541),
.B1(n_520),
.B2(n_530),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_582),
.A2(n_401),
.B1(n_472),
.B2(n_546),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_587),
.B(n_534),
.C(n_492),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_565),
.A2(n_530),
.B1(n_534),
.B2(n_535),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_564),
.Y(n_614)
);

AOI222xp33_ASAP7_75t_L g615 ( 
.A1(n_577),
.A2(n_448),
.B1(n_377),
.B2(n_374),
.C1(n_382),
.C2(n_465),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_401),
.B1(n_382),
.B2(n_465),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_569),
.B(n_535),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_561),
.A2(n_530),
.B1(n_513),
.B2(n_494),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_593),
.B(n_536),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_560),
.A2(n_513),
.B1(n_494),
.B2(n_550),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_576),
.A2(n_382),
.B1(n_460),
.B2(n_550),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_569),
.B(n_491),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_491),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_589),
.A2(n_401),
.B1(n_382),
.B2(n_460),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_592),
.A2(n_401),
.B1(n_382),
.B2(n_377),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_568),
.B1(n_575),
.B2(n_566),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_575),
.A2(n_401),
.B1(n_382),
.B2(n_377),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_574),
.A2(n_492),
.B1(n_489),
.B2(n_487),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_591),
.A2(n_550),
.B1(n_439),
.B2(n_426),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_401),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_566),
.A2(n_382),
.B1(n_381),
.B2(n_388),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_595),
.A2(n_597),
.B1(n_594),
.B2(n_382),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_594),
.A2(n_462),
.B1(n_375),
.B2(n_372),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_578),
.A2(n_381),
.B1(n_385),
.B2(n_388),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_562),
.B(n_462),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_595),
.C(n_598),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_633),
.B(n_598),
.C(n_596),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_609),
.B(n_590),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_606),
.A2(n_563),
.B1(n_572),
.B2(n_562),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_607),
.A2(n_567),
.B(n_563),
.Y(n_640)
);

OAI221xp5_ASAP7_75t_SL g641 ( 
.A1(n_632),
.A2(n_596),
.B1(n_590),
.B2(n_585),
.C(n_581),
.Y(n_641)
);

OA21x2_ASAP7_75t_L g642 ( 
.A1(n_608),
.A2(n_626),
.B(n_605),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_615),
.A2(n_578),
.B1(n_380),
.B2(n_375),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_601),
.B(n_562),
.Y(n_644)
);

AOI221xp5_ASAP7_75t_L g645 ( 
.A1(n_604),
.A2(n_372),
.B1(n_380),
.B2(n_581),
.C(n_585),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_610),
.A2(n_567),
.B(n_572),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_583),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_609),
.B(n_567),
.Y(n_648)
);

OAI21xp33_ASAP7_75t_L g649 ( 
.A1(n_613),
.A2(n_345),
.B(n_381),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_602),
.B(n_583),
.C(n_462),
.Y(n_650)
);

NAND4xp25_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_583),
.C(n_345),
.D(n_389),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_630),
.B(n_345),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_629),
.A2(n_488),
.B1(n_487),
.B2(n_486),
.Y(n_653)
);

AOI211xp5_ASAP7_75t_SL g654 ( 
.A1(n_628),
.A2(n_345),
.B(n_394),
.C(n_389),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_630),
.B(n_619),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_617),
.B(n_488),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_623),
.B(n_388),
.C(n_385),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_486),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_604),
.B(n_385),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_614),
.B(n_85),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_614),
.B(n_384),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_600),
.A2(n_394),
.B1(n_356),
.B2(n_355),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_599),
.B(n_384),
.C(n_356),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_603),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_659),
.Y(n_665)
);

AO21x2_ASAP7_75t_L g666 ( 
.A1(n_661),
.A2(n_599),
.B(n_635),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

OAI211xp5_ASAP7_75t_SL g668 ( 
.A1(n_640),
.A2(n_621),
.B(n_618),
.C(n_616),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_611),
.C(n_625),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_655),
.B(n_620),
.Y(n_670)
);

NOR2x1_ASAP7_75t_L g671 ( 
.A(n_636),
.B(n_356),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_634),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_638),
.B(n_627),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_642),
.A2(n_624),
.B1(n_631),
.B2(n_356),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_644),
.B(n_384),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_642),
.A2(n_355),
.B1(n_350),
.B2(n_91),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_648),
.B(n_88),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_642),
.A2(n_355),
.B1(n_350),
.B2(n_93),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_650),
.B(n_89),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_664),
.B(n_639),
.Y(n_680)
);

BUFx2_ASAP7_75t_SL g681 ( 
.A(n_664),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_665),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_670),
.B(n_648),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_665),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_670),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_667),
.Y(n_686)
);

XNOR2xp5_ASAP7_75t_L g687 ( 
.A(n_673),
.B(n_647),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_666),
.Y(n_689)
);

CKINVDCx14_ASAP7_75t_R g690 ( 
.A(n_677),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_682),
.Y(n_691)
);

XNOR2x2_ASAP7_75t_L g692 ( 
.A(n_680),
.B(n_669),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_685),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_681),
.Y(n_694)
);

XNOR2x2_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_683),
.Y(n_695)
);

XNOR2x2_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_671),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_SL g697 ( 
.A1(n_694),
.A2(n_690),
.B1(n_685),
.B2(n_689),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_694),
.B(n_690),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_691),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_693),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_699),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_698),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_699),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_696),
.Y(n_704)
);

AOI22x1_ASAP7_75t_L g705 ( 
.A1(n_704),
.A2(n_697),
.B1(n_693),
.B2(n_700),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_701),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_702),
.A2(n_692),
.B1(n_685),
.B2(n_668),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_701),
.A2(n_703),
.B1(n_685),
.B2(n_666),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_706),
.Y(n_709)
);

OAI211xp5_ASAP7_75t_L g710 ( 
.A1(n_705),
.A2(n_646),
.B(n_678),
.C(n_676),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_708),
.A2(n_654),
.B1(n_651),
.B2(n_663),
.Y(n_712)
);

AO22x2_ASAP7_75t_L g713 ( 
.A1(n_709),
.A2(n_711),
.B1(n_710),
.B2(n_712),
.Y(n_713)
);

NOR4xp25_ASAP7_75t_L g714 ( 
.A(n_712),
.B(n_688),
.C(n_686),
.D(n_684),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_711),
.A2(n_666),
.B1(n_672),
.B2(n_679),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_711),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_711),
.A2(n_674),
.B1(n_662),
.B2(n_649),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_711),
.A2(n_641),
.B1(n_643),
.B2(n_645),
.C(n_675),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_713),
.Y(n_719)
);

INVxp33_ASAP7_75t_SL g720 ( 
.A(n_714),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_715),
.A2(n_643),
.B1(n_658),
.B2(n_653),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_718),
.A2(n_652),
.B1(n_656),
.B2(n_660),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_717),
.B(n_652),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_713),
.A2(n_660),
.B1(n_657),
.B2(n_96),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_720),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_726)
);

AND4x1_ASAP7_75t_L g727 ( 
.A(n_722),
.B(n_99),
.C(n_100),
.D(n_101),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_719),
.Y(n_728)
);

AND4x1_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_103),
.C(n_104),
.D(n_106),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_724),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_723),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_721),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_722),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_722),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_SL g735 ( 
.A1(n_728),
.A2(n_726),
.B1(n_733),
.B2(n_734),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_731),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_732),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_727),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_729),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_728),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_742),
.B1(n_741),
.B2(n_739),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_736),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_735),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_737),
.B1(n_744),
.B2(n_746),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_749),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_748),
.B(n_124),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_751),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_752),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.C(n_127),
.Y(n_753)
);

AOI211xp5_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_128),
.B(n_129),
.C(n_130),
.Y(n_754)
);


endmodule