module fake_jpeg_25322_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_0),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_3),
.B(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_17),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_11),
.B(n_20),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_27),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_10),
.B1(n_2),
.B2(n_5),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_3),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.C(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_26),
.C(n_34),
.Y(n_43)
);

XOR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_2),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_7),
.B(n_35),
.C(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B(n_38),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_47),
.C(n_42),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_52),
.Y(n_55)
);


endmodule