module fake_jpeg_2287_n_195 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_1),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_1),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_62),
.B1(n_47),
.B2(n_48),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_62),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_90),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_45),
.B(n_49),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_94),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_55),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_48),
.C(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_51),
.B1(n_44),
.B2(n_43),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_46),
.B1(n_56),
.B2(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_118),
.B1(n_114),
.B2(n_61),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_120),
.Y(n_141)
);

OAI22x1_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_59),
.B1(n_61),
.B2(n_28),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_4),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_6),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_5),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_126),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_104),
.B1(n_100),
.B2(n_96),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_110),
.C(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_145),
.C(n_7),
.Y(n_149)
);

NAND2x1_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_91),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_7),
.B(n_10),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_31),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_59),
.B(n_61),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_25),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_59),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_12),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_26),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_154),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_125),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_161),
.C(n_37),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_35),
.C(n_41),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_158),
.C(n_20),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_29),
.C(n_40),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_126),
.B1(n_18),
.B2(n_19),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_21),
.B(n_39),
.C(n_14),
.D(n_15),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_164),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_13),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_173),
.C(n_153),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_13),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_158),
.C(n_149),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_157),
.B(n_156),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_179),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_185),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_169),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_170),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_189),
.A2(n_157),
.B(n_177),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_192),
.B(n_188),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_161),
.Y(n_195)
);


endmodule