module fake_netlist_6_2513_n_171 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_29, n_25, n_171);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_171;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

INVxp33_ASAP7_75t_SL g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_39),
.B1(n_48),
.B2(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_31),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

OR2x6_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_44),
.Y(n_88)
);

NAND2x1p5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_50),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_53),
.B1(n_51),
.B2(n_37),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_68),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_73),
.B1(n_66),
.B2(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_73),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_72),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_47),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_103),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_90),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_90),
.B1(n_57),
.B2(n_66),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_82),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_88),
.B(n_78),
.Y(n_111)
);

AOI221x1_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_85),
.B1(n_87),
.B2(n_51),
.C(n_72),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_99),
.B1(n_98),
.B2(n_35),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_104),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_97),
.B(n_95),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_109),
.B1(n_108),
.B2(n_98),
.C(n_110),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_112),
.B(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_113),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_108),
.B(n_109),
.C(n_34),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_100),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_122),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_122),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

AOI222xp33_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_54),
.B1(n_117),
.B2(n_64),
.C1(n_100),
.C2(n_92),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_89),
.C(n_117),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_119),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_86),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_134),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_138),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_148),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_153),
.B(n_151),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_154),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_135),
.C(n_155),
.Y(n_161)
);

OR2x6_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_126),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_6),
.B(n_10),
.C(n_126),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_15),
.C(n_16),
.Y(n_164)
);

NAND5xp2_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_162),
.C(n_22),
.D(n_25),
.E(n_29),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_102),
.C(n_104),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_86),
.B1(n_71),
.B2(n_102),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_64),
.B1(n_92),
.B2(n_71),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_167),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);


endmodule