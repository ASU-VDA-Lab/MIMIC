module fake_jpeg_25372_n_229 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_SL g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_15),
.B1(n_19),
.B2(n_14),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_40),
.B(n_16),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_15),
.B1(n_19),
.B2(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_31),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_60),
.B1(n_13),
.B2(n_55),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_60),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_57),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_59),
.B1(n_42),
.B2(n_13),
.Y(n_61)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_18),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_39),
.B1(n_33),
.B2(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_72),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_18),
.C(n_17),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_18),
.A3(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_39),
.B1(n_33),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_36),
.B1(n_35),
.B2(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_89),
.Y(n_96)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_53),
.B1(n_39),
.B2(n_33),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_77),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_64),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_94),
.B1(n_61),
.B2(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_88),
.B(n_79),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_108),
.B(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_91),
.B1(n_78),
.B2(n_87),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_108),
.B1(n_110),
.B2(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_95),
.B(n_77),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_23),
.B(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_102),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_69),
.C(n_81),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_128),
.C(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_107),
.C(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_93),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_96),
.C(n_102),
.D(n_108),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_149),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_140),
.B1(n_134),
.B2(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_21),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_66),
.C(n_71),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.C(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_71),
.C(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_104),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_20),
.C(n_21),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_104),
.B(n_1),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_117),
.B1(n_116),
.B2(n_126),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_148),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_128),
.C(n_123),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_163),
.C(n_150),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_164),
.B1(n_168),
.B2(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_123),
.C(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_114),
.B1(n_127),
.B2(n_121),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_113),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_113),
.B1(n_131),
.B2(n_35),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_136),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_182),
.C(n_17),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_143),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_18),
.B1(n_7),
.B2(n_8),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_161),
.C(n_158),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_113),
.B(n_149),
.C(n_2),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_159),
.B(n_1),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_0),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_173),
.C(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_189),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_5),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_183),
.B(n_5),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_201),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_183),
.B(n_8),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_202),
.B(n_194),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_198),
.A2(n_199),
.B(n_205),
.C(n_187),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_183),
.B(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_18),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_4),
.B(n_10),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_0),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_207),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_191),
.B(n_9),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_185),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_188),
.C(n_212),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_220),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_9),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_10),
.B(n_11),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.C(n_2),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_1),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_218),
.B(n_215),
.C(n_3),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);


endmodule