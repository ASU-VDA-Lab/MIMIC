module real_aes_7149_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_0), .A2(n_176), .B(n_177), .C(n_181), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_1), .B(n_170), .Y(n_183) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_3), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_4), .A2(n_164), .B(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_144), .B(n_161), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_6), .A2(n_164), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_7), .B(n_170), .Y(n_482) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_8), .A2(n_136), .B(n_258), .Y(n_257) );
AND2x6_ASAP7_75t_L g161 ( .A(n_9), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_10), .A2(n_144), .B(n_161), .C(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g573 ( .A(n_11), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_39), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_13), .B(n_180), .Y(n_522) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_15), .B(n_155), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_16), .A2(n_156), .B(n_531), .C(n_533), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_17), .B(n_170), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_18), .B(n_198), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_19), .A2(n_144), .B(n_190), .C(n_197), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_20), .A2(n_179), .B(n_232), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_21), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_22), .B(n_180), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_23), .B(n_180), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_24), .Y(n_500) );
INVx1_ASAP7_75t_L g470 ( .A(n_25), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_26), .A2(n_144), .B(n_197), .C(n_261), .Y(n_260) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_27), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_28), .Y(n_518) );
INVx1_ASAP7_75t_L g494 ( .A(n_29), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_30), .A2(n_164), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g146 ( .A(n_31), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_32), .A2(n_159), .B(n_213), .C(n_214), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_33), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_34), .A2(n_179), .B(n_479), .C(n_481), .Y(n_478) );
INVxp67_ASAP7_75t_L g495 ( .A(n_35), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_36), .B(n_263), .Y(n_262) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_37), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_38), .A2(n_144), .B(n_197), .C(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_40), .A2(n_181), .B(n_571), .C(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_41), .B(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_42), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_43), .B(n_155), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_44), .B(n_164), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_45), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_46), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_47), .A2(n_159), .B(n_213), .C(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g178 ( .A(n_48), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_49), .A2(n_125), .B1(n_439), .B2(n_440), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_49), .Y(n_439) );
INVx1_ASAP7_75t_L g242 ( .A(n_50), .Y(n_242) );
INVx1_ASAP7_75t_L g538 ( .A(n_51), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_52), .B(n_164), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_53), .A2(n_71), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_53), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_54), .Y(n_202) );
AOI222xp33_ASAP7_75t_SL g445 ( .A1(n_55), .A2(n_109), .B1(n_446), .B2(n_452), .C1(n_721), .C2(n_722), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g569 ( .A(n_56), .Y(n_569) );
INVx1_ASAP7_75t_L g162 ( .A(n_57), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_58), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_59), .B(n_170), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_60), .A2(n_151), .B(n_196), .C(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_61), .A2(n_70), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_61), .Y(n_450) );
INVx1_ASAP7_75t_L g140 ( .A(n_62), .Y(n_140) );
INVx1_ASAP7_75t_SL g480 ( .A(n_63), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_65), .B(n_155), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_66), .B(n_170), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_67), .B(n_156), .Y(n_229) );
INVx1_ASAP7_75t_L g503 ( .A(n_68), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_69), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_70), .Y(n_451) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_72), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_73), .A2(n_144), .B(n_149), .C(n_159), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_74), .Y(n_251) );
INVx1_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_76), .A2(n_164), .B(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_77), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_78), .A2(n_164), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_79), .A2(n_188), .B(n_490), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_80), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_81), .A2(n_447), .B1(n_448), .B2(n_449), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_81), .Y(n_447) );
INVx1_ASAP7_75t_L g529 ( .A(n_82), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_83), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_84), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_85), .A2(n_164), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g532 ( .A(n_86), .Y(n_532) );
INVx2_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
INVx1_ASAP7_75t_L g521 ( .A(n_88), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_89), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_90), .B(n_180), .Y(n_230) );
INVx2_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
OR2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_111), .Y(n_123) );
OR2x2_ASAP7_75t_L g456 ( .A(n_91), .B(n_112), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_92), .A2(n_144), .B(n_159), .C(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_93), .A2(n_104), .B1(n_115), .B2(n_726), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_94), .B(n_164), .Y(n_211) );
INVx1_ASAP7_75t_L g215 ( .A(n_95), .Y(n_215) );
INVxp67_ASAP7_75t_L g254 ( .A(n_96), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_97), .B(n_136), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g150 ( .A(n_99), .Y(n_150) );
INVx1_ASAP7_75t_L g225 ( .A(n_100), .Y(n_225) );
INVx2_ASAP7_75t_L g541 ( .A(n_101), .Y(n_541) );
AND2x2_ASAP7_75t_L g244 ( .A(n_102), .B(n_200), .Y(n_244) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g727 ( .A(n_105), .Y(n_727) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g720 ( .A(n_110), .B(n_112), .Y(n_720) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_444), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_117), .B(n_441), .C(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_124), .B(n_441), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_123), .Y(n_443) );
INVx1_ASAP7_75t_L g440 ( .A(n_125), .Y(n_440) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
INVx1_ASAP7_75t_L g453 ( .A(n_129), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_129), .A2(n_458), .B1(n_723), .B2(n_724), .Y(n_722) );
OR3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_347), .C(n_396), .Y(n_129) );
NAND5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_281), .C(n_310), .D(n_318), .E(n_333), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_204), .B(n_220), .C(n_265), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_184), .Y(n_132) );
AND2x2_ASAP7_75t_L g276 ( .A(n_133), .B(n_273), .Y(n_276) );
AND2x2_ASAP7_75t_L g309 ( .A(n_133), .B(n_185), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_133), .B(n_208), .Y(n_402) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
INVx2_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
BUFx2_ASAP7_75t_L g376 ( .A(n_134), .Y(n_376) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_167), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_135), .B(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_135), .B(n_219), .Y(n_218) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_135), .A2(n_224), .B(n_234), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_135), .B(n_473), .Y(n_472) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_135), .A2(n_499), .B(n_506), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_135), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_136), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_136), .A2(n_259), .B(n_260), .Y(n_258) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g236 ( .A(n_137), .Y(n_236) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_138), .B(n_139), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_163), .Y(n_142) );
INVx5_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
BUFx3_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx1_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_148), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_148), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx1_ASAP7_75t_L g263 ( .A(n_148), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .C(n_157), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_152), .A2(n_155), .B1(n_494), .B2(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_152), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_152), .B(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_155), .B(n_254), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_155), .A2(n_195), .B(n_470), .C(n_471), .Y(n_469) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_156), .B(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g481 ( .A(n_158), .Y(n_481) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_160), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_160), .A2(n_174), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_160), .A2(n_174), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_160), .A2(n_174), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_160), .A2(n_174), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_160), .A2(n_174), .B(n_538), .C(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_160), .A2(n_174), .B(n_569), .C(n_570), .Y(n_568) );
INVx4_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g164 ( .A(n_161), .B(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_161), .B(n_165), .Y(n_226) );
BUFx2_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
INVx1_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
AND2x2_ASAP7_75t_L g184 ( .A(n_169), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
AND2x2_ASAP7_75t_L g360 ( .A(n_169), .B(n_273), .Y(n_360) );
AND2x2_ASAP7_75t_L g415 ( .A(n_169), .B(n_207), .Y(n_415) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_169) );
INVx2_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_179), .B(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g571 ( .A(n_180), .Y(n_571) );
INVx2_ASAP7_75t_L g505 ( .A(n_181), .Y(n_505) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_182), .Y(n_217) );
INVx1_ASAP7_75t_L g533 ( .A(n_182), .Y(n_533) );
INVx1_ASAP7_75t_L g332 ( .A(n_184), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_184), .B(n_208), .Y(n_379) );
INVx5_ASAP7_75t_L g273 ( .A(n_185), .Y(n_273) );
AND2x4_ASAP7_75t_L g294 ( .A(n_185), .B(n_274), .Y(n_294) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_185), .Y(n_316) );
AND2x2_ASAP7_75t_L g391 ( .A(n_185), .B(n_376), .Y(n_391) );
AND2x2_ASAP7_75t_L g394 ( .A(n_185), .B(n_209), .Y(n_394) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_201), .Y(n_185) );
AOI21xp5_ASAP7_75t_SL g186 ( .A1(n_187), .A2(n_189), .B(n_198), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_195), .Y(n_190) );
INVx2_ASAP7_75t_L g194 ( .A(n_192), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_194), .A2(n_215), .B(n_216), .C(n_217), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_194), .A2(n_217), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_194), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_194), .A2(n_505), .B(n_521), .C(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_196), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_199), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g203 ( .A(n_200), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_200), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_200), .A2(n_239), .B(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_200), .A2(n_226), .B(n_467), .C(n_468), .Y(n_466) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_200), .A2(n_567), .B(n_574), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_203), .A2(n_517), .B(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_204), .B(n_274), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_204), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
AND2x2_ASAP7_75t_L g299 ( .A(n_206), .B(n_274), .Y(n_299) );
AND2x2_ASAP7_75t_L g317 ( .A(n_206), .B(n_209), .Y(n_317) );
INVx1_ASAP7_75t_L g337 ( .A(n_206), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_206), .B(n_273), .Y(n_382) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_206), .Y(n_424) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_208), .B(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_208), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_208), .A2(n_269), .B(n_330), .C(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g336 ( .A(n_208), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_208), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_208), .B(n_273), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_208), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g364 ( .A(n_208), .B(n_274), .Y(n_364) );
AND2x2_ASAP7_75t_L g414 ( .A(n_208), .B(n_415), .Y(n_414) );
INVx5_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx2_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
AND2x2_ASAP7_75t_L g319 ( .A(n_209), .B(n_272), .Y(n_319) );
AND2x2_ASAP7_75t_L g331 ( .A(n_209), .B(n_306), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_209), .B(n_360), .Y(n_378) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_245), .Y(n_220) );
INVx1_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_237), .Y(n_221) );
OR2x2_ASAP7_75t_L g269 ( .A(n_222), .B(n_237), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_222), .B(n_276), .C(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_222), .B(n_247), .Y(n_286) );
OR2x2_ASAP7_75t_L g301 ( .A(n_222), .B(n_289), .Y(n_301) );
AND2x2_ASAP7_75t_L g307 ( .A(n_222), .B(n_256), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_222), .B(n_438), .Y(n_437) );
INVx5_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_223), .B(n_247), .Y(n_304) );
AND2x2_ASAP7_75t_L g343 ( .A(n_223), .B(n_257), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_223), .B(n_256), .Y(n_371) );
OR2x2_ASAP7_75t_L g374 ( .A(n_223), .B(n_256), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_226), .A2(n_500), .B(n_501), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_226), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_262), .B(n_264), .Y(n_261) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g488 ( .A(n_236), .Y(n_488) );
INVx5_ASAP7_75t_SL g289 ( .A(n_237), .Y(n_289) );
OR2x2_ASAP7_75t_L g295 ( .A(n_237), .B(n_246), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_237), .B(n_312), .Y(n_311) );
AOI321xp33_ASAP7_75t_L g318 ( .A1(n_237), .A2(n_319), .A3(n_320), .B1(n_321), .B2(n_327), .C(n_329), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_237), .B(n_245), .Y(n_328) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_237), .Y(n_341) );
OR2x2_ASAP7_75t_L g388 ( .A(n_237), .B(n_286), .Y(n_388) );
AND2x2_ASAP7_75t_L g410 ( .A(n_237), .B(n_307), .Y(n_410) );
AND2x2_ASAP7_75t_L g429 ( .A(n_237), .B(n_247), .Y(n_429) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_256), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_247), .B(n_256), .Y(n_270) );
AND2x2_ASAP7_75t_L g279 ( .A(n_247), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g306 ( .A(n_247), .Y(n_306) );
AND2x2_ASAP7_75t_L g312 ( .A(n_247), .B(n_307), .Y(n_312) );
INVxp67_ASAP7_75t_L g342 ( .A(n_247), .Y(n_342) );
OR2x2_ASAP7_75t_L g384 ( .A(n_247), .B(n_289), .Y(n_384) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_255), .Y(n_247) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_248), .A2(n_475), .B(n_482), .Y(n_474) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_248), .A2(n_527), .B(n_534), .Y(n_526) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_248), .A2(n_536), .B(n_542), .Y(n_535) );
OR2x2_ASAP7_75t_L g266 ( .A(n_256), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_SL g280 ( .A(n_256), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_256), .B(n_269), .Y(n_313) );
AND2x2_ASAP7_75t_L g362 ( .A(n_256), .B(n_306), .Y(n_362) );
AND2x2_ASAP7_75t_L g400 ( .A(n_256), .B(n_289), .Y(n_400) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_257), .B(n_289), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B(n_271), .C(n_275), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_266), .A2(n_268), .B1(n_393), .B2(n_395), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_268), .A2(n_291), .B1(n_346), .B2(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_SL g420 ( .A(n_269), .Y(n_420) );
INVx1_ASAP7_75t_SL g320 ( .A(n_270), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_272), .B(n_292), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g333 ( .A1(n_272), .A2(n_313), .B1(n_320), .B2(n_334), .C1(n_338), .C2(n_344), .Y(n_333) );
AND2x2_ASAP7_75t_L g423 ( .A(n_272), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_273), .B(n_293), .Y(n_368) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_273), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_273), .B(n_317), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_273), .B(n_424), .Y(n_434) );
INVx1_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_274), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g416 ( .A1(n_276), .A2(n_417), .B(n_418), .C(n_421), .Y(n_416) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_278), .B(n_340), .C(n_343), .Y(n_339) );
OR2x2_ASAP7_75t_L g367 ( .A(n_278), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_278), .B(n_294), .Y(n_395) );
OR2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
AOI211xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B(n_290), .C(n_302), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_283), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g389 ( .A(n_284), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_285), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g303 ( .A(n_288), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_289), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g357 ( .A(n_289), .B(n_307), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_289), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_289), .B(n_306), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B1(n_296), .B2(n_300), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_292), .B(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_294), .B(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g358 ( .A1(n_295), .A2(n_359), .B1(n_361), .B2(n_363), .C(n_365), .Y(n_358) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g413 ( .A(n_298), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g426 ( .A(n_298), .B(n_415), .Y(n_426) );
INVx1_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g417 ( .A(n_300), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_301), .A2(n_384), .B(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_308), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI21xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_313), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_L g350 ( .A(n_311), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_312), .A2(n_398), .B1(n_401), .B2(n_403), .C(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_320), .A2(n_410), .B1(n_411), .B2(n_413), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g386 ( .A(n_322), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g390 ( .A(n_326), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_336), .B(n_360), .Y(n_412) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_342), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g435 ( .A(n_343), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI211xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_350), .B(n_351), .C(n_385), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_358), .C(n_377), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g438 ( .A(n_362), .Y(n_438) );
AND2x2_ASAP7_75t_L g375 ( .A(n_364), .B(n_376), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B1(n_373), .B2(n_375), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g383 ( .A(n_371), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g436 ( .A(n_372), .Y(n_436) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI31xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .A3(n_380), .B(n_383), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_389), .C(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
NAND5xp2_ASAP7_75t_L g396 ( .A(n_397), .B(n_409), .C(n_416), .D(n_430), .E(n_433), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_434), .B1(n_435), .B2(n_437), .Y(n_433) );
INVx1_ASAP7_75t_SL g432 ( .A(n_410), .Y(n_432) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_427), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g721 ( .A(n_446), .Y(n_721) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B1(n_457), .B2(n_720), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g723 ( .A(n_455), .Y(n_723) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR3x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_631), .C(n_678), .Y(n_458) );
NAND3xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_577), .C(n_602), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_515), .B1(n_543), .B2(n_546), .C(n_554), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_483), .B(n_508), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_463), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_463), .B(n_559), .Y(n_675) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AND2x2_ASAP7_75t_L g545 ( .A(n_464), .B(n_514), .Y(n_545) );
AND2x2_ASAP7_75t_L g595 ( .A(n_464), .B(n_513), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_464), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_464), .B(n_588), .Y(n_621) );
OR2x2_ASAP7_75t_L g629 ( .A(n_464), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g701 ( .A(n_464), .B(n_497), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_464), .B(n_650), .Y(n_715) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g560 ( .A(n_465), .B(n_474), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_465), .B(n_497), .Y(n_561) );
AND2x4_ASAP7_75t_L g583 ( .A(n_465), .B(n_514), .Y(n_583) );
AND2x2_ASAP7_75t_L g613 ( .A(n_465), .B(n_485), .Y(n_613) );
AND2x2_ASAP7_75t_L g622 ( .A(n_465), .B(n_612), .Y(n_622) );
AND2x2_ASAP7_75t_L g638 ( .A(n_465), .B(n_498), .Y(n_638) );
OR2x2_ASAP7_75t_L g647 ( .A(n_465), .B(n_630), .Y(n_647) );
AND2x2_ASAP7_75t_L g653 ( .A(n_465), .B(n_588), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_465), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g667 ( .A(n_465), .B(n_510), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_465), .B(n_556), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_465), .B(n_617), .Y(n_706) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
INVx2_ASAP7_75t_L g514 ( .A(n_474), .Y(n_514) );
AND2x2_ASAP7_75t_L g612 ( .A(n_474), .B(n_497), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_498), .Y(n_617) );
INVx1_ASAP7_75t_L g673 ( .A(n_474), .Y(n_673) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g582 ( .A(n_484), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_497), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_485), .B(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
OR2x2_ASAP7_75t_L g630 ( .A(n_485), .B(n_497), .Y(n_630) );
OR2x2_ASAP7_75t_L g691 ( .A(n_485), .B(n_598), .Y(n_691) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B(n_496), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_487), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g511 ( .A(n_489), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_496), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_497), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g650 ( .A(n_497), .B(n_510), .Y(n_650) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g589 ( .A(n_498), .Y(n_589) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_509), .A2(n_695), .B1(n_699), .B2(n_702), .C(n_703), .Y(n_694) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx1_ASAP7_75t_SL g557 ( .A(n_510), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_510), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_545), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_513), .B(n_559), .Y(n_681) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g592 ( .A(n_515), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_515), .B(n_598), .Y(n_628) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
AND2x2_ASAP7_75t_L g553 ( .A(n_516), .B(n_526), .Y(n_553) );
INVx4_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
BUFx3_ASAP7_75t_L g608 ( .A(n_516), .Y(n_608) );
AND3x2_ASAP7_75t_L g623 ( .A(n_516), .B(n_624), .C(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g705 ( .A(n_525), .B(n_619), .Y(n_705) );
AND2x2_ASAP7_75t_L g713 ( .A(n_525), .B(n_598), .Y(n_713) );
INVx1_ASAP7_75t_SL g718 ( .A(n_525), .Y(n_718) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
INVx1_ASAP7_75t_SL g576 ( .A(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_565), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_526), .B(n_549), .Y(n_601) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_526), .Y(n_641) );
OR2x2_ASAP7_75t_L g646 ( .A(n_526), .B(n_565), .Y(n_646) );
INVx2_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
AND2x2_ASAP7_75t_L g586 ( .A(n_535), .B(n_566), .Y(n_586) );
OR2x2_ASAP7_75t_L g606 ( .A(n_535), .B(n_566), .Y(n_606) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_535), .Y(n_626) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_544), .A2(n_585), .B(n_677), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_546), .A2(n_556), .A3(n_583), .B1(n_713), .B2(n_714), .C1(n_716), .C2(n_719), .Y(n_712) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_548), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_549), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g575 ( .A(n_550), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_565), .Y(n_643) );
AND2x2_ASAP7_75t_L g710 ( .A(n_551), .B(n_566), .Y(n_710) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g651 ( .A(n_553), .B(n_605), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .A3(n_561), .B(n_562), .Y(n_554) );
AND2x2_ASAP7_75t_L g610 ( .A(n_556), .B(n_588), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_556), .B(n_580), .Y(n_692) );
AND2x2_ASAP7_75t_L g711 ( .A(n_556), .B(n_616), .Y(n_711) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_559), .B(n_588), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_559), .B(n_617), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_559), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_559), .B(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_560), .B(n_617), .Y(n_649) );
INVx1_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_575), .Y(n_563) );
INVxp67_ASAP7_75t_L g645 ( .A(n_564), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_565), .B(n_576), .Y(n_581) );
INVx1_ASAP7_75t_L g687 ( .A(n_565), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_565), .B(n_664), .Y(n_698) );
BUFx3_ASAP7_75t_L g598 ( .A(n_566), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_576), .Y(n_624) );
INVx2_ASAP7_75t_L g664 ( .A(n_566), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_575), .B(n_697), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_582), .B(n_584), .C(n_593), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_579), .A2(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_580), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_580), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g660 ( .A(n_581), .B(n_606), .Y(n_660) );
INVx3_ASAP7_75t_L g591 ( .A(n_583), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B1(n_590), .B2(n_592), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_586), .A2(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g635 ( .A(n_586), .B(n_599), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_586), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g590 ( .A(n_589), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g659 ( .A(n_589), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_590), .A2(n_604), .B(n_609), .Y(n_603) );
OAI22xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B1(n_600), .B2(n_601), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_595), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g619 ( .A(n_598), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_641), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_614), .C(n_627), .Y(n_602) );
OAI22xp5_ASAP7_75t_SL g669 ( .A1(n_604), .A2(n_670), .B1(n_674), .B2(n_675), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g674 ( .A(n_606), .B(n_607), .Y(n_674) );
AND2x2_ASAP7_75t_L g682 ( .A(n_607), .B(n_663), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_SL g690 ( .A1(n_608), .A2(n_691), .B(n_692), .C(n_693), .Y(n_690) );
OR2x2_ASAP7_75t_L g717 ( .A(n_608), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B(n_620), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_616), .A2(n_653), .B(n_654), .C(n_657), .Y(n_652) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_622), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g685 ( .A(n_624), .B(n_643), .Y(n_685) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g663 ( .A(n_626), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_628), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_652), .C(n_665), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_636), .C(n_644), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g702 ( .A(n_639), .Y(n_702) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_641), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_647), .C(n_648), .Y(n_644) );
INVx2_ASAP7_75t_SL g656 ( .A(n_646), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_647), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_657) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_669), .C(n_676), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp33_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g719 ( .A(n_673), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_694), .C(n_707), .D(n_712), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B(n_683), .C(n_690), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_688), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g703 ( .A1(n_684), .A2(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_691), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g725 ( .A(n_720), .Y(n_725) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
endmodule