module fake_jpeg_6567_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_31),
.Y(n_57)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_52),
.B1(n_24),
.B2(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_54),
.Y(n_75)
);

AO22x2_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_32),
.B1(n_19),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_28),
.B1(n_17),
.B2(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_39),
.B1(n_46),
.B2(n_56),
.Y(n_70)
);

AO21x2_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_0),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_76),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_39),
.A3(n_30),
.B1(n_36),
.B2(n_20),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_32),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_18),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_29),
.B1(n_16),
.B2(n_19),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_60),
.B1(n_25),
.B2(n_19),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_76),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_59),
.B1(n_32),
.B2(n_25),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_99),
.B1(n_103),
.B2(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_29),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_105),
.CI(n_82),
.CON(n_128),
.SN(n_128)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_82),
.B(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_14),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_0),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_3),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_81),
.C(n_70),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_118),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_123),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_96),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_70),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_133),
.B1(n_106),
.B2(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_81),
.C(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_96),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_147),
.B1(n_152),
.B2(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_106),
.B(n_103),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_150),
.B(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_104),
.B1(n_103),
.B2(n_99),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_123),
.B1(n_97),
.B2(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_95),
.B(n_105),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_107),
.B(n_102),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_91),
.B1(n_108),
.B2(n_89),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_124),
.B1(n_98),
.B2(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_138),
.B1(n_137),
.B2(n_141),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_131),
.C(n_129),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_90),
.C(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_135),
.C(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_98),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_165),
.B(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_86),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_86),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_146),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_176),
.Y(n_182)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_157),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_173),
.B(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_3),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_164),
.B(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_160),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_154),
.B(n_156),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_181),
.B1(n_169),
.B2(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_165),
.B1(n_180),
.B2(n_178),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_185),
.B(n_182),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_187),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.C(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_200),
.C(n_7),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_200),
.B(n_7),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);


endmodule