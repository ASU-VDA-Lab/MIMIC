module fake_netlist_6_762_n_1529 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1529);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1529;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_SL g145 ( 
.A(n_16),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_53),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_46),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_8),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_31),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_25),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_38),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_20),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_99),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_85),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_15),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_92),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_130),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx8_ASAP7_75t_SL g171 ( 
.A(n_31),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_12),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_30),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_47),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_64),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_1),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_42),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_35),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_29),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_50),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_68),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_13),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_67),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_28),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_20),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_37),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_84),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_59),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_30),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_97),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_43),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_13),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_39),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_61),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_132),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_24),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_79),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_66),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_81),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_1),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_123),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_75),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_6),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_37),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_44),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_46),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_122),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_126),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_6),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_26),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_103),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_49),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_91),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_136),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_2),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_114),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_18),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_116),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_72),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_14),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_17),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_40),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_77),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_60),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_96),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_78),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_69),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_21),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_113),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_102),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_29),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_86),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_10),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_265),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_171),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_151),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_187),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_151),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_151),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_187),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_204),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_204),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_204),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_221),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_225),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_171),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_204),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_245),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_147),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_251),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_204),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_167),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

INVx4_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_181),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_233),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_150),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_233),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_233),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_185),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_156),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_284),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_174),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_175),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_198),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_188),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_263),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_223),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_155),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_263),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_172),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_155),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_279),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_279),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_195),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_146),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_268),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_191),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_148),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_148),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_203),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_234),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_292),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_219),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_168),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_356),
.B(n_202),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_295),
.B(n_168),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_311),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_312),
.A2(n_241),
.B1(n_202),
.B2(n_145),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_R g381 ( 
.A(n_311),
.B(n_320),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_321),
.B(n_153),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_296),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_296),
.B(n_170),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_290),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_291),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_298),
.A2(n_196),
.B(n_179),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_297),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_179),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_300),
.B(n_196),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_326),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_302),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_294),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_276),
.B(n_226),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_361),
.B(n_330),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_309),
.B(n_306),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_153),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_154),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_330),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_309),
.B(n_226),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_313),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_337),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_299),
.A2(n_241),
.B1(n_285),
.B2(n_283),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_316),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_350),
.B(n_157),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_249),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_297),
.B(n_146),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_317),
.B(n_154),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_317),
.B(n_276),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_301),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_167),
.Y(n_430)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_374),
.B(n_167),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_420),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_381),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_365),
.B(n_359),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_363),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_364),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_374),
.B(n_167),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_359),
.B1(n_249),
.B2(n_346),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_374),
.A2(n_325),
.B1(n_176),
.B2(n_336),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_325),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_420),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_392),
.B(n_331),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_405),
.B(n_352),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_289),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_404),
.A2(n_166),
.B(n_163),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_418),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_374),
.B(n_186),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_405),
.B(n_186),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_385),
.B(n_186),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_391),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_377),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_385),
.B(n_186),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_385),
.B(n_333),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_375),
.B(n_328),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_371),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_370),
.B(n_289),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_385),
.B(n_217),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_393),
.B(n_334),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_402),
.B(n_324),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_369),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_375),
.B(n_329),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_397),
.B(n_201),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_378),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_370),
.B(n_308),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_369),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_393),
.B(n_217),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_399),
.Y(n_497)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

INVx11_ASAP7_75t_L g499 ( 
.A(n_373),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_406),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_393),
.B(n_217),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_414),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_308),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_394),
.A2(n_335),
.B1(n_340),
.B2(n_338),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_415),
.B(n_305),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_419),
.B(n_357),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_394),
.B(n_217),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_394),
.B(n_286),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_390),
.B(n_426),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_369),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_394),
.B(n_286),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_409),
.B(n_307),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_380),
.B(n_157),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

OAI22xp33_ASAP7_75t_L g526 ( 
.A1(n_373),
.A2(n_180),
.B1(n_215),
.B2(n_208),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_428),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_411),
.B(n_310),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_387),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_380),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_369),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_376),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_240),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_388),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_412),
.B(n_339),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_149),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_407),
.B(n_286),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_343),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_388),
.B(n_286),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_376),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_407),
.B(n_173),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_407),
.B(n_177),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_388),
.B(n_178),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_413),
.B(n_357),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_390),
.B(n_152),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_376),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_390),
.B(n_348),
.Y(n_553)
);

AO21x2_ASAP7_75t_L g554 ( 
.A1(n_389),
.A2(n_224),
.B(n_190),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_388),
.B(n_183),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_422),
.A2(n_351),
.B1(n_353),
.B2(n_280),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_395),
.B(n_164),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_396),
.B(n_165),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_376),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_396),
.B(n_349),
.Y(n_561)
);

INVxp33_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_396),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_422),
.B(n_261),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_379),
.B(n_169),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_425),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_564),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_473),
.A2(n_403),
.B(n_400),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_454),
.B(n_351),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_434),
.B(n_158),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_449),
.B(n_403),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_453),
.B(n_158),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_522),
.B(n_425),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_522),
.B(n_425),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_438),
.B(n_425),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_437),
.B(n_358),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_159),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_425),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_560),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_427),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_491),
.B(n_358),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_454),
.B(n_353),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_432),
.B(n_427),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_455),
.B(n_159),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_489),
.A2(n_227),
.B1(n_206),
.B2(n_200),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_435),
.B(n_427),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_441),
.B(n_427),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_442),
.B(n_427),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_448),
.B(n_450),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_459),
.B(n_427),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_462),
.B(n_429),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_454),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_463),
.B(n_467),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_446),
.B(n_161),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_429),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_492),
.B(n_160),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_561),
.B(n_160),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_477),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_475),
.B(n_429),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_494),
.B(n_429),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_429),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_523),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_443),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_451),
.B(n_344),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_505),
.B(n_429),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_458),
.A2(n_214),
.B1(n_197),
.B2(n_194),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_447),
.B(n_162),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_379),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_528),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_477),
.B(n_345),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_460),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_489),
.A2(n_400),
.B1(n_389),
.B2(n_252),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_532),
.B(n_379),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_446),
.B(n_345),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_553),
.A2(n_216),
.B1(n_184),
.B2(n_192),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_485),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_541),
.B(n_379),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_506),
.B(n_189),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_SL g626 ( 
.A(n_497),
.B(n_161),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_542),
.B(n_400),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_465),
.B(n_282),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_210),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_513),
.B(n_199),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_461),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_478),
.B(n_488),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_517),
.B(n_400),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_510),
.B(n_211),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_499),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_461),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_521),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_540),
.A2(n_218),
.B1(n_274),
.B2(n_273),
.Y(n_639)
);

AND2x6_ASAP7_75t_SL g640 ( 
.A(n_534),
.B(n_347),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_465),
.B(n_193),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_474),
.B(n_205),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_524),
.A2(n_253),
.B1(n_256),
.B2(n_270),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_445),
.B(n_490),
.C(n_564),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_538),
.A2(n_209),
.B1(n_272),
.B2(n_266),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_486),
.B(n_213),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_486),
.A2(n_207),
.B1(n_264),
.B2(n_262),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_466),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_512),
.B(n_426),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_536),
.B(n_222),
.Y(n_651)
);

OAI221xp5_ASAP7_75t_L g652 ( 
.A1(n_556),
.A2(n_524),
.B1(n_507),
.B2(n_547),
.C(n_546),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_486),
.B(n_526),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_481),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_486),
.A2(n_254),
.B1(n_228),
.B2(n_232),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_536),
.Y(n_656)
);

O2A1O1Ixp5_ASAP7_75t_L g657 ( 
.A1(n_471),
.A2(n_347),
.B(n_318),
.C(n_146),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_557),
.B(n_376),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_549),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_527),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_498),
.A2(n_248),
.B1(n_231),
.B2(n_235),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_464),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_558),
.B(n_382),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_529),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_471),
.A2(n_239),
.B(n_242),
.C(n_255),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_464),
.B(n_382),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_498),
.B(n_382),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_550),
.B(n_382),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_565),
.B(n_382),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_500),
.B(n_257),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_500),
.B(n_509),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_527),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_547),
.B(n_260),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_433),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_481),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_433),
.B(n_278),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_444),
.B(n_212),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_452),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_530),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_468),
.B(n_267),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_468),
.B(n_212),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_452),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_530),
.B(n_259),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_452),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_482),
.B(n_258),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_534),
.B(n_212),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_SL g687 ( 
.A1(n_534),
.A2(n_250),
.B1(n_247),
.B2(n_246),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_543),
.B(n_243),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_472),
.A2(n_237),
.B1(n_236),
.B2(n_230),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_452),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_472),
.B(n_135),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_534),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_554),
.A2(n_238),
.B1(n_229),
.B2(n_4),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_501),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_430),
.A2(n_134),
.B1(n_124),
.B2(n_117),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_503),
.B(n_108),
.Y(n_697)
);

NAND2x1p5_ASAP7_75t_L g698 ( 
.A(n_476),
.B(n_88),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_476),
.A2(n_496),
.B(n_516),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_504),
.B(n_87),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_SL g701 ( 
.A(n_493),
.B(n_0),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_554),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_508),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_439),
.B(n_3),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_430),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_493),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_511),
.B(n_76),
.Y(n_707)
);

AND3x1_ASAP7_75t_SL g708 ( 
.A(n_580),
.B(n_7),
.C(n_9),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_633),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_578),
.B(n_519),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_607),
.B(n_496),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_569),
.A2(n_627),
.B(n_669),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_585),
.B(n_519),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_594),
.B(n_567),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_615),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_597),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_656),
.B(n_515),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_585),
.B(n_601),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_SL g721 ( 
.A(n_601),
.B(n_516),
.C(n_539),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_656),
.B(n_691),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_607),
.B(n_539),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_656),
.B(n_515),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_602),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_656),
.B(n_566),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_614),
.B(n_520),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_603),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_674),
.B(n_551),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_621),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_678),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_SL g732 ( 
.A(n_653),
.B(n_520),
.C(n_16),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_619),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_582),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_678),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_660),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_622),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_656),
.B(n_439),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_694),
.A2(n_484),
.B1(n_502),
.B2(n_514),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_609),
.Y(n_741)
);

BUFx4f_ASAP7_75t_L g742 ( 
.A(n_631),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_678),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_672),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_609),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_570),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_614),
.B(n_11),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_645),
.Y(n_749)
);

AND2x6_ASAP7_75t_SL g750 ( 
.A(n_683),
.B(n_17),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_682),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_635),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_664),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_682),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_694),
.A2(n_514),
.B1(n_502),
.B2(n_484),
.Y(n_755)
);

BUFx4f_ASAP7_75t_L g756 ( 
.A(n_631),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_691),
.B(n_535),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_616),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_572),
.B(n_559),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_629),
.B(n_440),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_586),
.A2(n_555),
.B(n_548),
.C(n_544),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_596),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_702),
.A2(n_514),
.B1(n_484),
.B2(n_502),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_576),
.B(n_440),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_682),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_603),
.B(n_439),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_480),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_642),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_644),
.A2(n_555),
.B1(n_548),
.B2(n_470),
.Y(n_769)
);

AND2x6_ASAP7_75t_SL g770 ( 
.A(n_631),
.B(n_19),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_687),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_659),
.B(n_470),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_570),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_583),
.B(n_552),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_583),
.B(n_552),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_632),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_702),
.A2(n_514),
.B1(n_484),
.B2(n_502),
.Y(n_777)
);

AO22x1_ASAP7_75t_L g778 ( 
.A1(n_647),
.A2(n_502),
.B1(n_484),
.B2(n_514),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_659),
.B(n_22),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_679),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_552),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_634),
.A2(n_545),
.B(n_533),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_635),
.B(n_545),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_637),
.Y(n_784)
);

BUFx12f_ASAP7_75t_SL g785 ( 
.A(n_671),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_705),
.A2(n_544),
.B1(n_545),
.B2(n_533),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_684),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_705),
.A2(n_533),
.B1(n_456),
.B2(n_518),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_684),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_636),
.B(n_518),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_568),
.B(n_518),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_693),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_568),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_684),
.Y(n_794)
);

OR2x2_ASAP7_75t_SL g795 ( 
.A(n_593),
.B(n_23),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_649),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_652),
.A2(n_457),
.B1(n_480),
.B2(n_531),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_703),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_679),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_690),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_695),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_652),
.A2(n_457),
.B1(n_531),
.B2(n_493),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_571),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_593),
.Y(n_804)
);

NOR2x1p5_ASAP7_75t_L g805 ( 
.A(n_676),
.B(n_531),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_600),
.B(n_487),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_688),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_630),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_579),
.B(n_487),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_573),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_690),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_599),
.B(n_23),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_581),
.B(n_487),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_577),
.B(n_24),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_685),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_643),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_688),
.B(n_479),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_643),
.B(n_57),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_686),
.B(n_33),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_625),
.B(n_479),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_654),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_675),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_600),
.B(n_479),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_630),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_680),
.Y(n_825)
);

CKINVDCx8_ASAP7_75t_R g826 ( 
.A(n_640),
.Y(n_826)
);

AND2x6_ASAP7_75t_SL g827 ( 
.A(n_704),
.B(n_33),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_613),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

NOR2x2_ASAP7_75t_L g830 ( 
.A(n_662),
.B(n_34),
.Y(n_830)
);

NOR2x2_ASAP7_75t_L g831 ( 
.A(n_662),
.B(n_34),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_617),
.B(n_574),
.Y(n_832)
);

BUFx12f_ASAP7_75t_SL g833 ( 
.A(n_626),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_617),
.B(n_479),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_677),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_655),
.B(n_35),
.C(n_41),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_628),
.B(n_42),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_575),
.B(n_611),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_699),
.B(n_431),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_623),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_692),
.B(n_62),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_699),
.B(n_431),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_681),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_620),
.B(n_431),
.Y(n_844)
);

CKINVDCx11_ASAP7_75t_R g845 ( 
.A(n_689),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_584),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_587),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_690),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_670),
.B(n_44),
.Y(n_849)
);

NOR2x1p5_ASAP7_75t_L g850 ( 
.A(n_666),
.B(n_591),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_588),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_706),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_589),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_639),
.B(n_431),
.C(n_436),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_692),
.A2(n_45),
.B1(n_71),
.B2(n_74),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_592),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_648),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_612),
.B(n_436),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_706),
.B(n_436),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_701),
.A2(n_45),
.B1(n_436),
.B2(n_698),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_641),
.B(n_651),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_598),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_604),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_673),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_657),
.B(n_661),
.C(n_665),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_646),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_605),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_720),
.A2(n_650),
.B1(n_667),
.B2(n_698),
.Y(n_868)
);

BUFx6f_ASAP7_75t_SL g869 ( 
.A(n_780),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_722),
.A2(n_668),
.B(n_663),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_752),
.B(n_606),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_832),
.A2(n_610),
.B(n_658),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_752),
.A2(n_657),
.B(n_697),
.C(n_700),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_740),
.B(n_755),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_807),
.B(n_762),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_712),
.B(n_707),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_793),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_818),
.B(n_696),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_723),
.B(n_815),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_812),
.A2(n_819),
.B(n_849),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_785),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_746),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_818),
.A2(n_757),
.B1(n_755),
.B2(n_740),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_709),
.B(n_734),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_731),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_731),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_709),
.B(n_866),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_749),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_804),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_793),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_763),
.A2(n_777),
.B1(n_727),
.B2(n_802),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_812),
.A2(n_849),
.B(n_819),
.C(n_772),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_731),
.Y(n_893)
);

BUFx2_ASAP7_75t_SL g894 ( 
.A(n_736),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_748),
.A2(n_816),
.B(n_779),
.C(n_732),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_816),
.A2(n_732),
.B(n_836),
.C(n_814),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_728),
.A2(n_738),
.B(n_760),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_731),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_782),
.A2(n_797),
.B(n_838),
.Y(n_899)
);

XNOR2xp5_ASAP7_75t_L g900 ( 
.A(n_857),
.B(n_768),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_808),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_764),
.A2(n_724),
.B(n_719),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_837),
.A2(n_718),
.B1(n_737),
.B2(n_730),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_772),
.A2(n_810),
.B(n_803),
.C(n_825),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_735),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_824),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_861),
.A2(n_783),
.B(n_725),
.C(n_739),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_846),
.B(n_847),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_721),
.A2(n_840),
.B1(n_828),
.B2(n_829),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_851),
.B(n_853),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_747),
.B(n_773),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_711),
.Y(n_912)
);

INVx8_ASAP7_75t_L g913 ( 
.A(n_735),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_745),
.B(n_716),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_856),
.B(n_862),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_836),
.A2(n_729),
.B(n_721),
.C(n_753),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_744),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_834),
.A2(n_766),
.B(n_710),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_SL g919 ( 
.A(n_771),
.B(n_717),
.C(n_790),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_795),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_741),
.B(n_864),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_735),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_863),
.B(n_867),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_742),
.B(n_756),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_763),
.A2(n_777),
.B(n_761),
.C(n_860),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_860),
.A2(n_714),
.B1(n_786),
.B2(n_788),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_726),
.A2(n_817),
.B(n_781),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_767),
.A2(n_713),
.B(n_842),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_751),
.B(n_794),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_790),
.B(n_774),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_845),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_839),
.A2(n_809),
.B(n_813),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_774),
.B(n_775),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_835),
.A2(n_843),
.B1(n_775),
.B2(n_841),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_786),
.A2(n_788),
.B1(n_850),
.B2(n_765),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_799),
.B(n_841),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_833),
.B(n_791),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_742),
.B(n_756),
.Y(n_938)
);

OAI22x1_ASAP7_75t_L g939 ( 
.A1(n_830),
.A2(n_831),
.B1(n_805),
.B2(n_791),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_715),
.B(n_858),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_735),
.B(n_787),
.Y(n_941)
);

OAI22x1_ASAP7_75t_L g942 ( 
.A1(n_769),
.A2(n_827),
.B1(n_708),
.B2(n_770),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_SL g943 ( 
.A(n_855),
.B(n_826),
.C(n_865),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_750),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_792),
.B(n_798),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_787),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_761),
.A2(n_865),
.B(n_822),
.C(n_801),
.Y(n_947)
);

BUFx10_ASAP7_75t_L g948 ( 
.A(n_858),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_758),
.A2(n_784),
.B(n_821),
.C(n_796),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_787),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_787),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_776),
.B(n_848),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_789),
.B(n_811),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_743),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_743),
.B(n_754),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_754),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_855),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_844),
.A2(n_806),
.B(n_823),
.C(n_859),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_854),
.A2(n_806),
.B(n_820),
.C(n_852),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_789),
.B(n_811),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_751),
.B(n_794),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_789),
.Y(n_962)
);

AO32x1_ASAP7_75t_L g963 ( 
.A1(n_708),
.A2(n_800),
.A3(n_759),
.B1(n_778),
.B2(n_859),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_SL g964 ( 
.A1(n_800),
.A2(n_789),
.B1(n_811),
.B2(n_759),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_811),
.B(n_759),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_759),
.A2(n_720),
.B(n_653),
.C(n_812),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_759),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_SL g968 ( 
.A1(n_720),
.A2(n_586),
.B(n_807),
.C(n_752),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_722),
.A2(n_603),
.B(n_498),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_752),
.B(n_807),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_720),
.A2(n_807),
.B1(n_722),
.B2(n_752),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_752),
.B(n_607),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_733),
.B(n_633),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_746),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_720),
.A2(n_807),
.B1(n_722),
.B2(n_752),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_768),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_720),
.B(n_752),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_720),
.A2(n_653),
.B(n_752),
.C(n_812),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_722),
.A2(n_603),
.B(n_498),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_752),
.B(n_807),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_731),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_720),
.A2(n_653),
.B(n_812),
.C(n_578),
.Y(n_982)
);

AND3x1_ASAP7_75t_SL g983 ( 
.A(n_830),
.B(n_831),
.C(n_745),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_722),
.A2(n_603),
.B(n_498),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_720),
.A2(n_807),
.B1(n_722),
.B2(n_752),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_746),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_768),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_720),
.A2(n_653),
.B(n_812),
.C(n_578),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_899),
.A2(n_870),
.B(n_927),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_882),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_977),
.B(n_982),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_988),
.A2(n_968),
.B(n_892),
.Y(n_992)
);

BUFx2_ASAP7_75t_SL g993 ( 
.A(n_869),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_928),
.A2(n_932),
.B(n_902),
.Y(n_994)
);

NOR4xp25_ASAP7_75t_L g995 ( 
.A(n_880),
.B(n_978),
.C(n_943),
.D(n_896),
.Y(n_995)
);

OAI21x1_ASAP7_75t_SL g996 ( 
.A1(n_958),
.A2(n_909),
.B(n_916),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_955),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_872),
.A2(n_897),
.B(n_868),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_888),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_973),
.B(n_972),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_976),
.B(n_987),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_966),
.A2(n_925),
.B(n_926),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_917),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_940),
.B(n_936),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_908),
.B(n_910),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_878),
.A2(n_895),
.B(n_883),
.C(n_907),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_893),
.B(n_905),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_969),
.A2(n_984),
.B(n_979),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_876),
.A2(n_873),
.B(n_891),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_SL g1010 ( 
.A(n_935),
.B(n_915),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_909),
.A2(n_904),
.B(n_975),
.C(n_971),
.Y(n_1011)
);

OAI21xp33_ASAP7_75t_L g1012 ( 
.A1(n_903),
.A2(n_879),
.B(n_957),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_894),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_930),
.A2(n_965),
.B(n_952),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_940),
.B(n_936),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_913),
.B(n_936),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_941),
.A2(n_953),
.B(n_985),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_875),
.B(n_970),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_900),
.B(n_937),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_874),
.A2(n_959),
.B(n_923),
.Y(n_1020)
);

AOI221x1_ASAP7_75t_L g1021 ( 
.A1(n_942),
.A2(n_939),
.B1(n_964),
.B2(n_967),
.C(n_945),
.Y(n_1021)
);

BUFx2_ASAP7_75t_R g1022 ( 
.A(n_924),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_980),
.B(n_887),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_871),
.A2(n_933),
.B(n_949),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_919),
.B(n_884),
.C(n_921),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_974),
.A2(n_986),
.B(n_934),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_946),
.A2(n_950),
.B(n_981),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_954),
.A2(n_956),
.B(n_962),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_L g1029 ( 
.A(n_960),
.B(n_913),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_913),
.A2(n_963),
.B(n_961),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_877),
.B(n_906),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_SL g1032 ( 
.A1(n_920),
.A2(n_938),
.B(n_914),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_950),
.A2(n_981),
.B(n_929),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_931),
.A2(n_911),
.B1(n_881),
.B2(n_983),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_911),
.B(n_889),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_912),
.B(n_890),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_948),
.A2(n_893),
.B(n_905),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_948),
.A2(n_951),
.B(n_885),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_901),
.B(n_885),
.C(n_886),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_885),
.A2(n_886),
.B(n_898),
.C(n_922),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_886),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_944),
.A2(n_898),
.B(n_922),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_922),
.A2(n_951),
.B(n_869),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_897),
.A2(n_918),
.B(n_928),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_917),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_880),
.A2(n_720),
.B(n_988),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_928),
.A2(n_947),
.A3(n_932),
.B(n_966),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_880),
.A2(n_629),
.B(n_653),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_877),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_928),
.A2(n_932),
.B(n_902),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_880),
.B(n_607),
.Y(n_1051)
);

AO31x2_ASAP7_75t_L g1052 ( 
.A1(n_928),
.A2(n_947),
.A3(n_932),
.B(n_966),
.Y(n_1052)
);

NAND2x1p5_ASAP7_75t_L g1053 ( 
.A(n_893),
.B(n_905),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_894),
.B(n_913),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_SL g1055 ( 
.A1(n_971),
.A2(n_586),
.B(n_985),
.C(n_975),
.Y(n_1055)
);

AO31x2_ASAP7_75t_L g1056 ( 
.A1(n_928),
.A2(n_947),
.A3(n_932),
.B(n_966),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_977),
.B(n_752),
.Y(n_1057)
);

NOR4xp25_ASAP7_75t_L g1058 ( 
.A(n_880),
.B(n_988),
.C(n_982),
.D(n_892),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_977),
.B(n_752),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_SL g1060 ( 
.A1(n_958),
.A2(n_909),
.B(n_916),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_SL g1061 ( 
.A1(n_977),
.A2(n_720),
.B(n_861),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_977),
.B(n_752),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_SL g1063 ( 
.A1(n_977),
.A2(n_720),
.B(n_861),
.Y(n_1063)
);

AO32x2_ASAP7_75t_L g1064 ( 
.A1(n_926),
.A2(n_985),
.A3(n_975),
.B1(n_971),
.B2(n_935),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_889),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_977),
.B(n_752),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_973),
.B(n_633),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_880),
.A2(n_943),
.B1(n_653),
.B2(n_878),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_925),
.A2(n_818),
.B1(n_926),
.B2(n_740),
.Y(n_1069)
);

INVx8_ASAP7_75t_L g1070 ( 
.A(n_913),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_L g1071 ( 
.A1(n_982),
.A2(n_720),
.B(n_988),
.C(n_892),
.Y(n_1071)
);

AO21x2_ASAP7_75t_L g1072 ( 
.A1(n_899),
.A2(n_928),
.B(n_932),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_899),
.A2(n_928),
.B(n_947),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_982),
.A2(n_988),
.B(n_899),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_882),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_977),
.B(n_752),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_880),
.B(n_752),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_917),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_882),
.Y(n_1079)
);

AOI221x1_ASAP7_75t_L g1080 ( 
.A1(n_880),
.A2(n_988),
.B1(n_982),
.B2(n_892),
.C(n_943),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_982),
.A2(n_988),
.B(n_899),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_977),
.B(n_752),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_982),
.A2(n_988),
.B(n_899),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_885),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_973),
.B(n_633),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_882),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_982),
.A2(n_988),
.B(n_899),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_977),
.B(n_982),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_928),
.A2(n_947),
.A3(n_932),
.B(n_966),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_925),
.A2(n_818),
.B1(n_926),
.B2(n_740),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_894),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_894),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_973),
.B(n_633),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_977),
.B(n_752),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_928),
.A2(n_947),
.A3(n_932),
.B(n_966),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_977),
.B(n_752),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_877),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_917),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_977),
.B(n_752),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_977),
.B(n_752),
.Y(n_1100)
);

CKINVDCx11_ASAP7_75t_R g1101 ( 
.A(n_931),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1048),
.B(n_991),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1008),
.A2(n_1050),
.B(n_994),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_990),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_997),
.B(n_1004),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_999),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1003),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_998),
.B(n_1074),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1051),
.B(n_1012),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_989),
.A2(n_1009),
.B(n_992),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1068),
.A2(n_1046),
.B1(n_1087),
.B2(n_1074),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_1070),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1081),
.A2(n_1087),
.B(n_1083),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_1037),
.B(n_1038),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1046),
.A2(n_1020),
.B(n_1055),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1005),
.A2(n_1025),
.B1(n_1018),
.B2(n_1059),
.Y(n_1116)
);

CKINVDCx11_ASAP7_75t_R g1117 ( 
.A(n_1101),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1013),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_R g1119 ( 
.A(n_1070),
.B(n_1029),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_1001),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1006),
.A2(n_1069),
.B(n_1090),
.C(n_1002),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1075),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1079),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_996),
.A2(n_1060),
.B(n_1002),
.Y(n_1124)
);

BUFx5_ASAP7_75t_L g1125 ( 
.A(n_1086),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1000),
.B(n_1067),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_997),
.B(n_1004),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1033),
.B(n_1027),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1084),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1085),
.B(n_1093),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1058),
.A2(n_1024),
.B(n_1088),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1010),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1078),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1005),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1028),
.Y(n_1135)
);

OAI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_995),
.A2(n_1025),
.B1(n_1032),
.B2(n_1034),
.C(n_1023),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1084),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1069),
.A2(n_1090),
.B1(n_1077),
.B2(n_1088),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1057),
.A2(n_1100),
.B1(n_1062),
.B2(n_1066),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_1072),
.A2(n_1011),
.B(n_1030),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1076),
.B(n_1099),
.Y(n_1141)
);

AO221x2_ASAP7_75t_L g1142 ( 
.A1(n_1032),
.A2(n_995),
.B1(n_1026),
.B2(n_1042),
.C(n_1021),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_993),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_1063),
.B(n_1061),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1098),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1026),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1073),
.A2(n_1014),
.B(n_1040),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1043),
.A2(n_1007),
.B(n_1053),
.Y(n_1148)
);

BUFx2_ASAP7_75t_SL g1149 ( 
.A(n_1065),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1036),
.Y(n_1150)
);

AOI332xp33_ASAP7_75t_L g1151 ( 
.A1(n_1082),
.A2(n_1094),
.A3(n_1096),
.B1(n_1015),
.B2(n_1041),
.B3(n_1064),
.C1(n_1049),
.C2(n_1022),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1098),
.A2(n_1097),
.B1(n_1045),
.B2(n_1092),
.C(n_1091),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1015),
.A2(n_1054),
.B1(n_1042),
.B2(n_1016),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1039),
.A2(n_1019),
.B(n_1031),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1039),
.A2(n_1035),
.B(n_1054),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1047),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1064),
.A2(n_1016),
.B1(n_1084),
.B2(n_1052),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1047),
.A2(n_1052),
.A3(n_1056),
.B(n_1089),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1016),
.A2(n_1064),
.B(n_1052),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1095),
.A2(n_1056),
.B(n_1089),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1056),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1089),
.A2(n_1008),
.B(n_1044),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1095),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1037),
.B(n_967),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1037),
.B(n_967),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1048),
.A2(n_880),
.B(n_629),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_990),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_1067),
.Y(n_1168)
);

AND2x6_ASAP7_75t_L g1169 ( 
.A(n_1088),
.B(n_965),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1000),
.B(n_1067),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_992),
.A2(n_998),
.B(n_1074),
.Y(n_1171)
);

BUFx2_ASAP7_75t_SL g1172 ( 
.A(n_1003),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1003),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1098),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1069),
.A2(n_818),
.B1(n_299),
.B2(n_301),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1008),
.A2(n_1044),
.B(n_994),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1048),
.B(n_880),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1003),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1008),
.A2(n_1050),
.B(n_994),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_990),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1048),
.A2(n_880),
.B1(n_1068),
.B2(n_653),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1071),
.A2(n_720),
.B(n_982),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1071),
.A2(n_720),
.B(n_982),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_990),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1008),
.A2(n_1050),
.B(n_994),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_992),
.A2(n_998),
.B(n_1074),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_992),
.A2(n_998),
.B(n_1074),
.Y(n_1188)
);

BUFx2_ASAP7_75t_SL g1189 ( 
.A(n_1003),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_990),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_998),
.A2(n_1080),
.A3(n_989),
.B(n_1011),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1098),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1068),
.A2(n_607),
.B1(n_614),
.B2(n_720),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_990),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1003),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1048),
.A2(n_880),
.B(n_818),
.C(n_982),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1005),
.B(n_1094),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1048),
.A2(n_880),
.B1(n_1068),
.B2(n_653),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1048),
.A2(n_880),
.B1(n_1068),
.B2(n_653),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1068),
.A2(n_607),
.B1(n_614),
.B2(n_720),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1003),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1107),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1175),
.A2(n_1139),
.B1(n_1199),
.B2(n_1198),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1175),
.A2(n_1166),
.B(n_1177),
.C(n_1109),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1170),
.B(n_1130),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1141),
.B(n_1139),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1181),
.A2(n_1199),
.B1(n_1198),
.B2(n_1136),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1173),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1178),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1195),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1105),
.B(n_1127),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1134),
.B(n_1197),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1154),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1105),
.B(n_1127),
.Y(n_1214)
);

AND2x6_ASAP7_75t_L g1215 ( 
.A(n_1146),
.B(n_1163),
.Y(n_1215)
);

OA22x2_ASAP7_75t_L g1216 ( 
.A1(n_1116),
.A2(n_1155),
.B1(n_1200),
.B2(n_1193),
.Y(n_1216)
);

INVx8_ASAP7_75t_L g1217 ( 
.A(n_1118),
.Y(n_1217)
);

NAND2x1_ASAP7_75t_L g1218 ( 
.A(n_1169),
.B(n_1135),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1115),
.A2(n_1131),
.B(n_1160),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1124),
.B(n_1138),
.Y(n_1220)
);

AND2x6_ASAP7_75t_L g1221 ( 
.A(n_1156),
.B(n_1161),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_1121),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1111),
.A2(n_1196),
.B1(n_1153),
.B2(n_1121),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1124),
.B(n_1138),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1145),
.B(n_1174),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1117),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1162),
.A2(n_1147),
.B(n_1144),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1153),
.B(n_1148),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1142),
.A2(n_1151),
.B(n_1113),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1150),
.B(n_1104),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_1117),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1192),
.B(n_1122),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1142),
.A2(n_1113),
.B(n_1132),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1110),
.A2(n_1171),
.B(n_1186),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1106),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1177),
.A2(n_1152),
.B1(n_1132),
.B2(n_1143),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1133),
.B(n_1201),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1191),
.A2(n_1188),
.B(n_1186),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1123),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1172),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1102),
.B(n_1169),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1167),
.B(n_1194),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1143),
.A2(n_1120),
.B1(n_1189),
.B2(n_1157),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1180),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1184),
.B(n_1190),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1120),
.A2(n_1157),
.B1(n_1149),
.B2(n_1118),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1187),
.A2(n_1188),
.B1(n_1108),
.B2(n_1171),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1112),
.A2(n_1137),
.B1(n_1129),
.B2(n_1159),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1169),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_1119),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1169),
.B(n_1125),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1164),
.A2(n_1165),
.B1(n_1114),
.B2(n_1128),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1140),
.B(n_1125),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1114),
.A2(n_1164),
.B(n_1165),
.C(n_1128),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1125),
.B(n_1158),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1125),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1176),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1103),
.A2(n_1179),
.B(n_1185),
.Y(n_1258)
);

BUFx8_ASAP7_75t_SL g1259 ( 
.A(n_1118),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1175),
.A2(n_1068),
.B1(n_1139),
.B2(n_1025),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1196),
.A2(n_892),
.B(n_926),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1175),
.A2(n_880),
.B1(n_671),
.B2(n_653),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1175),
.A2(n_771),
.B1(n_819),
.B2(n_653),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1126),
.B(n_1168),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1219),
.B(n_1255),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1234),
.B(n_1253),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1218),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1257),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1241),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1247),
.B(n_1251),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1224),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1227),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1256),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1220),
.B(n_1224),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1241),
.B(n_1249),
.Y(n_1275)
);

INVx5_ASAP7_75t_SL g1276 ( 
.A(n_1228),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1261),
.B(n_1222),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1227),
.Y(n_1278)
);

BUFx2_ASAP7_75t_R g1279 ( 
.A(n_1259),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1215),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1206),
.B(n_1212),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1221),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1249),
.A2(n_1239),
.B(n_1235),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1215),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1252),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1212),
.B(n_1223),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1204),
.B(n_1207),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1258),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1244),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1242),
.B(n_1214),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1232),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1248),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1238),
.A2(n_1213),
.B(n_1233),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1254),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1254),
.A2(n_1203),
.B(n_1260),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1246),
.A2(n_1243),
.B(n_1262),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1271),
.B(n_1230),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1291),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1283),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1268),
.B(n_1225),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1289),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1289),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1287),
.A2(n_1263),
.B1(n_1277),
.B2(n_1216),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1268),
.B(n_1210),
.Y(n_1304)
);

INVx5_ASAP7_75t_L g1305 ( 
.A(n_1277),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1288),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1273),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1283),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1283),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1265),
.B(n_1205),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1283),
.Y(n_1311)
);

OAI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1287),
.A2(n_1216),
.B1(n_1236),
.B2(n_1240),
.C(n_1208),
.Y(n_1312)
);

OAI222xp33_ASAP7_75t_L g1313 ( 
.A1(n_1287),
.A2(n_1229),
.B1(n_1250),
.B2(n_1245),
.C1(n_1226),
.C2(n_1264),
.Y(n_1313)
);

AND2x2_ASAP7_75t_SL g1314 ( 
.A(n_1284),
.B(n_1229),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1283),
.Y(n_1315)
);

AND2x4_ASAP7_75t_SL g1316 ( 
.A(n_1282),
.B(n_1211),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1266),
.B(n_1209),
.Y(n_1317)
);

AOI221xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1312),
.A2(n_1313),
.B1(n_1299),
.B2(n_1308),
.C(n_1315),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1314),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1309),
.A2(n_1278),
.B(n_1272),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1303),
.A2(n_1277),
.B1(n_1286),
.B2(n_1284),
.Y(n_1321)
);

OAI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1303),
.A2(n_1277),
.B1(n_1286),
.B2(n_1281),
.C(n_1292),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1301),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1312),
.A2(n_1277),
.B1(n_1296),
.B2(n_1295),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1304),
.B(n_1269),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1304),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1302),
.Y(n_1327)
);

OAI31xp33_ASAP7_75t_L g1328 ( 
.A1(n_1313),
.A2(n_1286),
.A3(n_1292),
.B(n_1285),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1316),
.B(n_1282),
.Y(n_1329)
);

OAI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1305),
.A2(n_1277),
.B1(n_1281),
.B2(n_1292),
.C(n_1269),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_L g1331 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1314),
.A2(n_1292),
.B(n_1284),
.C(n_1280),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_R g1333 ( 
.A(n_1298),
.B(n_1231),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1310),
.B(n_1276),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1314),
.A2(n_1277),
.B1(n_1295),
.B2(n_1296),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1298),
.Y(n_1336)
);

AND3x1_ASAP7_75t_L g1337 ( 
.A(n_1317),
.B(n_1279),
.C(n_1267),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1314),
.B(n_1290),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1305),
.A2(n_1296),
.B1(n_1295),
.B2(n_1285),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1305),
.A2(n_1296),
.B1(n_1295),
.B2(n_1275),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1307),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1297),
.B(n_1202),
.Y(n_1342)
);

NAND4xp25_ASAP7_75t_L g1343 ( 
.A(n_1300),
.B(n_1274),
.C(n_1270),
.D(n_1275),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_L g1344 ( 
.A(n_1308),
.B(n_1294),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1308),
.A2(n_1295),
.B1(n_1274),
.B2(n_1291),
.C(n_1275),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1320),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1343),
.B(n_1315),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1323),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_SL g1349 ( 
.A(n_1324),
.B(n_1315),
.C(n_1311),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1323),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1331),
.B(n_1305),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1320),
.Y(n_1352)
);

INVx4_ASAP7_75t_SL g1353 ( 
.A(n_1329),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_SL g1354 ( 
.A(n_1328),
.B(n_1279),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1319),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1344),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1331),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1329),
.Y(n_1358)
);

AND2x6_ASAP7_75t_SL g1359 ( 
.A(n_1333),
.B(n_1217),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1335),
.B(n_1324),
.C(n_1318),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1344),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1337),
.Y(n_1362)
);

INVx5_ASAP7_75t_L g1363 ( 
.A(n_1319),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1336),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_SL g1365 ( 
.A(n_1345),
.B(n_1309),
.C(n_1311),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1327),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1329),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1326),
.B(n_1306),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1341),
.B(n_1310),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1339),
.A2(n_1293),
.B(n_1294),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1352),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1352),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1347),
.B(n_1369),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1357),
.B(n_1334),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1362),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1359),
.B(n_1217),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1348),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1350),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1359),
.B(n_1217),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1353),
.B(n_1334),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1353),
.B(n_1358),
.Y(n_1381)
);

INVx5_ASAP7_75t_L g1382 ( 
.A(n_1355),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1352),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1347),
.B(n_1369),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1353),
.B(n_1319),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1365),
.B(n_1325),
.Y(n_1386)
);

AND2x2_ASAP7_75t_SL g1387 ( 
.A(n_1362),
.B(n_1337),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1338),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1352),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1366),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1365),
.B(n_1300),
.Y(n_1391)
);

NOR2x1_ASAP7_75t_SL g1392 ( 
.A(n_1349),
.B(n_1355),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1360),
.B(n_1327),
.Y(n_1393)
);

AND2x2_ASAP7_75t_SL g1394 ( 
.A(n_1354),
.B(n_1340),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1353),
.B(n_1329),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1346),
.Y(n_1396)
);

CKINVDCx14_ASAP7_75t_R g1397 ( 
.A(n_1355),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1356),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1353),
.B(n_1332),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1382),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1387),
.B(n_1358),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1379),
.B(n_1364),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1375),
.B(n_1364),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1387),
.B(n_1354),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1390),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1393),
.B(n_1360),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1387),
.B(n_1367),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1393),
.B(n_1349),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1375),
.B(n_1367),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1373),
.B(n_1368),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1375),
.B(n_1367),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1399),
.B(n_1367),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1398),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1399),
.B(n_1355),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1390),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_L g1416 ( 
.A1(n_1394),
.A2(n_1370),
.B(n_1322),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1399),
.B(n_1355),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1385),
.B(n_1355),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1394),
.A2(n_1295),
.B1(n_1321),
.B2(n_1296),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1394),
.A2(n_1370),
.B1(n_1363),
.B2(n_1330),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1398),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1395),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1382),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1388),
.B(n_1374),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1377),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1373),
.B(n_1368),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1377),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1395),
.B(n_1355),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1388),
.B(n_1342),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1380),
.B(n_1351),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1378),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1378),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1406),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1413),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1401),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1421),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1406),
.B(n_1374),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1402),
.B(n_1404),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1422),
.B(n_1380),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1401),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_SL g1444 ( 
.A(n_1400),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1407),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1424),
.B(n_1384),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1407),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1405),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1410),
.B(n_1384),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1415),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1428),
.B(n_1381),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1415),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1400),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1410),
.B(n_1386),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1418),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1433),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1433),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1409),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1444),
.A2(n_1408),
.B1(n_1419),
.B2(n_1420),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1456),
.B(n_1416),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1445),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1434),
.A2(n_1416),
.B1(n_1419),
.B2(n_1408),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1441),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1440),
.B(n_1376),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1454),
.A2(n_1423),
.B(n_1430),
.Y(n_1467)
);

OAI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1445),
.A2(n_1418),
.B(n_1417),
.Y(n_1468)
);

XOR2xp5_ASAP7_75t_L g1469 ( 
.A(n_1437),
.B(n_1428),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1436),
.B(n_1414),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1434),
.A2(n_1386),
.B1(n_1363),
.B2(n_1391),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1439),
.A2(n_1417),
.B(n_1414),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1443),
.A2(n_1431),
.B1(n_1412),
.B2(n_1411),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1452),
.Y(n_1476)
);

OAI21xp33_ASAP7_75t_L g1477 ( 
.A1(n_1446),
.A2(n_1431),
.B(n_1411),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1463),
.B(n_1435),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1474),
.B(n_1435),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1467),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1467),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1465),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1470),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1448),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_L g1488 ( 
.A1(n_1479),
.A2(n_1461),
.B(n_1471),
.C(n_1464),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1479),
.A2(n_1462),
.B(n_1464),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1487),
.A2(n_1477),
.B1(n_1473),
.B2(n_1469),
.C(n_1460),
.Y(n_1490)
);

AOI21xp33_ASAP7_75t_L g1491 ( 
.A1(n_1480),
.A2(n_1475),
.B(n_1455),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1481),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1486),
.A2(n_1452),
.B1(n_1459),
.B2(n_1455),
.Y(n_1493)
);

AOI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1478),
.A2(n_1459),
.B(n_1449),
.C(n_1453),
.Y(n_1494)
);

AOI222xp33_ASAP7_75t_L g1495 ( 
.A1(n_1482),
.A2(n_1392),
.B1(n_1453),
.B2(n_1451),
.C1(n_1449),
.C2(n_1442),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1484),
.A2(n_1451),
.B1(n_1442),
.B2(n_1458),
.C(n_1457),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1490),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1493),
.B(n_1485),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1492),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1489),
.A2(n_1483),
.B(n_1392),
.Y(n_1500)
);

XOR2xp5_ASAP7_75t_L g1501 ( 
.A(n_1491),
.B(n_1450),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1500),
.A2(n_1488),
.B(n_1495),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1501),
.B(n_1450),
.Y(n_1503)
);

NOR2x1_ASAP7_75t_L g1504 ( 
.A(n_1499),
.B(n_1457),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1498),
.B(n_1494),
.Y(n_1505)
);

NAND2xp33_ASAP7_75t_L g1506 ( 
.A(n_1497),
.B(n_1423),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1498),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1503),
.A2(n_1382),
.B1(n_1391),
.B2(n_1361),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1507),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1505),
.B(n_1496),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1504),
.Y(n_1511)
);

NAND4xp75_ASAP7_75t_L g1512 ( 
.A(n_1502),
.B(n_1458),
.C(n_1412),
.D(n_1381),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1511),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1509),
.B(n_1426),
.Y(n_1514)
);

NOR3x1_ASAP7_75t_L g1515 ( 
.A(n_1512),
.B(n_1506),
.C(n_1427),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1514),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1516),
.Y(n_1517)
);

XNOR2xp5_ASAP7_75t_L g1518 ( 
.A(n_1517),
.B(n_1513),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1517),
.A2(n_1510),
.B(n_1508),
.Y(n_1519)
);

XNOR2xp5_ASAP7_75t_L g1520 ( 
.A(n_1518),
.B(n_1515),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1519),
.A2(n_1432),
.B1(n_1427),
.B2(n_1425),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1520),
.A2(n_1432),
.B1(n_1425),
.B2(n_1430),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1521),
.A2(n_1430),
.B1(n_1426),
.B2(n_1382),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1522),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1524),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1525),
.A2(n_1523),
.B(n_1372),
.Y(n_1526)
);

AOI322xp5_ASAP7_75t_L g1527 ( 
.A1(n_1526),
.A2(n_1382),
.A3(n_1389),
.B1(n_1372),
.B2(n_1371),
.C1(n_1383),
.C2(n_1396),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1527),
.A2(n_1383),
.B1(n_1372),
.B2(n_1371),
.Y(n_1528)
);

AOI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1528),
.A2(n_1237),
.B(n_1383),
.C(n_1389),
.Y(n_1529)
);


endmodule