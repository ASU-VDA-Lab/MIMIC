module fake_jpeg_29494_n_156 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_18),
.B1(n_45),
.B2(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_64),
.B1(n_63),
.B2(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx2_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_71),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_63),
.B1(n_61),
.B2(n_4),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_55),
.B1(n_53),
.B2(n_52),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_91),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_57),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_61),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_1),
.CI(n_3),
.CON(n_98),
.SN(n_98)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_75),
.B1(n_61),
.B2(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_99),
.B1(n_106),
.B2(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_56),
.B1(n_68),
.B2(n_60),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_101),
.B1(n_110),
.B2(n_27),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_88),
.B1(n_90),
.B2(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_66),
.C(n_58),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_9),
.C(n_10),
.Y(n_127)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_51),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_20),
.B(n_43),
.Y(n_109)
);

NAND2x1p5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_9),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_19),
.B1(n_42),
.B2(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_16),
.B1(n_17),
.B2(n_28),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_106),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_12),
.C(n_13),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_47),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_139),
.B1(n_124),
.B2(n_117),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_30),
.B(n_34),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_127),
.B(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_144),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_146),
.B(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_148),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_130),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_149),
.B1(n_129),
.B2(n_142),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_136),
.B1(n_134),
.B2(n_132),
.Y(n_156)
);


endmodule