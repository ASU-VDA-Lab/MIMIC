module fake_jpeg_27990_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.C(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_16),
.B1(n_11),
.B2(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_22),
.B1(n_11),
.B2(n_16),
.Y(n_54)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_57),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_25),
.C(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_30),
.B1(n_27),
.B2(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_9),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_10),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_11),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_67),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_24),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_54),
.B1(n_50),
.B2(n_58),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_4),
.B(n_6),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_59),
.B(n_64),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_77),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_20),
.C(n_26),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_41),
.B1(n_57),
.B2(n_48),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_68),
.C(n_69),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_31),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_86),
.B(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_43),
.B1(n_44),
.B2(n_26),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_44),
.B1(n_31),
.B2(n_20),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_73),
.B1(n_78),
.B2(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_87),
.C(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_95),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_82),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_20),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_89),
.C(n_93),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_97),
.C(n_44),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_2),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_103),
.B(n_8),
.C(n_10),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.Y(n_107)
);


endmodule