module real_jpeg_22046_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_0),
.A2(n_31),
.B1(n_42),
.B2(n_50),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_0),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_2),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_2),
.A2(n_14),
.B(n_46),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_2),
.A2(n_42),
.B1(n_50),
.B2(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_78),
.B1(n_217),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_27),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_2),
.A2(n_27),
.B(n_244),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_132),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_132),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_3),
.A2(n_42),
.B1(n_50),
.B2(n_132),
.Y(n_251)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_5),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_158),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_158),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_5),
.A2(n_42),
.B1(n_50),
.B2(n_158),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_34),
.B1(n_42),
.B2(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_6),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_124)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_123),
.B(n_171),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_42),
.B1(n_50),
.B2(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_11),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_11),
.A2(n_42),
.B1(n_50),
.B2(n_164),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_164),
.Y(n_217)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_110),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_91),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_65),
.C(n_74),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_20),
.B(n_65),
.CI(n_74),
.CON(n_136),
.SN(n_136)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_21),
.A2(n_22),
.B1(n_93),
.B2(n_106),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_39),
.C(n_53),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_23),
.A2(n_28),
.B1(n_87),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_23),
.A2(n_87),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_23),
.B(n_162),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_23),
.A2(n_87),
.B1(n_131),
.B2(n_177),
.Y(n_288)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_25),
.B(n_30),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_24),
.B(n_89),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_24),
.A2(n_35),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_25),
.B(n_27),
.Y(n_168)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_36),
.B1(n_161),
.B2(n_168),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g243 ( 
.A1(n_26),
.A2(n_42),
.A3(n_57),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_56),
.Y(n_58)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g161 ( 
.A(n_30),
.B(n_162),
.CON(n_161),
.SN(n_161)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_39),
.A2(n_40),
.B1(n_98),
.B2(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_48),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_41),
.A2(n_44),
.B1(n_83),
.B2(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_41),
.A2(n_48),
.B(n_84),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_41),
.A2(n_44),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_41),
.A2(n_44),
.B1(n_213),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_41),
.A2(n_44),
.B1(n_235),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_41),
.A2(n_69),
.B(n_251),
.Y(n_266)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_44),
.A2(n_71),
.B(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_44),
.B(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_45),
.B(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_79),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_47),
.A2(n_50),
.B(n_162),
.C(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_70),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_50),
.B(n_56),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_60),
.B(n_63),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_54),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_54),
.A2(n_100),
.B(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_54),
.A2(n_63),
.B(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_55),
.A2(n_59),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_55),
.A2(n_59),
.B1(n_157),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_55),
.A2(n_59),
.B1(n_189),
.B2(n_248),
.Y(n_247)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_59),
.A2(n_67),
.B(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_59),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_64),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_85),
.B(n_86),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_76),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_85),
.B1(n_86),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_77),
.A2(n_82),
.B1(n_85),
.B2(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_78),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_78),
.A2(n_147),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_78),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_78),
.A2(n_172),
.B1(n_203),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_78),
.A2(n_125),
.B(n_205),
.Y(n_236)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_124),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_81),
.A2(n_149),
.B(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_90),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_107),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_105),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_101),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_137),
.B(n_314),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_136),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_112),
.B(n_136),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_113),
.B(n_117),
.Y(n_312)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_118),
.A2(n_119),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.C(n_134),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_120),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_121),
.B(n_127),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_126),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_200)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_136),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_308),
.B(n_313),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_296),
.B(n_307),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_193),
.B(n_275),
.C(n_295),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_182),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_141),
.B(n_182),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_165),
.B2(n_181),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_152),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_144),
.B(n_152),
.C(n_181),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_145),
.B(n_151),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_160),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_162),
.B(n_172),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_166),
.B(n_174),
.C(n_179),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_183),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_187),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_188),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_190),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_274),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_268),
.B(n_273),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_256),
.B(n_267),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_238),
.B(n_255),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_226),
.B(n_237),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_214),
.B(n_225),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_206),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_219),
.B(n_224),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_240),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_246),
.B1(n_253),
.B2(n_254),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_258),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_277),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_293),
.B2(n_294),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_283),
.C(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_292),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_290),
.C(n_292),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_298),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_304),
.C(n_306),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);


endmodule