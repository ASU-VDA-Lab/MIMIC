module fake_ariane_1256_n_1417 (n_295, n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_289, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_294, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_299, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_291, n_20, n_292, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_297, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_290, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_302, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_301, n_184, n_177, n_135, n_258, n_73, n_77, n_293, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_303, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_300, n_14, n_163, n_88, n_186, n_141, n_296, n_298, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1417);

input n_295;
input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_289;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_294;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_299;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_291;
input n_20;
input n_292;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_297;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_290;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_302;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_301;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_293;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_303;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_300;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_296;
input n_298;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1417;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_383;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_99),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_21),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_23),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_146),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_75),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_84),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_17),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_59),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_118),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_74),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_88),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_152),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_248),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_217),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_134),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_62),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_58),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_69),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_160),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_176),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_231),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_208),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_233),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_18),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_220),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_43),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_199),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_162),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_27),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_81),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_89),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_105),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_198),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_239),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_7),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_25),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_255),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_91),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_295),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_151),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_237),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_243),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_100),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_202),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_7),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_213),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_109),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_226),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_256),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_83),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_14),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_194),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_124),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_56),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_144),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_79),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_283),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_30),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_212),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_4),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_171),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_190),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_204),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_155),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_94),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_258),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_113),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_97),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_48),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_264),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_294),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_296),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_127),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_200),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_282),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_254),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_286),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_238),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_224),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_279),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_261),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_47),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_266),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_299),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_78),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_19),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_242),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_227),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_253),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_247),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_276),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_17),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_236),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_18),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_230),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_77),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_125),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_175),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_271),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_138),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_85),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_133),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_27),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_82),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_22),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_222),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_240),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_29),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_107),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_76),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_285),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_158),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_25),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_263),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_137),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_189),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_104),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_267),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_9),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_117),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_301),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_132),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_281),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_183),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_44),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_139),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_96),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_98),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_182),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_114),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_93),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_31),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_303),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_46),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_61),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_9),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_111),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_169),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_136),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_165),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_140),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_177),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_149),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_270),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_28),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_249),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_287),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_298),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_47),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_277),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_120),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_252),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_259),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_72),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_37),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_173),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_278),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_2),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_167),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_43),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_153),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_221),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_49),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_150),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_244),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_101),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_215),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_26),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_207),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_157),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_95),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_51),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g488 ( 
.A(n_290),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_250),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_161),
.Y(n_490)
);

BUFx10_ASAP7_75t_L g491 ( 
.A(n_156),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_24),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_184),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_195),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_4),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_33),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_49),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_143),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_35),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_147),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_193),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_268),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_209),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_232),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_8),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_273),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_280),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_274),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_192),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_178),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_284),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_80),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_6),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_219),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_70),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_73),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_225),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_71),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_128),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_112),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_289),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_126),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_141),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_64),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_6),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_170),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_241),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_154),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_55),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_447),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_344),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_418),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_373),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_306),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_354),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_397),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_347),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_513),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_305),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_344),
.Y(n_541)
);

INVxp33_ASAP7_75t_SL g542 ( 
.A(n_335),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_373),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_346),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_350),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_358),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_373),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_352),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_407),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_423),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_353),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_373),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_460),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_433),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_445),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_463),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_468),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_311),
.B(n_0),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_498),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_497),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_501),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g564 ( 
.A(n_337),
.B(n_0),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_318),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_311),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_340),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_332),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_332),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_420),
.Y(n_570)
);

INVxp33_ASAP7_75t_SL g571 ( 
.A(n_348),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_307),
.B(n_1),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_364),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_367),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_371),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_384),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_432),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_401),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_409),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_428),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_309),
.B(n_1),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_434),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_462),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_462),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_440),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_385),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_491),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_491),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_451),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_470),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_475),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_509),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_478),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_310),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_385),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_483),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_313),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_315),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_487),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_2),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_495),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_316),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_394),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_322),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_323),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_499),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_324),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_505),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_394),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_525),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_529),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_398),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_304),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_410),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_308),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_398),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_317),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_408),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_408),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_484),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_484),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_515),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_319),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_320),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_515),
.Y(n_632)
);

INVxp33_ASAP7_75t_SL g633 ( 
.A(n_314),
.Y(n_633)
);

INVxp33_ASAP7_75t_L g634 ( 
.A(n_321),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_327),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_325),
.Y(n_636)
);

CKINVDCx14_ASAP7_75t_R g637 ( 
.A(n_329),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_330),
.B(n_3),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_339),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_328),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_333),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_334),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_343),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_357),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_361),
.Y(n_645)
);

INVxp33_ASAP7_75t_SL g646 ( 
.A(n_336),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_338),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_342),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_376),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_378),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_345),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_349),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_410),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_387),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_389),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_326),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_351),
.Y(n_657)
);

CKINVDCx16_ASAP7_75t_R g658 ( 
.A(n_328),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_355),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_359),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_328),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_360),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_390),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_392),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_363),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_366),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_396),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_368),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_465),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_369),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_399),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_406),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_370),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_374),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_422),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_375),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_425),
.B(n_3),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_377),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_427),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_430),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_379),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_380),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_435),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_439),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_534),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_543),
.Y(n_686)
);

INVx6_ASAP7_75t_L g687 ( 
.A(n_640),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_532),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_600),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_312),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_583),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_535),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_621),
.B(n_490),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_602),
.B(n_443),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_537),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_656),
.B(n_341),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_538),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_532),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_550),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_584),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_559),
.B(n_328),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_553),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_557),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_634),
.B(n_412),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_586),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_592),
.B(n_365),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_602),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_628),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_593),
.B(n_372),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_541),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_331),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_530),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_601),
.B(n_446),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_566),
.B(n_474),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_531),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_634),
.B(n_480),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_600),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_672),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_604),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_672),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_658),
.B(n_356),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_565),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_570),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_609),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_611),
.B(n_467),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_572),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_612),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_661),
.B(n_362),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_614),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_636),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_633),
.B(n_414),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_545),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_639),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_643),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_645),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_653),
.B(n_417),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_638),
.B(n_431),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_649),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_622),
.B(n_438),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_548),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_650),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_654),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_SL g757 ( 
.A(n_619),
.B(n_482),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_655),
.B(n_331),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_544),
.B(n_521),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

OA21x2_ASAP7_75t_L g761 ( 
.A1(n_667),
.A2(n_502),
.B(n_494),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_539),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_671),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_581),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_675),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_679),
.Y(n_766)
);

AND2x2_ASAP7_75t_SL g767 ( 
.A(n_607),
.B(n_444),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_680),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_683),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_616),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_629),
.B(n_503),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_664),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_594),
.B(n_381),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_596),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_624),
.B(n_455),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_603),
.A2(n_507),
.B1(n_523),
.B2(n_518),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_599),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_646),
.B(n_508),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_669),
.B(n_527),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_549),
.B(n_500),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_585),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_630),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_SL g784 ( 
.A(n_619),
.B(n_331),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_677),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_631),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_641),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_647),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_610),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_714),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_688),
.B(n_623),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_701),
.B(n_564),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_SL g793 ( 
.A(n_787),
.B(n_635),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_710),
.B(n_637),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_693),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_693),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_761),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_727),
.B(n_637),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_767),
.A2(n_623),
.B1(n_626),
.B2(n_625),
.Y(n_799)
);

AND2x6_ASAP7_75t_SL g800 ( 
.A(n_779),
.B(n_603),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_765),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_721),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_786),
.B(n_542),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_765),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_779),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_746),
.B(n_551),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_740),
.B(n_651),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_740),
.B(n_657),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_720),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_787),
.B(n_659),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_728),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_740),
.B(n_662),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_754),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_761),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_693),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_714),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_736),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_700),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_765),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_766),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_770),
.B(n_571),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_687),
.B(n_725),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_723),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_736),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_766),
.Y(n_826)
);

BUFx10_ASAP7_75t_L g827 ( 
.A(n_787),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_687),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_723),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_759),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_766),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_694),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_736),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_685),
.B(n_582),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_688),
.B(n_665),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_700),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_696),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_704),
.B(n_627),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_689),
.B(n_555),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_785),
.A2(n_632),
.B1(n_618),
.B2(n_615),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_713),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_715),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_686),
.B(n_666),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_696),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_783),
.B(n_331),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_704),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_719),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_719),
.B(n_668),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_717),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_690),
.B(n_695),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_711),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_782),
.B(n_673),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_728),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_762),
.Y(n_855)
);

BUFx4f_ASAP7_75t_L g856 ( 
.A(n_783),
.Y(n_856)
);

INVx5_ASAP7_75t_L g857 ( 
.A(n_720),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_729),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_697),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_772),
.B(n_556),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_696),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_729),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_691),
.B(n_670),
.Y(n_864)
);

AND3x1_ASAP7_75t_L g865 ( 
.A(n_777),
.B(n_536),
.C(n_678),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_782),
.B(n_674),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_782),
.B(n_676),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_702),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_703),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_788),
.B(n_681),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_698),
.B(n_682),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_706),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_698),
.B(n_567),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_705),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_708),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_764),
.B(n_573),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_692),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_699),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_706),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_699),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_730),
.Y(n_881)
);

OR2x2_ASAP7_75t_SL g882 ( 
.A(n_762),
.B(n_536),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_725),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_734),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_735),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_881),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_881),
.Y(n_887)
);

AO22x2_ASAP7_75t_L g888 ( 
.A1(n_865),
.A2(n_789),
.B1(n_777),
.B2(n_742),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_811),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_878),
.B(n_880),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_878),
.B(n_733),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_842),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_843),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_854),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_840),
.B(n_724),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_884),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_850),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_850),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_802),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_859),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_828),
.B(n_554),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_868),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_869),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_874),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_875),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_828),
.B(n_558),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_885),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_L g908 ( 
.A(n_883),
.B(n_575),
.C(n_574),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_823),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_829),
.B(n_732),
.Y(n_910)
);

AO22x2_ASAP7_75t_L g911 ( 
.A1(n_864),
.A2(n_742),
.B1(n_745),
.B2(n_691),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_829),
.B(n_732),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_833),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_833),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_852),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_871),
.B(n_771),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_821),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_826),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_863),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_863),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_814),
.Y(n_922)
);

OAI221xp5_ASAP7_75t_L g923 ( 
.A1(n_873),
.A2(n_780),
.B1(n_771),
.B2(n_745),
.C(n_750),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_832),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_801),
.Y(n_925)
);

BUFx8_ASAP7_75t_L g926 ( 
.A(n_837),
.Y(n_926)
);

AO22x2_ASAP7_75t_L g927 ( 
.A1(n_864),
.A2(n_712),
.B1(n_718),
.B2(n_753),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_847),
.B(n_848),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_801),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_847),
.B(n_726),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_855),
.B(n_773),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_804),
.Y(n_932)
);

AO22x2_ASAP7_75t_L g933 ( 
.A1(n_831),
.A2(n_712),
.B1(n_718),
.B2(n_753),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_839),
.B(n_560),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_791),
.B(n_709),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_827),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_791),
.B(n_562),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_848),
.B(n_707),
.Y(n_938)
);

OAI221xp5_ASAP7_75t_L g939 ( 
.A1(n_794),
.A2(n_780),
.B1(n_750),
.B2(n_776),
.C(n_739),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_806),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_856),
.B(n_774),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_804),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_860),
.Y(n_943)
);

BUFx8_ASAP7_75t_L g944 ( 
.A(n_793),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_820),
.Y(n_945)
);

OAI221xp5_ASAP7_75t_L g946 ( 
.A1(n_798),
.A2(n_776),
.B1(n_739),
.B2(n_722),
.C(n_716),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_820),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_797),
.A2(n_757),
.B1(n_707),
.B2(n_751),
.Y(n_948)
);

AND2x6_ASAP7_75t_L g949 ( 
.A(n_797),
.B(n_775),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_799),
.A2(n_751),
.B1(n_533),
.B2(n_781),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_851),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_841),
.B(n_724),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_818),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_825),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_840),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_SL g956 ( 
.A(n_877),
.B(n_642),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_856),
.B(n_648),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_853),
.B(n_707),
.Y(n_958)
);

OR2x6_ASAP7_75t_SL g959 ( 
.A(n_866),
.B(n_576),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_819),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_834),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_838),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_845),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_822),
.A2(n_835),
.B1(n_844),
.B2(n_803),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_867),
.B(n_587),
.C(n_580),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_805),
.B(n_807),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_861),
.Y(n_967)
);

OAI221xp5_ASAP7_75t_L g968 ( 
.A1(n_792),
.A2(n_722),
.B1(n_731),
.B2(n_741),
.C(n_738),
.Y(n_968)
);

OAI221xp5_ASAP7_75t_L g969 ( 
.A1(n_808),
.A2(n_756),
.B1(n_763),
.B2(n_748),
.C(n_744),
.Y(n_969)
);

OAI221xp5_ASAP7_75t_L g970 ( 
.A1(n_812),
.A2(n_769),
.B1(n_768),
.B2(n_743),
.C(n_747),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_876),
.A2(n_810),
.B1(n_870),
.B2(n_660),
.Y(n_971)
);

AO22x2_ASAP7_75t_L g972 ( 
.A1(n_800),
.A2(n_533),
.B1(n_882),
.B2(n_781),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_836),
.A2(n_652),
.B1(n_784),
.B2(n_707),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_858),
.B(n_724),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_849),
.A2(n_769),
.B1(n_768),
.B2(n_590),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_805),
.B(n_595),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_862),
.B(n_737),
.Y(n_977)
);

AO22x2_ASAP7_75t_L g978 ( 
.A1(n_815),
.A2(n_568),
.B1(n_577),
.B2(n_569),
.Y(n_978)
);

AO22x2_ASAP7_75t_L g979 ( 
.A1(n_815),
.A2(n_589),
.B1(n_579),
.B2(n_749),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_790),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_830),
.B(n_597),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_916),
.B(n_830),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_964),
.B(n_790),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_931),
.B(n_598),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_951),
.B(n_813),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_966),
.B(n_890),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_973),
.B(n_813),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_940),
.B(n_813),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_936),
.B(n_817),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_976),
.B(n_817),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_922),
.B(n_824),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_975),
.B(n_824),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_891),
.B(n_606),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_974),
.B(n_608),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_960),
.B(n_943),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_617),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_908),
.B(n_956),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_971),
.B(n_752),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_981),
.B(n_755),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_965),
.B(n_760),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_909),
.B(n_778),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_889),
.B(n_778),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_894),
.B(n_872),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_901),
.B(n_809),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_930),
.B(n_941),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_887),
.B(n_846),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_899),
.B(n_846),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_935),
.B(n_879),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_958),
.B(n_809),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_937),
.B(n_809),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_906),
.B(n_795),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_SL g1012 ( 
.A(n_957),
.B(n_796),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_910),
.B(n_857),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_912),
.B(n_816),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_900),
.B(n_382),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_934),
.B(n_386),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_902),
.B(n_388),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_920),
.B(n_519),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_903),
.B(n_391),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_904),
.B(n_393),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_905),
.B(n_846),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_952),
.B(n_400),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_923),
.B(n_720),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_938),
.B(n_928),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_926),
.B(n_403),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_917),
.B(n_980),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_SL g1027 ( 
.A(n_925),
.B(n_404),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_892),
.B(n_405),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_893),
.B(n_411),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_897),
.B(n_413),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_898),
.B(n_415),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_913),
.B(n_416),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_915),
.B(n_720),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_914),
.B(n_419),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_948),
.B(n_421),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_SL g1036 ( 
.A(n_929),
.B(n_424),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_SL g1037 ( 
.A(n_932),
.B(n_426),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_921),
.B(n_528),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_939),
.B(n_758),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_946),
.B(n_758),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_942),
.B(n_429),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_945),
.B(n_947),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_955),
.B(n_436),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_955),
.B(n_437),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_SL g1045 ( 
.A(n_918),
.B(n_441),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_933),
.B(n_758),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_977),
.B(n_442),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_919),
.B(n_448),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_924),
.B(n_450),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_933),
.B(n_911),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_907),
.B(n_452),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_896),
.B(n_453),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_895),
.B(n_5),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_953),
.B(n_454),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_927),
.B(n_5),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_954),
.B(n_488),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_SL g1057 ( 
.A(n_984),
.B(n_944),
.Y(n_1057)
);

NAND4xp25_ASAP7_75t_SL g1058 ( 
.A(n_1055),
.B(n_968),
.C(n_969),
.D(n_888),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_SL g1059 ( 
.A1(n_982),
.A2(n_962),
.B(n_961),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_995),
.B(n_888),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_1011),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_986),
.B(n_911),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_993),
.A2(n_970),
.B(n_967),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1056),
.A2(n_963),
.B(n_949),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_997),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1004),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_1050),
.A2(n_949),
.A3(n_927),
.B(n_950),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_1046),
.A2(n_949),
.A3(n_950),
.B(n_979),
.Y(n_1068)
);

NAND2x1_ASAP7_75t_L g1069 ( 
.A(n_1006),
.B(n_758),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_1039),
.A2(n_979),
.A3(n_959),
.B(n_972),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_996),
.A2(n_978),
.B(n_972),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_SL g1072 ( 
.A1(n_1040),
.A2(n_1023),
.B(n_1021),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_994),
.B(n_978),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_983),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_1053),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_SL g1076 ( 
.A(n_1005),
.B(n_383),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1009),
.A2(n_488),
.B(n_63),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1026),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1022),
.B(n_456),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1024),
.A2(n_458),
.B(n_457),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_998),
.B(n_10),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_991),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_SL g1083 ( 
.A1(n_985),
.A2(n_488),
.B(n_395),
.C(n_402),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_988),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1007),
.A2(n_488),
.A3(n_395),
.B(n_402),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1018),
.A2(n_488),
.B(n_65),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_1015),
.B(n_459),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1008),
.B(n_11),
.Y(n_1088)
);

BUFx8_ASAP7_75t_L g1089 ( 
.A(n_1025),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1001),
.B(n_461),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1002),
.B(n_11),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_999),
.B(n_466),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_1012),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1003),
.B(n_12),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1018),
.A2(n_66),
.B(n_60),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1010),
.B(n_12),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_987),
.A2(n_395),
.B(n_383),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1038),
.A2(n_68),
.B(n_67),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1038),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1016),
.B(n_469),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1045),
.B(n_526),
.Y(n_1101)
);

AO32x2_ASAP7_75t_L g1102 ( 
.A1(n_992),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1033),
.A2(n_1014),
.B(n_1035),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_1042),
.A2(n_383),
.A3(n_476),
.B(n_402),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1000),
.A2(n_472),
.B(n_471),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1028),
.A2(n_479),
.B(n_477),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_990),
.A2(n_383),
.A3(n_476),
.B(n_402),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1043),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1029),
.A2(n_524),
.B1(n_522),
.B2(n_520),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_989),
.B(n_19),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1030),
.A2(n_485),
.B(n_481),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1027),
.A2(n_517),
.B1(n_516),
.B2(n_514),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1036),
.A2(n_512),
.B(n_511),
.C(n_510),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1041),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1017),
.B(n_20),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1054),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1031),
.A2(n_489),
.B(n_486),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1072),
.A2(n_1013),
.B(n_1047),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_1064),
.A2(n_1034),
.B(n_1032),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_1059),
.A2(n_1049),
.B(n_1048),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1078),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_1057),
.B(n_476),
.Y(n_1122)
);

BUFx5_ASAP7_75t_L g1123 ( 
.A(n_1074),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1062),
.B(n_1060),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1077),
.A2(n_1051),
.B(n_1020),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1089),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_1097),
.A2(n_1063),
.B(n_1076),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_1103),
.A2(n_1019),
.B(n_1044),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1066),
.B(n_86),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1099),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_1086),
.A2(n_1037),
.B(n_1052),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1061),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1067),
.B(n_21),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1081),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1083),
.A2(n_90),
.B(n_87),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1069),
.A2(n_476),
.B(n_493),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1083),
.A2(n_1098),
.B(n_1095),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1066),
.B(n_92),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1058),
.B(n_504),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1065),
.B(n_22),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_1093),
.B(n_23),
.Y(n_1141)
);

AO21x2_ASAP7_75t_L g1142 ( 
.A1(n_1088),
.A2(n_1080),
.B(n_1115),
.Y(n_1142)
);

CKINVDCx6p67_ASAP7_75t_R g1143 ( 
.A(n_1075),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1067),
.B(n_24),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1071),
.A2(n_1073),
.B1(n_1091),
.B2(n_1116),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1099),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1094),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1105),
.A2(n_506),
.B(n_26),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1079),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1070),
.B(n_32),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1096),
.A2(n_103),
.B(n_102),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1113),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1108),
.B(n_32),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1104),
.A2(n_188),
.B(n_297),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1087),
.A2(n_187),
.B(n_293),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1101),
.A2(n_186),
.B(n_292),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1082),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1102),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1090),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1102),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1085),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1085),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1093),
.Y(n_1163)
);

AO21x2_ASAP7_75t_L g1164 ( 
.A1(n_1106),
.A2(n_191),
.B(n_291),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1070),
.B(n_36),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1082),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1068),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1100),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1109),
.A2(n_1092),
.B1(n_1112),
.B2(n_1084),
.C(n_1111),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1084),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1068),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1107),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1107),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1167),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1123),
.Y(n_1175)
);

CKINVDCx11_ASAP7_75t_R g1176 ( 
.A(n_1126),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1171),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1137),
.A2(n_1117),
.B(n_197),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1139),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1158),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1132),
.B(n_41),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1160),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1123),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1139),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1172),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1134),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1161),
.A2(n_45),
.B(n_46),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1123),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1161),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1131),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1166),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1123),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1162),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1123),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1123),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1121),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1163),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1129),
.B(n_106),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1149),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1133),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1162),
.A2(n_50),
.B(n_53),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1135),
.A2(n_201),
.B(n_288),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1173),
.Y(n_1203)
);

INVx6_ASAP7_75t_SL g1204 ( 
.A(n_1129),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1124),
.B(n_53),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1144),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1144),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1163),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1154),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1154),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1147),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1119),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1119),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1138),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1130),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1128),
.Y(n_1216)
);

AOI222xp33_ASAP7_75t_L g1217 ( 
.A1(n_1140),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.C1(n_57),
.C2(n_108),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1128),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1127),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1149),
.A2(n_57),
.B(n_110),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1148),
.A2(n_115),
.B(n_116),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1150),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1118),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1165),
.B(n_119),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1140),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1138),
.B(n_129),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1131),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_L g1228 ( 
.A(n_1163),
.B(n_130),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1214),
.B(n_1141),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1186),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_R g1231 ( 
.A(n_1198),
.B(n_1141),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_R g1232 ( 
.A(n_1176),
.B(n_1143),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_R g1233 ( 
.A(n_1198),
.B(n_1141),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1211),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1226),
.B(n_1130),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_1197),
.B(n_1122),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1197),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1208),
.B(n_1170),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1208),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1205),
.B(n_1153),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1205),
.B(n_1157),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_R g1242 ( 
.A(n_1187),
.B(n_1146),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_R g1243 ( 
.A(n_1228),
.B(n_1122),
.Y(n_1243)
);

XNOR2xp5_ASAP7_75t_L g1244 ( 
.A(n_1225),
.B(n_1145),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1181),
.B(n_1152),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1200),
.B(n_1130),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1215),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_R g1248 ( 
.A(n_1187),
.B(n_1155),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1191),
.B(n_1142),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1196),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_R g1251 ( 
.A(n_1201),
.B(n_1156),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1224),
.B(n_1159),
.Y(n_1252)
);

NAND2xp33_ASAP7_75t_SL g1253 ( 
.A(n_1204),
.B(n_1120),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1179),
.B(n_1169),
.Y(n_1254)
);

BUFx5_ASAP7_75t_L g1255 ( 
.A(n_1223),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_R g1256 ( 
.A(n_1201),
.B(n_1151),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1206),
.B(n_1168),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1174),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1207),
.B(n_1169),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1222),
.B(n_1125),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1177),
.B(n_1164),
.Y(n_1261)
);

XNOR2xp5_ASAP7_75t_L g1262 ( 
.A(n_1199),
.B(n_1184),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1204),
.B(n_1148),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1203),
.B(n_1164),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1174),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1185),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_1189),
.B(n_131),
.Y(n_1267)
);

CKINVDCx14_ASAP7_75t_R g1268 ( 
.A(n_1180),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1180),
.B(n_1136),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1182),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1230),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1268),
.B(n_1182),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1270),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1250),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1244),
.A2(n_1220),
.B1(n_1217),
.B2(n_1183),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1234),
.B(n_1189),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1245),
.B(n_1175),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1237),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1258),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1229),
.B(n_1188),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1247),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1240),
.B(n_1193),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1265),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1266),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1246),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1249),
.B(n_1216),
.Y(n_1287)
);

BUFx5_ASAP7_75t_L g1288 ( 
.A(n_1264),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1229),
.B(n_1192),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1235),
.B(n_1192),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1257),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1238),
.B(n_1218),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1254),
.A2(n_1194),
.B1(n_1195),
.B2(n_1223),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1269),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1262),
.A2(n_1195),
.B1(n_1210),
.B2(n_1213),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1260),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1241),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1242),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1261),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1235),
.B(n_1190),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1239),
.B(n_1190),
.Y(n_1301)
);

OR2x2_ASAP7_75t_SL g1302 ( 
.A(n_1231),
.B(n_1212),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1255),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1252),
.B(n_1263),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1283),
.B(n_1271),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1291),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1277),
.B(n_1255),
.Y(n_1307)
);

NOR2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1304),
.B(n_1233),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1271),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1272),
.B(n_1255),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1303),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1282),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1296),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1273),
.Y(n_1314)
);

AND2x2_ASAP7_75t_SL g1315 ( 
.A(n_1298),
.B(n_1267),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1276),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1282),
.Y(n_1317)
);

AOI33xp33_ASAP7_75t_L g1318 ( 
.A1(n_1284),
.A2(n_1210),
.A3(n_1212),
.B1(n_1256),
.B2(n_1248),
.B3(n_1251),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1294),
.B(n_1227),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1280),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1286),
.B(n_1227),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1276),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1275),
.A2(n_1221),
.B1(n_1243),
.B2(n_1253),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1285),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1295),
.A2(n_1209),
.B(n_1219),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1299),
.B(n_1219),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1279),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1301),
.B(n_1178),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1306),
.B(n_1290),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1316),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1306),
.B(n_1297),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1312),
.B(n_1300),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1312),
.B(n_1292),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1314),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1314),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1309),
.B(n_1317),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1320),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1310),
.B(n_1274),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1320),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1322),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1319),
.B(n_1281),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1322),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1324),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1307),
.B(n_1289),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1305),
.Y(n_1345)
);

INVxp33_ASAP7_75t_L g1346 ( 
.A(n_1329),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1330),
.B(n_1321),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1331),
.B(n_1318),
.Y(n_1348)
);

AO221x2_ASAP7_75t_L g1349 ( 
.A1(n_1334),
.A2(n_1275),
.B1(n_1327),
.B2(n_1295),
.C(n_1315),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1336),
.Y(n_1350)
);

INVxp33_ASAP7_75t_SL g1351 ( 
.A(n_1329),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1345),
.A2(n_1315),
.B1(n_1323),
.B2(n_1308),
.Y(n_1352)
);

CKINVDCx8_ASAP7_75t_R g1353 ( 
.A(n_1333),
.Y(n_1353)
);

NOR2x1_ASAP7_75t_L g1354 ( 
.A(n_1333),
.B(n_1327),
.Y(n_1354)
);

AO221x2_ASAP7_75t_L g1355 ( 
.A1(n_1335),
.A2(n_1232),
.B1(n_1293),
.B2(n_1302),
.C(n_1278),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_L g1356 ( 
.A(n_1333),
.B(n_1311),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1337),
.Y(n_1357)
);

CKINVDCx8_ASAP7_75t_R g1358 ( 
.A(n_1341),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1348),
.B(n_1340),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1357),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1354),
.B(n_1332),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1350),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1358),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1347),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1351),
.B(n_1343),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1346),
.B(n_1342),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1349),
.B(n_1339),
.Y(n_1367)
);

NAND3xp33_ASAP7_75t_L g1368 ( 
.A(n_1355),
.B(n_1311),
.C(n_1293),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1356),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1352),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1353),
.B(n_1332),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1363),
.B(n_1355),
.Y(n_1372)
);

AOI211xp5_ASAP7_75t_L g1373 ( 
.A1(n_1367),
.A2(n_1368),
.B(n_1359),
.C(n_1370),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1363),
.A2(n_1341),
.B(n_1338),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1360),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1363),
.B(n_1371),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1360),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1375),
.B(n_1364),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1376),
.B(n_1371),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1372),
.B(n_1361),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1377),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1373),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1379),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1378),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1380),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1383),
.B(n_1365),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1382),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1380),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1380),
.Y(n_1390)
);

NOR4xp25_ASAP7_75t_L g1391 ( 
.A(n_1387),
.B(n_1381),
.C(n_1362),
.D(n_1365),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1385),
.A2(n_1369),
.B(n_1366),
.C(n_1325),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1384),
.B(n_1366),
.Y(n_1393)
);

NOR3x1_ASAP7_75t_L g1394 ( 
.A(n_1389),
.B(n_1178),
.C(n_1287),
.Y(n_1394)
);

NOR4xp75_ASAP7_75t_L g1395 ( 
.A(n_1386),
.B(n_1313),
.C(n_1328),
.D(n_1344),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1388),
.Y(n_1396)
);

NOR2x1_ASAP7_75t_SL g1397 ( 
.A(n_1390),
.B(n_1325),
.Y(n_1397)
);

AOI322xp5_ASAP7_75t_L g1398 ( 
.A1(n_1393),
.A2(n_1396),
.A3(n_1391),
.B1(n_1392),
.B2(n_1394),
.C1(n_1395),
.C2(n_1397),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1393),
.B(n_1326),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1399),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_SL g1401 ( 
.A(n_1398),
.B(n_1236),
.C(n_1202),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1399),
.B(n_135),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1400),
.B(n_1401),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1402),
.B(n_142),
.C(n_145),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1401),
.B(n_1288),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1403),
.A2(n_1288),
.B1(n_1185),
.B2(n_148),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1404),
.B(n_302),
.C(n_163),
.Y(n_1407)
);

OAI211xp5_ASAP7_75t_L g1408 ( 
.A1(n_1406),
.A2(n_1405),
.B(n_166),
.C(n_168),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1407),
.A2(n_172),
.B1(n_174),
.B2(n_179),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1408),
.B(n_180),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1409),
.A2(n_181),
.B(n_196),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1410),
.A2(n_206),
.B1(n_210),
.B2(n_214),
.Y(n_1412)
);

OAI322xp33_ASAP7_75t_L g1413 ( 
.A1(n_1412),
.A2(n_1411),
.A3(n_223),
.B1(n_228),
.B2(n_229),
.C1(n_234),
.C2(n_235),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1413),
.A2(n_245),
.B(n_246),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1414),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1415),
.A2(n_251),
.B1(n_260),
.B2(n_262),
.C(n_265),
.Y(n_1416)
);

AOI211xp5_ASAP7_75t_L g1417 ( 
.A1(n_1416),
.A2(n_269),
.B(n_272),
.C(n_275),
.Y(n_1417)
);


endmodule