module fake_netlist_1_5739_n_41 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_25;
wire n_26;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g16 ( .A(n_11), .B(n_13), .Y(n_16) );
OR2x6_ASAP7_75t_L g17 ( .A(n_2), .B(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_4), .B(n_7), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_12), .B(n_6), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_5), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_0), .A2(n_3), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_21), .B(n_1), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_21), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_24), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_27), .B(n_23), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_17), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_29), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_17), .B1(n_25), .B2(n_19), .Y(n_33) );
OAI21xp33_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_22), .B(n_17), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_22), .B(n_19), .Y(n_35) );
NOR2x1_ASAP7_75t_L g36 ( .A(n_35), .B(n_17), .Y(n_36) );
NAND4xp75_ASAP7_75t_L g37 ( .A(n_34), .B(n_20), .C(n_16), .D(n_4), .Y(n_37) );
OAI21xp5_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_21), .B(n_20), .Y(n_38) );
OAI21x1_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_8), .B(n_9), .Y(n_39) );
OAI21xp5_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_1), .B(n_2), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .B1(n_10), .B2(n_14), .Y(n_41) );
endmodule