module fake_netlist_5_2290_n_1075 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1075);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1075;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_568;
wire n_509;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_696;
wire n_255;
wire n_522;
wire n_897;
wire n_798;
wire n_350;
wire n_1020;
wire n_662;
wire n_459;
wire n_646;
wire n_1062;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_685;
wire n_598;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_969;
wire n_1069;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1028;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_632;
wire n_489;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_647;
wire n_679;
wire n_425;
wire n_513;
wire n_710;
wire n_407;
wire n_527;
wire n_707;
wire n_480;
wire n_832;
wire n_795;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

BUFx2_ASAP7_75t_R g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_174),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_94),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_22),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_201),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_211),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_48),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_123),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_107),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_71),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_85),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_140),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_138),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_164),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_154),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_180),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_67),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_98),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_173),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_181),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_30),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_89),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_244),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_90),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_205),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_99),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_159),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_86),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_163),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_17),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_104),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_183),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_184),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_88),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_142),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_147),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_130),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_242),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_84),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_56),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_102),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_218),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_122),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_76),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_0),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_252),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_304),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_50),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_51),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_307),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_0),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_249),
.B(n_1),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_1),
.Y(n_333)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_52),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

BUFx8_ASAP7_75t_SL g337 ( 
.A(n_264),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

BUFx8_ASAP7_75t_SL g339 ( 
.A(n_264),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_2),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_2),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_254),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_256),
.B(n_3),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_3),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_270),
.B(n_53),
.Y(n_349)
);

BUFx12f_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_246),
.B(n_4),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_272),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_274),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_251),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_345),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_300),
.B1(n_285),
.B2(n_287),
.Y(n_356)
);

AO22x2_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_292),
.B1(n_299),
.B2(n_275),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_251),
.B1(n_310),
.B2(n_287),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_248),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_321),
.A2(n_300),
.B1(n_285),
.B2(n_255),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_253),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_257),
.Y(n_367)
);

NAND3x1_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_303),
.C(n_301),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g369 ( 
.A1(n_335),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_259),
.B1(n_260),
.B2(n_258),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_269),
.B1(n_273),
.B2(n_267),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_276),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_322),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_282),
.B1(n_283),
.B2(n_281),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_R g378 ( 
.A1(n_348),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_322),
.A2(n_324),
.B1(n_331),
.B2(n_326),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_284),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_286),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_288),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_327),
.A2(n_297),
.B1(n_298),
.B2(n_296),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_327),
.A2(n_308),
.B1(n_11),
.B2(n_9),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_338),
.A2(n_350),
.B1(n_346),
.B2(n_322),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_324),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g394 ( 
.A(n_324),
.B(n_13),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_338),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_L g396 ( 
.A1(n_350),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_314),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_349),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_399)
);

AO22x2_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_326),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g402 ( 
.A(n_332),
.B(n_24),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_54),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_332),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_332),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_337),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_397),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_394),
.B(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

NAND2x1p5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_399),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_355),
.B(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

BUFx6f_ASAP7_75t_SL g425 ( 
.A(n_359),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_332),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_317),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_382),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_386),
.B(n_339),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_373),
.B(n_339),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_317),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_372),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_371),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_387),
.B(n_336),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_341),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_377),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

XNOR2x2_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_330),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_341),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_401),
.B(n_333),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_374),
.Y(n_458)
);

OR2x2_ASAP7_75t_SL g459 ( 
.A(n_378),
.B(n_340),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_358),
.B(n_340),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_370),
.B(n_341),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_395),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_340),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_359),
.B(n_341),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_379),
.A2(n_341),
.B(n_313),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_356),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_340),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_440),
.B(n_312),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_25),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_412),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_334),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_447),
.A2(n_334),
.B(n_313),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_431),
.B(n_312),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_334),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_334),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_334),
.Y(n_491)
);

AND2x2_ASAP7_75t_SL g492 ( 
.A(n_417),
.B(n_319),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_319),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_447),
.B(n_319),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_410),
.B(n_456),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_409),
.B(n_319),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_453),
.B(n_441),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_320),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_460),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_411),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_445),
.B(n_411),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_320),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_466),
.A2(n_313),
.B(n_312),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_457),
.B(n_320),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_320),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_469),
.B(n_27),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_442),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_446),
.B(n_55),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_448),
.B(n_312),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_449),
.B(n_312),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_316),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_468),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_313),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_469),
.A2(n_316),
.B1(n_315),
.B2(n_313),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_450),
.B(n_315),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_455),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_465),
.B(n_454),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_455),
.B(n_315),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_458),
.B(n_58),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_462),
.B(n_59),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_420),
.B(n_315),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_315),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_465),
.B(n_316),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_463),
.B(n_316),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_316),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_468),
.B(n_60),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_407),
.B(n_61),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_444),
.B(n_62),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_432),
.A2(n_413),
.B(n_64),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_444),
.B(n_63),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_459),
.B(n_65),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_527),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_501),
.B(n_422),
.Y(n_547)
);

BUFx8_ASAP7_75t_SL g548 ( 
.A(n_539),
.Y(n_548)
);

BUFx6f_ASAP7_75t_SL g549 ( 
.A(n_540),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_501),
.B(n_433),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_497),
.B(n_435),
.Y(n_551)
);

INVx8_ASAP7_75t_L g552 ( 
.A(n_543),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_435),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_502),
.B(n_490),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_500),
.B(n_425),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_477),
.B(n_66),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_500),
.B(n_425),
.Y(n_557)
);

AND2x2_ASAP7_75t_SL g558 ( 
.A(n_530),
.B(n_27),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_68),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_477),
.B(n_504),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_514),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_69),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_514),
.B(n_28),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_543),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_483),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_505),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_497),
.B(n_70),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_477),
.B(n_72),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_530),
.B(n_29),
.Y(n_571)
);

BUFx4f_ASAP7_75t_L g572 ( 
.A(n_543),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_530),
.B(n_29),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_506),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_478),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_497),
.B(n_73),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_495),
.B(n_516),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_506),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_506),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_495),
.B(n_74),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_75),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_538),
.B(n_30),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_531),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_538),
.B(n_31),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_518),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_513),
.B(n_77),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_492),
.B(n_476),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_473),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_513),
.B(n_78),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_492),
.B(n_31),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_478),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_473),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_518),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_528),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_474),
.Y(n_603)
);

NAND2x1_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_79),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_564),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_554),
.B(n_527),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_564),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_546),
.Y(n_611)
);

INVx6_ASAP7_75t_L g612 ( 
.A(n_569),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_545),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx4_ASAP7_75t_SL g616 ( 
.A(n_559),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_553),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_548),
.Y(n_620)
);

INVx6_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_578),
.B(n_516),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_551),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_578),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

NAND2x1p5_ASAP7_75t_L g627 ( 
.A(n_586),
.B(n_478),
.Y(n_627)
);

BUFx2_ASAP7_75t_SL g628 ( 
.A(n_549),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_590),
.A2(n_492),
.B1(n_540),
.B2(n_543),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_583),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_567),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_546),
.Y(n_635)
);

BUFx2_ASAP7_75t_R g636 ( 
.A(n_596),
.Y(n_636)
);

NAND2x1p5_ASAP7_75t_L g637 ( 
.A(n_586),
.B(n_479),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_565),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_563),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_563),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_568),
.Y(n_642)
);

INVx3_ASAP7_75t_SL g643 ( 
.A(n_558),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_574),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_550),
.Y(n_645)
);

NAND2x1p5_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_588),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_576),
.Y(n_647)
);

INVx5_ASAP7_75t_SL g648 ( 
.A(n_583),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_555),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

INVx5_ASAP7_75t_SL g651 ( 
.A(n_579),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_579),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_559),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_555),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

BUFx4f_ASAP7_75t_SL g656 ( 
.A(n_601),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_595),
.Y(n_657)
);

BUFx6f_ASAP7_75t_SL g658 ( 
.A(n_601),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_549),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_601),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_575),
.Y(n_661)
);

BUFx12f_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_557),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_587),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_580),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_664),
.A2(n_571),
.B1(n_573),
.B2(n_587),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_609),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_608),
.B(n_602),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_656),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_660),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_664),
.A2(n_543),
.B1(n_539),
.B2(n_542),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_666),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_633),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_609),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_616),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_643),
.A2(n_571),
.B1(n_573),
.B2(n_585),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_666),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_640),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_642),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_658),
.Y(n_682)
);

INVx6_ASAP7_75t_L g683 ( 
.A(n_616),
.Y(n_683)
);

BUFx12f_ASAP7_75t_L g684 ( 
.A(n_659),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_644),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_620),
.Y(n_686)
);

BUFx4_ASAP7_75t_R g687 ( 
.A(n_607),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_661),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_649),
.A2(n_593),
.B1(n_542),
.B2(n_531),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_L g690 ( 
.A1(n_643),
.A2(n_593),
.B1(n_602),
.B2(n_586),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_650),
.A2(n_531),
.B1(n_517),
.B2(n_532),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_620),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

INVx6_ASAP7_75t_L g695 ( 
.A(n_616),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_629),
.A2(n_531),
.B1(n_517),
.B2(n_532),
.Y(n_696)
);

CKINVDCx11_ASAP7_75t_R g697 ( 
.A(n_624),
.Y(n_697)
);

BUFx8_ASAP7_75t_L g698 ( 
.A(n_658),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_645),
.A2(n_531),
.B1(n_517),
.B2(n_533),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_614),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_641),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_617),
.A2(n_531),
.B1(n_533),
.B2(n_595),
.Y(n_703)
);

BUFx8_ASAP7_75t_SL g704 ( 
.A(n_659),
.Y(n_704)
);

BUFx4f_ASAP7_75t_SL g705 ( 
.A(n_624),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_639),
.A2(n_531),
.B1(n_552),
.B2(n_498),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_614),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_639),
.A2(n_531),
.B1(n_552),
.B2(n_562),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_SL g709 ( 
.A1(n_649),
.A2(n_552),
.B1(n_566),
.B2(n_562),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_613),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_612),
.A2(n_621),
.B1(n_610),
.B2(n_607),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_632),
.A2(n_566),
.B1(n_572),
.B2(n_471),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_632),
.A2(n_572),
.B1(n_512),
.B2(n_570),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_628),
.Y(n_715)
);

CKINVDCx11_ASAP7_75t_R g716 ( 
.A(n_634),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_655),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_529),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_672),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_613),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_623),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_667),
.A2(n_634),
.B1(n_654),
.B2(n_638),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_675),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_678),
.B(n_657),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_680),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_673),
.A2(n_626),
.B1(n_631),
.B2(n_619),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_687),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_689),
.A2(n_696),
.B1(n_690),
.B2(n_638),
.Y(n_729)
);

BUFx8_ASAP7_75t_SL g730 ( 
.A(n_686),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_692),
.A2(n_615),
.B1(n_663),
.B2(n_541),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_702),
.B(n_648),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_681),
.A2(n_541),
.B1(n_481),
.B2(n_610),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

CKINVDCx11_ASAP7_75t_R g735 ( 
.A(n_693),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_711),
.B(n_648),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_705),
.A2(n_619),
.B1(n_631),
.B2(n_626),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_700),
.A2(n_648),
.B1(n_621),
.B2(n_612),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_687),
.B(n_622),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_712),
.A2(n_621),
.B1(n_612),
.B2(n_622),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_688),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_668),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_715),
.A2(n_626),
.B1(n_631),
.B2(n_619),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_703),
.A2(n_481),
.B1(n_625),
.B2(n_653),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_714),
.A2(n_625),
.B1(n_622),
.B2(n_619),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_674),
.B(n_652),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_674),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_677),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_SL g749 ( 
.A(n_682),
.B(n_636),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_697),
.A2(n_653),
.B1(n_489),
.B2(n_499),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_SL g751 ( 
.A1(n_706),
.A2(n_509),
.B(n_484),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_713),
.A2(n_662),
.B1(n_651),
.B2(n_652),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_697),
.A2(n_653),
.B1(n_489),
.B2(n_499),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_716),
.A2(n_486),
.B1(n_662),
.B2(n_591),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_709),
.A2(n_631),
.B1(n_626),
.B2(n_651),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_716),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_676),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_679),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_679),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_708),
.A2(n_651),
.B1(n_570),
.B2(n_556),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_SL g762 ( 
.A1(n_717),
.A2(n_484),
.B(n_556),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_693),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_670),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_698),
.A2(n_665),
.B1(n_528),
.B2(n_512),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_670),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_682),
.B(n_710),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_677),
.A2(n_600),
.B1(n_584),
.B2(n_592),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_691),
.Y(n_770)
);

OAI22x1_ASAP7_75t_SL g771 ( 
.A1(n_686),
.A2(n_507),
.B1(n_486),
.B2(n_515),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_694),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_682),
.A2(n_472),
.B1(n_485),
.B2(n_665),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_699),
.A2(n_599),
.B1(n_603),
.B2(n_582),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_677),
.A2(n_600),
.B1(n_584),
.B2(n_592),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_699),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_698),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_694),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_701),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_731),
.A2(n_475),
.B1(n_684),
.B2(n_507),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_720),
.B(n_701),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_SL g783 ( 
.A(n_733),
.B(n_494),
.C(n_535),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_723),
.A2(n_677),
.B1(n_695),
.B2(n_683),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_742),
.Y(n_785)
);

OAI222xp33_ASAP7_75t_L g786 ( 
.A1(n_723),
.A2(n_494),
.B1(n_707),
.B2(n_589),
.C1(n_606),
.C2(n_598),
.Y(n_786)
);

OAI221xp5_ASAP7_75t_L g787 ( 
.A1(n_731),
.A2(n_733),
.B1(n_765),
.B2(n_755),
.C(n_754),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_749),
.A2(n_684),
.B1(n_695),
.B2(n_683),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_758),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_728),
.A2(n_695),
.B1(n_683),
.B2(n_589),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_725),
.A2(n_475),
.B1(n_482),
.B2(n_508),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_728),
.A2(n_475),
.B1(n_482),
.B2(n_508),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_721),
.B(n_707),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_729),
.A2(n_508),
.B1(n_522),
.B2(n_515),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_729),
.A2(n_522),
.B1(n_695),
.B2(n_683),
.Y(n_796)
);

OAI221xp5_ASAP7_75t_SL g797 ( 
.A1(n_750),
.A2(n_754),
.B1(n_751),
.B2(n_755),
.C(n_744),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_744),
.A2(n_581),
.B1(n_491),
.B2(n_521),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_739),
.A2(n_510),
.B1(n_717),
.B2(n_521),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_524),
.C(n_491),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_753),
.A2(n_646),
.B1(n_637),
.B2(n_627),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_739),
.A2(n_510),
.B1(n_535),
.B2(n_710),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_727),
.A2(n_479),
.B1(n_493),
.B2(n_630),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_750),
.A2(n_646),
.B1(n_637),
.B2(n_627),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_780),
.B(n_710),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_740),
.A2(n_630),
.B1(n_536),
.B2(n_710),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_774),
.A2(n_536),
.B1(n_479),
.B2(n_655),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_SL g808 ( 
.A1(n_756),
.A2(n_588),
.B(n_611),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_736),
.A2(n_479),
.B1(n_525),
.B2(n_605),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_771),
.A2(n_493),
.B1(n_487),
.B2(n_480),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_726),
.B(n_710),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_745),
.A2(n_488),
.B1(n_537),
.B2(n_704),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_757),
.A2(n_537),
.B1(n_704),
.B2(n_503),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_761),
.A2(n_503),
.B1(n_605),
.B2(n_594),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_764),
.A2(n_525),
.B1(n_594),
.B2(n_635),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_778),
.A2(n_766),
.B1(n_776),
.B2(n_769),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_778),
.A2(n_503),
.B1(n_671),
.B2(n_534),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_767),
.A2(n_773),
.B1(n_779),
.B2(n_732),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_735),
.A2(n_503),
.B1(n_671),
.B2(n_534),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_730),
.A2(n_671),
.B1(n_611),
.B2(n_635),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_779),
.A2(n_611),
.B1(n_671),
.B2(n_660),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_763),
.A2(n_660),
.B1(n_529),
.B2(n_526),
.Y(n_822)
);

AO22x1_ASAP7_75t_L g823 ( 
.A1(n_724),
.A2(n_526),
.B1(n_520),
.B2(n_519),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_734),
.A2(n_480),
.B1(n_487),
.B2(n_496),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_737),
.A2(n_520),
.B1(n_519),
.B2(n_511),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_780),
.B(n_32),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_SL g827 ( 
.A1(n_741),
.A2(n_496),
.B1(n_33),
.B2(n_34),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_746),
.A2(n_523),
.B1(n_511),
.B2(n_518),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_775),
.A2(n_511),
.B1(n_523),
.B2(n_34),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_743),
.A2(n_523),
.B1(n_511),
.B2(n_35),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_SL g831 ( 
.A(n_748),
.B(n_32),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_748),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_768),
.A2(n_759),
.B1(n_770),
.B2(n_722),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_782),
.B(n_794),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_791),
.B(n_742),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_790),
.B(n_747),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_827),
.B(n_762),
.C(n_775),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_SL g838 ( 
.A1(n_810),
.A2(n_777),
.B1(n_772),
.B2(n_760),
.C(n_752),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_832),
.B(n_752),
.C(n_747),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_787),
.A2(n_768),
.B1(n_772),
.B2(n_777),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_SL g841 ( 
.A1(n_816),
.A2(n_760),
.B(n_36),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_SL g842 ( 
.A1(n_781),
.A2(n_830),
.B1(n_796),
.B2(n_813),
.C(n_800),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_799),
.B(n_80),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_831),
.B(n_37),
.C(n_38),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_811),
.B(n_37),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_805),
.B(n_38),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_805),
.B(n_39),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_818),
.B(n_39),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_789),
.B(n_40),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_SL g850 ( 
.A1(n_788),
.A2(n_40),
.B(n_41),
.Y(n_850)
);

AND4x1_ASAP7_75t_L g851 ( 
.A(n_820),
.B(n_41),
.C(n_42),
.D(n_43),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_789),
.B(n_42),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_826),
.B(n_44),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_826),
.B(n_44),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_785),
.B(n_833),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_831),
.B(n_45),
.C(n_46),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_785),
.B(n_45),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_795),
.B(n_46),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_792),
.B(n_47),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_802),
.B(n_47),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_812),
.B(n_48),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_797),
.B(n_822),
.C(n_819),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_823),
.B(n_49),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_823),
.B(n_49),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_786),
.B(n_81),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_806),
.B(n_82),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_83),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_783),
.A2(n_87),
.B(n_91),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_798),
.B(n_824),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_801),
.B(n_92),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_793),
.B(n_93),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_784),
.B(n_95),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_809),
.B(n_96),
.Y(n_873)
);

AOI221xp5_ASAP7_75t_L g874 ( 
.A1(n_829),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.C(n_103),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_817),
.B(n_105),
.C(n_106),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_803),
.B(n_807),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_815),
.B(n_821),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_828),
.B(n_108),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_825),
.B(n_109),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_110),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_SL g881 ( 
.A1(n_808),
.A2(n_111),
.B(n_112),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_808),
.B(n_113),
.C(n_114),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_790),
.B(n_115),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_782),
.B(n_116),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_117),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_L g886 ( 
.A(n_827),
.B(n_118),
.C(n_119),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_836),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_855),
.B(n_863),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_848),
.B(n_845),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_834),
.B(n_120),
.Y(n_890)
);

AO21x1_ASAP7_75t_SL g891 ( 
.A1(n_864),
.A2(n_121),
.B(n_124),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_855),
.B(n_125),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_851),
.B(n_126),
.C(n_127),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_863),
.B(n_128),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_843),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_843),
.B(n_133),
.C(n_134),
.Y(n_896)
);

NAND4xp75_ASAP7_75t_L g897 ( 
.A(n_860),
.B(n_135),
.C(n_136),
.D(n_137),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_862),
.A2(n_837),
.B1(n_861),
.B2(n_860),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_SL g899 ( 
.A(n_850),
.B(n_139),
.C(n_141),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_868),
.A2(n_143),
.B(n_144),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_844),
.B(n_145),
.C(n_146),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_841),
.B(n_148),
.C(n_149),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_852),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_857),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_846),
.B(n_150),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_847),
.B(n_151),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_835),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_856),
.B(n_153),
.C(n_155),
.Y(n_909)
);

AO21x2_ASAP7_75t_L g910 ( 
.A1(n_840),
.A2(n_156),
.B(n_157),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_877),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_883),
.Y(n_912)
);

OAI211xp5_ASAP7_75t_SL g913 ( 
.A1(n_853),
.A2(n_158),
.B(n_160),
.C(n_161),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_854),
.B(n_166),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_835),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_881),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_917)
);

NOR2x1_ASAP7_75t_SL g918 ( 
.A(n_882),
.B(n_171),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_873),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_865),
.B(n_172),
.C(n_175),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_888),
.B(n_861),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_908),
.Y(n_922)
);

NAND4xp75_ASAP7_75t_L g923 ( 
.A(n_917),
.B(n_872),
.C(n_865),
.D(n_874),
.Y(n_923)
);

AND4x1_ASAP7_75t_L g924 ( 
.A(n_893),
.B(n_886),
.C(n_875),
.D(n_839),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_888),
.B(n_880),
.Y(n_925)
);

XOR2x2_ASAP7_75t_L g926 ( 
.A(n_898),
.B(n_842),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_911),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_887),
.Y(n_928)
);

XNOR2x2_ASAP7_75t_L g929 ( 
.A(n_899),
.B(n_872),
.Y(n_929)
);

NAND4xp75_ASAP7_75t_L g930 ( 
.A(n_895),
.B(n_870),
.C(n_866),
.D(n_879),
.Y(n_930)
);

XNOR2x2_ASAP7_75t_L g931 ( 
.A(n_889),
.B(n_869),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_910),
.Y(n_932)
);

NAND4xp75_ASAP7_75t_L g933 ( 
.A(n_915),
.B(n_858),
.C(n_878),
.D(n_859),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_887),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_904),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_903),
.Y(n_936)
);

XNOR2xp5_ASAP7_75t_L g937 ( 
.A(n_898),
.B(n_884),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_912),
.B(n_876),
.Y(n_938)
);

NAND4xp75_ASAP7_75t_SL g939 ( 
.A(n_889),
.B(n_878),
.C(n_867),
.D(n_838),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_902),
.A2(n_867),
.B1(n_871),
.B2(n_885),
.Y(n_940)
);

XNOR2x2_ASAP7_75t_L g941 ( 
.A(n_897),
.B(n_176),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_919),
.B(n_177),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_912),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_919),
.B(n_179),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_907),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_892),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_945),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_935),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_927),
.Y(n_950)
);

XOR2x2_ASAP7_75t_L g951 ( 
.A(n_926),
.B(n_920),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_936),
.Y(n_952)
);

XOR2x2_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_894),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_938),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_945),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_931),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_946),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_928),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_934),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_947),
.Y(n_960)
);

XOR2x2_ASAP7_75t_L g961 ( 
.A(n_931),
.B(n_896),
.Y(n_961)
);

XOR2x2_ASAP7_75t_L g962 ( 
.A(n_937),
.B(n_901),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_921),
.B(n_892),
.Y(n_963)
);

OA22x2_ASAP7_75t_L g964 ( 
.A1(n_956),
.A2(n_932),
.B1(n_922),
.B2(n_921),
.Y(n_964)
);

AOI22x1_ASAP7_75t_L g965 ( 
.A1(n_956),
.A2(n_932),
.B1(n_941),
.B2(n_929),
.Y(n_965)
);

XNOR2xp5_ASAP7_75t_L g966 ( 
.A(n_953),
.B(n_923),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_950),
.Y(n_967)
);

OA22x2_ASAP7_75t_L g968 ( 
.A1(n_954),
.A2(n_932),
.B1(n_922),
.B2(n_940),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_949),
.Y(n_969)
);

OAI22x1_ASAP7_75t_L g970 ( 
.A1(n_948),
.A2(n_955),
.B1(n_947),
.B2(n_961),
.Y(n_970)
);

XNOR2xp5_ASAP7_75t_L g971 ( 
.A(n_951),
.B(n_933),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_960),
.Y(n_972)
);

OA22x2_ASAP7_75t_L g973 ( 
.A1(n_951),
.A2(n_943),
.B1(n_925),
.B2(n_894),
.Y(n_973)
);

OA22x2_ASAP7_75t_L g974 ( 
.A1(n_961),
.A2(n_963),
.B1(n_962),
.B2(n_952),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_958),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_962),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_971),
.Y(n_977)
);

AOI322xp5_ASAP7_75t_L g978 ( 
.A1(n_976),
.A2(n_958),
.A3(n_929),
.B1(n_914),
.B2(n_957),
.C1(n_928),
.C2(n_941),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_969),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_975),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_967),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_972),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_971),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_970),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_979),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_977),
.A2(n_965),
.B1(n_966),
.B2(n_974),
.Y(n_986)
);

AO22x2_ASAP7_75t_L g987 ( 
.A1(n_977),
.A2(n_966),
.B1(n_968),
.B2(n_964),
.Y(n_987)
);

OAI31xp33_ASAP7_75t_L g988 ( 
.A1(n_983),
.A2(n_965),
.A3(n_913),
.B(n_909),
.Y(n_988)
);

AND4x1_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_905),
.C(n_906),
.D(n_973),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_985),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_986),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_988),
.A2(n_984),
.B(n_980),
.C(n_978),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_987),
.A2(n_982),
.B1(n_959),
.B2(n_944),
.C(n_942),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_987),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_990),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_991),
.B(n_989),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_994),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_SL g998 ( 
.A1(n_992),
.A2(n_924),
.B1(n_890),
.B2(n_939),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_993),
.A2(n_930),
.B1(n_910),
.B2(n_900),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_910),
.B1(n_900),
.B2(n_906),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_990),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_996),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_995),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_1001),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_905),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1002),
.A2(n_999),
.B1(n_900),
.B2(n_891),
.Y(n_1008)
);

NOR4xp75_ASAP7_75t_L g1009 ( 
.A(n_1003),
.B(n_918),
.C(n_185),
.D(n_186),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1007),
.A2(n_1006),
.B1(n_1005),
.B2(n_1004),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1007),
.A2(n_182),
.B(n_187),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1003),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1003),
.Y(n_1013)
);

AO22x2_ASAP7_75t_L g1014 ( 
.A1(n_1002),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1003),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1014),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1013),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1012),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1015),
.B(n_191),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1010),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_1011),
.B(n_192),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1009),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1008),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1013),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1013),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1014),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1014),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1013),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1013),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1013),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1013),
.B(n_193),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1020),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1022),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1017),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1016),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1026),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1027),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_1023),
.A2(n_204),
.B1(n_206),
.B2(n_208),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_1021),
.Y(n_1039)
);

AO22x2_ASAP7_75t_L g1040 ( 
.A1(n_1024),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1031),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1025),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1028),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1029),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1030),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1018),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1021),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1019),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1039),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1032),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1037),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1034),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1046),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1047),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1041),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1042),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1040),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1043),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1059),
.A2(n_1049),
.B1(n_1035),
.B2(n_1036),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1052),
.A2(n_1038),
.B1(n_1033),
.B2(n_1048),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1054),
.A2(n_1040),
.B1(n_1044),
.B2(n_1045),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_SL g1063 ( 
.A1(n_1051),
.A2(n_1053),
.B1(n_1050),
.B2(n_1058),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1055),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1056),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1062),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1063),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1060),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1064),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1067),
.A2(n_1061),
.B1(n_1057),
.B2(n_1065),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1066),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1070),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1071),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1072),
.A2(n_1068),
.B1(n_1069),
.B2(n_236),
.C(n_237),
.Y(n_1074)
);

AOI211xp5_ASAP7_75t_L g1075 ( 
.A1(n_1074),
.A2(n_1073),
.B(n_238),
.C(n_239),
.Y(n_1075)
);


endmodule