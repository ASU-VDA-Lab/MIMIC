module real_jpeg_7047_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_1),
.B(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_1),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_4),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_5),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_5),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_5),
.B(n_306),
.Y(n_305)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_8),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_9),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_9),
.B(n_27),
.Y(n_223)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_13),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_13),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_14),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_14),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_15),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_15),
.B(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_200),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_198),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_154),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_19),
.B(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.C(n_138),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_20),
.B(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_65),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_21),
.B(n_66),
.C(n_83),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_54),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_22),
.B(n_226),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_22),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_30),
.CI(n_34),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_23),
.B(n_30),
.C(n_34),
.Y(n_153)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_27),
.Y(n_281)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_28),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_36),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_37),
.Y(n_127)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_37),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_38),
.A2(n_54),
.B1(n_55),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_38),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.C(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_39),
.A2(n_51),
.B1(n_176),
.B2(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_40),
.B(n_163),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_40),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_43),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_44),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_45),
.B(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_50),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_51),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_51),
.Y(n_176)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_224)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_59),
.Y(n_300)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_83),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_75),
.C(n_80),
.Y(n_189)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_72),
.Y(n_259)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_75),
.A2(n_82),
.B1(n_123),
.B2(n_124),
.Y(n_264)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_85),
.B(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_84),
.B(n_93),
.C(n_95),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_91),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_96),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_96),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_96),
.B(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_100),
.B(n_138),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_118),
.C(n_120),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_101),
.A2(n_118),
.B1(n_119),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_117),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_107),
.C(n_113),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_105),
.Y(n_245)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_105),
.Y(n_263)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_120),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.C(n_134),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_121),
.A2(n_122),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_337)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_153),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_141),
.C(n_153),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_145),
.C(n_148),
.Y(n_159)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_184),
.B1(n_196),
.B2(n_197),
.Y(n_156)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_173),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_172),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_177),
.A2(n_180),
.B1(n_256),
.B2(n_257),
.Y(n_275)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_180),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_228),
.B(n_345),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_203),
.B(n_205),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_225),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_206),
.A2(n_207),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_210),
.B(n_225),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_224),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_211),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_214),
.B(n_224),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.C(n_223),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_339),
.B(n_344),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_324),
.B(n_338),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_276),
.B(n_323),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_265),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_232),
.B(n_265),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_254),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_250),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_250),
.C(n_254),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_241),
.C(n_246),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_236),
.B1(n_241),
.B2(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_255),
.B(n_333),
.C(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.C(n_275),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_268),
.A2(n_275),
.B1(n_315),
.B2(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_317),
.B(n_322),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_302),
.B(n_316),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_286),
.B(n_301),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_297),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_297),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_292),
.B(n_296),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_292),
.Y(n_296)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_307),
.B(n_310),
.Y(n_318)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B(n_315),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_326),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_332),
.C(n_335),
.Y(n_340)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_341),
.Y(n_344)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);


endmodule