module fake_netlist_6_4302_n_317 (n_52, n_16, n_1, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_317);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_317;

wire n_91;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_125;
wire n_168;
wire n_297;
wire n_106;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_142;
wire n_143;
wire n_180;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_108;
wire n_280;
wire n_287;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_107;
wire n_103;
wire n_272;
wire n_185;
wire n_293;
wire n_232;
wire n_163;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_152;
wire n_92;
wire n_105;
wire n_227;
wire n_132;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_231;
wire n_240;
wire n_139;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_149;
wire n_195;
wire n_285;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_12),
.B(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_14),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_42),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_2),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_4),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_20),
.B(n_3),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_52),
.A2(n_51),
.B1(n_22),
.B2(n_1),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_40),
.A2(n_74),
.B(n_17),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_33),
.A2(n_60),
.B(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_18),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_7),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_5),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_15),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_47),
.B(n_38),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_0),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_30),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_55),
.B(n_6),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_48),
.A2(n_44),
.B1(n_45),
.B2(n_25),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_28),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_16),
.B(n_5),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_26),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_21),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_53),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_86),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_11),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_82),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_145),
.C(n_140),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_115),
.B(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_117),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_155),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_133),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_99),
.B(n_116),
.C(n_119),
.Y(n_185)
);

BUFx6f_ASAP7_75t_SL g186 ( 
.A(n_137),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_L g187 ( 
.A(n_113),
.B(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_154),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_128),
.Y(n_199)
);

AO221x1_ASAP7_75t_L g200 ( 
.A1(n_122),
.A2(n_138),
.B1(n_125),
.B2(n_157),
.C(n_153),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_160),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_135),
.A2(n_158),
.B(n_124),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_102),
.B(n_151),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_102),
.B(n_151),
.Y(n_205)
);

AOI221xp5_ASAP7_75t_L g206 ( 
.A1(n_139),
.A2(n_157),
.B1(n_134),
.B2(n_125),
.C(n_122),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_102),
.B(n_151),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_103),
.B(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_103),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_103),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_199),
.B(n_181),
.C(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_144),
.B1(n_94),
.B2(n_98),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_163),
.B(n_153),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_113),
.B1(n_138),
.B2(n_141),
.Y(n_217)
);

CKINVDCx8_ASAP7_75t_R g218 ( 
.A(n_203),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_178),
.B(n_188),
.C(n_198),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_120),
.B(n_96),
.C(n_100),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_198),
.B(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_113),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

O2A1O1Ixp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_92),
.B(n_105),
.C(n_111),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_138),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_192),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_190),
.A2(n_118),
.B(n_141),
.C(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_189),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_169),
.B(n_205),
.C(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_195),
.B(n_185),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_187),
.A2(n_171),
.B(n_207),
.C(n_185),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_186),
.B(n_166),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_171),
.A2(n_173),
.B(n_199),
.C(n_181),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_139),
.B1(n_206),
.B2(n_181),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_183),
.B(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_165),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_166),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_206),
.B(n_163),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_172),
.B(n_184),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_180),
.B(n_181),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_203),
.A2(n_120),
.B(n_96),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_239),
.B1(n_213),
.B2(n_249),
.Y(n_253)
);

NAND2x1p5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_252),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_227),
.B(n_230),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_222),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_224),
.A2(n_217),
.B1(n_215),
.B2(n_211),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_219),
.B(n_241),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_228),
.B(n_212),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_238),
.B(n_209),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

BUFx2_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_245),
.B1(n_234),
.B2(n_238),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_242),
.B1(n_214),
.B2(n_247),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_233),
.B1(n_248),
.B2(n_274),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

CKINVDCx8_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_270),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_273),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_262),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_264),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_261),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_260),
.C(n_259),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_278),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_254),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_277),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_265),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_268),
.Y(n_301)
);

NAND4xp25_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_272),
.C(n_255),
.D(n_254),
.Y(n_302)
);

AOI211xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_279),
.B(n_288),
.C(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_302),
.B(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_297),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_300),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_295),
.Y(n_311)
);

AOI211xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_301),
.B(n_288),
.C(n_287),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_307),
.Y(n_313)
);

AOI211xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_312),
.B(n_306),
.C(n_285),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_281),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_302),
.Y(n_316)
);

OR2x6_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_308),
.Y(n_317)
);


endmodule