module fake_jpeg_22021_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_1),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_40),
.C(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_21),
.C(n_16),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_51),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_61),
.C(n_19),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_69),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_34),
.C(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_23),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_29),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_18),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_1),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_38),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_31),
.B1(n_28),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_38),
.B1(n_16),
.B2(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_82),
.B1(n_70),
.B2(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_37),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_37),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_122),
.Y(n_137)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g113 ( 
.A(n_109),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_107),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_83),
.A3(n_66),
.B1(n_71),
.B2(n_81),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_90),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_22),
.Y(n_148)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_120),
.Y(n_132)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_85),
.B1(n_79),
.B2(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_72),
.B1(n_62),
.B2(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_125),
.B(n_131),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_72),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_100),
.B1(n_108),
.B2(n_105),
.C(n_32),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_74),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_78),
.B1(n_32),
.B2(n_22),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_148),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_96),
.B1(n_98),
.B2(n_103),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_107),
.B1(n_92),
.B2(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_131),
.B1(n_123),
.B2(n_118),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_140),
.B(n_143),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_94),
.A3(n_104),
.B1(n_102),
.B2(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_114),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_108),
.C(n_37),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.C(n_147),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_2),
.B(n_3),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_32),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_3),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_150),
.B(n_117),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_10),
.C(n_14),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_143),
.C(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_10),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_14),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_153),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_142),
.C(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.C(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_148),
.B1(n_138),
.B2(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_139),
.C(n_144),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_15),
.C(n_9),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_175),
.B(n_164),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_181),
.C(n_13),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_153),
.B1(n_157),
.B2(n_155),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_168),
.B(n_170),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_154),
.B(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_4),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_174),
.B1(n_167),
.B2(n_11),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_185),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_191),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_13),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_197),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_180),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_180),
.B1(n_189),
.B2(n_4),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_188),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_4),
.B1(n_5),
.B2(n_199),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_203),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_201),
.Y(n_205)
);


endmodule