module fake_jpeg_30487_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_38),
.B1(n_5),
.B2(n_4),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_18),
.B1(n_6),
.B2(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_4),
.B1(n_11),
.B2(n_12),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_51),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_74),
.B(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_49),
.C(n_54),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_73),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_47),
.B(n_21),
.C(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_47),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_61),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_61),
.B(n_25),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_66),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_77),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_80),
.B(n_75),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_72),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_29),
.CI(n_28),
.CON(n_88),
.SN(n_88)
);


endmodule