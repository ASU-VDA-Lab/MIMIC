module fake_ariane_268_n_2286 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_381, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_389, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_393, n_359, n_155, n_127, n_2286);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2286;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_436;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_552;
wire n_670;
wire n_1826;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_2075;
wire n_1726;
wire n_699;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1975;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1733;
wire n_1856;
wire n_463;
wire n_1476;
wire n_1524;
wire n_640;
wire n_2016;
wire n_1258;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_586;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_550;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1806;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1777;
wire n_1477;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_1474;
wire n_937;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_311),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_138),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_222),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_308),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_225),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_333),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_201),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_117),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_28),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_188),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_24),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_214),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_353),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_256),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_223),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_306),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_124),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_45),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_289),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_283),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_391),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_373),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_113),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_21),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_139),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_375),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_181),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_6),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_98),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_43),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_298),
.Y(n_428)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_50),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_41),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_2),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_216),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_106),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_91),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_266),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_287),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_178),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_33),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_202),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_203),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_132),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_142),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_326),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_128),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_265),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_310),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_71),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_254),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_4),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_210),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_58),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_365),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_180),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_220),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_161),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_337),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_261),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_341),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_41),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_372),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_163),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_274),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_344),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_123),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_121),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_293),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_183),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_52),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_350),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_89),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_172),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_63),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_47),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_72),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_107),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_385),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_158),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_366),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_354),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_307),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_98),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_338),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_95),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_273),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_94),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_95),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_110),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_329),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_108),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_103),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_340),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_65),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_80),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_251),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_312),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_393),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_131),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_313),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_386),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_381),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_0),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_150),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_115),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_147),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_263),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_57),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_277),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_24),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_46),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_292),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_145),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_208),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_40),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_10),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_130),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_226),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_27),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_302),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_331),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_194),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_320),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_295),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_296),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_215),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_315),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_347),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_280),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_357),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_63),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_318),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_196),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_190),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_327),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_177),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_348),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_314),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_361),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_198),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_22),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_143),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_362),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_75),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_290),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_69),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_89),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_3),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_309),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_179),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_30),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_319),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_170),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_275),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_305),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_352),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_288),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_78),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_83),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_176),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_384),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_269),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_346),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_300),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_377),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_245),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_165),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_371),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_205),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_279),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_299),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_69),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_382),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_243),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_109),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_213),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_33),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_246),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_136),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_378),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_61),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_10),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_102),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_355),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_388),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_247),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_343),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_284),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_29),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_191),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_48),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_155),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_18),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_159),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_16),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_325),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_21),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_78),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_316),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_193),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_133),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_324),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_96),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_252),
.Y(n_605)
);

CKINVDCx14_ASAP7_75t_R g606 ( 
.A(n_167),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_231),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_66),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_140),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_168),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_364),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_282),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_368),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_379),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_211),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_13),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_126),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_370),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_207),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_270),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_141),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_60),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_60),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_358),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_367),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_43),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_212),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_376),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_86),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_152),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_342),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_387),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_239),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_317),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_27),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_91),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_30),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_96),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_339),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_197),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_9),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_334),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_52),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_82),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_359),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_58),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_233),
.Y(n_647)
);

CKINVDCx14_ASAP7_75t_R g648 ( 
.A(n_14),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_230),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_389),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_276),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_356),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_31),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_77),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_104),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_169),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_40),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_227),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_294),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_1),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_285),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_73),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_72),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_74),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_267),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_86),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_84),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_1),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_250),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_257),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_20),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_303),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_291),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_48),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_83),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_236),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_297),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_330),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_304),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_44),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_221),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_157),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_322),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_37),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_146),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_224),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_49),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_0),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_248),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_363),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_101),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_9),
.Y(n_692)
);

BUFx8_ASAP7_75t_SL g693 ( 
.A(n_237),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_262),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_301),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_88),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_74),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_17),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_380),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_35),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_76),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_37),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_160),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_321),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_390),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_28),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_54),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_336),
.Y(n_708)
);

CKINVDCx14_ASAP7_75t_R g709 ( 
.A(n_85),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_187),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_281),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_71),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_260),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_17),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_349),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_323),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_328),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_204),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_173),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_192),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_35),
.Y(n_721)
);

BUFx2_ASAP7_75t_SL g722 ( 
.A(n_3),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_360),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_127),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_199),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_20),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_39),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_88),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_114),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_286),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_335),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_648),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_424),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_420),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_648),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_430),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_693),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_420),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_472),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_438),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_495),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_495),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_511),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_511),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_582),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_693),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_582),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_429),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_429),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_429),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_429),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_429),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_429),
.Y(n_754)
);

INVxp33_ASAP7_75t_SL g755 ( 
.A(n_504),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_405),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_449),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_509),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_410),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_425),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_426),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_461),
.Y(n_762)
);

INVxp33_ASAP7_75t_SL g763 ( 
.A(n_722),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_512),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_470),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_545),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_709),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_486),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_424),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_709),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_517),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_520),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_592),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_622),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_431),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_396),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_416),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_431),
.Y(n_779)
);

INVxp33_ASAP7_75t_SL g780 ( 
.A(n_407),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_641),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_664),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_666),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_667),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_437),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_451),
.Y(n_787)
);

INVxp33_ASAP7_75t_SL g788 ( 
.A(n_414),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_442),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_688),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_692),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_463),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_696),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_702),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_478),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_458),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_714),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_721),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_451),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_635),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_701),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_545),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_545),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_548),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_545),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_490),
.Y(n_810)
);

CKINVDCx16_ASAP7_75t_R g811 ( 
.A(n_527),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_584),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_642),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_655),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_704),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_469),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_435),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_421),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_501),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_643),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_673),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_434),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_434),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_472),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_508),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_508),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_515),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_706),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_421),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_519),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_515),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_652),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_652),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_665),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_665),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_556),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_708),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_708),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_556),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_482),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_482),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_580),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_472),
.B(n_2),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_580),
.Y(n_844)
);

INVxp33_ASAP7_75t_SL g845 ( 
.A(n_439),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_482),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_605),
.Y(n_847)
);

INVxp33_ASAP7_75t_SL g848 ( 
.A(n_453),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_609),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_474),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_620),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_427),
.B(n_4),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_661),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_730),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_445),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_424),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_730),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_690),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_731),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_718),
.Y(n_861)
);

INVxp33_ASAP7_75t_L g862 ( 
.A(n_445),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_731),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_661),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_537),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_731),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_401),
.Y(n_867)
);

CKINVDCx14_ASAP7_75t_R g868 ( 
.A(n_606),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_408),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_411),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_475),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_412),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_419),
.Y(n_873)
);

INVxp33_ASAP7_75t_SL g874 ( 
.A(n_476),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_422),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_432),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_484),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_488),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_433),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_444),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_489),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_529),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_606),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_448),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_456),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_465),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_467),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_471),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_496),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_532),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_477),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_537),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_481),
.Y(n_893)
);

INVxp33_ASAP7_75t_SL g894 ( 
.A(n_516),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_491),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_572),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_547),
.Y(n_897)
);

INVxp33_ASAP7_75t_SL g898 ( 
.A(n_560),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_549),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_492),
.Y(n_900)
);

INVxp33_ASAP7_75t_L g901 ( 
.A(n_572),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_494),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_573),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_503),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_578),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_583),
.Y(n_906)
);

CKINVDCx14_ASAP7_75t_R g907 ( 
.A(n_552),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_506),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_513),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_594),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_514),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_521),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_522),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_535),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_536),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_546),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_598),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_555),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_599),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_567),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_604),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_608),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_569),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_570),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_577),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_585),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_588),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_559),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_595),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_607),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_616),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_615),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_617),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_629),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_424),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_633),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_639),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_645),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_637),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_623),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_649),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_650),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_466),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_628),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_672),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_677),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_679),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_682),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_685),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_705),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_638),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_646),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_716),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_626),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_466),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_725),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_729),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_628),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_653),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_654),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_657),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_660),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_662),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_663),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_675),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_680),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_394),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_684),
.Y(n_968)
);

INVxp33_ASAP7_75t_L g969 ( 
.A(n_651),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_466),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_687),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_697),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_698),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_668),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_700),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_712),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_726),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_727),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_728),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_395),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_397),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_651),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_542),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_656),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_724),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_398),
.Y(n_986)
);

INVxp33_ASAP7_75t_L g987 ( 
.A(n_656),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_703),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_703),
.Y(n_989)
);

XOR2xp5_ASAP7_75t_L g990 ( 
.A(n_671),
.B(n_5),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_720),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_466),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_720),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_447),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_399),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_613),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_596),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_678),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_400),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_402),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_403),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_479),
.Y(n_1002)
);

CKINVDCx14_ASAP7_75t_R g1003 ( 
.A(n_404),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_406),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_413),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_415),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_417),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_418),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_423),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_769),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_749),
.Y(n_1011)
);

OA21x2_ASAP7_75t_L g1012 ( 
.A1(n_750),
.A2(n_436),
.B(n_428),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_751),
.A2(n_443),
.B(n_441),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_769),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_769),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_741),
.B(n_409),
.Y(n_1016)
);

AOI22x1_ASAP7_75t_SL g1017 ( 
.A1(n_890),
.A2(n_446),
.B1(n_452),
.B2(n_450),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_928),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_797),
.B(n_440),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_837),
.B(n_502),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_752),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_1002),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_983),
.Y(n_1023)
);

CKINVDCx11_ASAP7_75t_R g1024 ( 
.A(n_931),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_753),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_983),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_997),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_754),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1002),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_967),
.B(n_589),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_982),
.A2(n_455),
.B(n_454),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_1002),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_934),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_734),
.Y(n_1034)
);

INVx6_ASAP7_75t_L g1035 ( 
.A(n_766),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_766),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_756),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_985),
.Y(n_1038)
);

OA21x2_ASAP7_75t_L g1039 ( 
.A1(n_984),
.A2(n_459),
.B(n_457),
.Y(n_1039)
);

BUFx8_ASAP7_75t_SL g1040 ( 
.A(n_940),
.Y(n_1040)
);

OAI22x1_ASAP7_75t_R g1041 ( 
.A1(n_954),
.A2(n_462),
.B1(n_464),
.B2(n_460),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_734),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_806),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_755),
.A2(n_824),
.B1(n_811),
.B2(n_777),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_822),
.B(n_683),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_738),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_734),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_997),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_843),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_757),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_734),
.Y(n_1051)
);

OAI22x1_ASAP7_75t_SL g1052 ( 
.A1(n_974),
.A2(n_473),
.B1(n_480),
.B2(n_468),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_988),
.A2(n_485),
.B(n_483),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_818),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_760),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_836),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_857),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_758),
.Y(n_1058)
);

INVx6_ASAP7_75t_L g1059 ( 
.A(n_933),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_747),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_877),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_807),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_857),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_989),
.A2(n_493),
.B(n_487),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_878),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_823),
.B(n_479),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_857),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_881),
.Y(n_1068)
);

BUFx8_ASAP7_75t_SL g1069 ( 
.A(n_830),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_857),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_1004),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_809),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_847),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_999),
.B(n_497),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_935),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_844),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_829),
.B(n_498),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_993),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_889),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_897),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_935),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_903),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_935),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_935),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_SL g1085 ( 
.A1(n_859),
.A2(n_500),
.B1(n_507),
.B2(n_499),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_943),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_943),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_853),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_761),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_980),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_824),
.A2(n_518),
.B1(n_523),
.B2(n_510),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_765),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_943),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_759),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_955),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_955),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_905),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_825),
.B(n_479),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_955),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_768),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_981),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_986),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_SL g1104 ( 
.A1(n_778),
.A2(n_525),
.B1(n_526),
.B2(n_524),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_786),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_829),
.B(n_528),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_790),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_958),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_793),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_955),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_883),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_917),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_886),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1000),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_839),
.B(n_530),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_839),
.B(n_531),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_970),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_882),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_867),
.A2(n_870),
.B(n_869),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_970),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_970),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_919),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_796),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_810),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1001),
.B(n_533),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_887),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_826),
.B(n_479),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_842),
.B(n_534),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_771),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_772),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1007),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_970),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_735),
.Y(n_1134)
);

BUFx8_ASAP7_75t_L g1135 ( 
.A(n_740),
.Y(n_1135)
);

CKINVDCx16_ASAP7_75t_R g1136 ( 
.A(n_899),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_739),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_842),
.B(n_864),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_992),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_773),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_992),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_921),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_774),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_780),
.A2(n_538),
.B1(n_540),
.B2(n_539),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_872),
.B(n_505),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_992),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_922),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_827),
.B(n_505),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_992),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1005),
.B(n_543),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_776),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_802),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_803),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_804),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_939),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_805),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_849),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_742),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_744),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_781),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_904),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_873),
.A2(n_550),
.B(n_544),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_782),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_951),
.Y(n_1164)
);

AND2x2_ASAP7_75t_SL g1165 ( 
.A(n_852),
.B(n_505),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_783),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_745),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_864),
.B(n_551),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_733),
.B(n_505),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_851),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_746),
.Y(n_1171)
);

BUFx8_ASAP7_75t_L g1172 ( 
.A(n_831),
.Y(n_1172)
);

BUFx8_ASAP7_75t_SL g1173 ( 
.A(n_861),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_732),
.B(n_553),
.Y(n_1174)
);

AND2x6_ASAP7_75t_L g1175 ( 
.A(n_875),
.B(n_541),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_911),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_748),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_832),
.B(n_541),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_968),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1006),
.B(n_554),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_916),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_920),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_762),
.Y(n_1183)
);

INVxp33_ASAP7_75t_L g1184 ( 
.A(n_817),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_833),
.B(n_541),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_855),
.B(n_557),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_936),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_949),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_950),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_953),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_784),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_971),
.Y(n_1192)
);

BUFx8_ASAP7_75t_L g1193 ( 
.A(n_834),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_785),
.Y(n_1194)
);

BUFx8_ASAP7_75t_L g1195 ( 
.A(n_1095),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1180),
.B(n_1003),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1152),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1138),
.B(n_1008),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1152),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1026),
.B(n_862),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1045),
.B(n_840),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1076),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1186),
.B(n_868),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1158),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1167),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1171),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1177),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1021),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1152),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1021),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1183),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1077),
.B(n_1009),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1120),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1045),
.B(n_841),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1011),
.A2(n_879),
.B(n_876),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1153),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1190),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1153),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1153),
.Y(n_1219)
);

NAND2x1_ASAP7_75t_L g1220 ( 
.A(n_1145),
.B(n_541),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1037),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1055),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1020),
.B(n_846),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1090),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1154),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1154),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1093),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1183),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1154),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1101),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1014),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1027),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1030),
.B(n_591),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1130),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1048),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1156),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1117),
.B(n_901),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1140),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1054),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1023),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1103),
.B(n_978),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1054),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1129),
.B(n_969),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1143),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1151),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1056),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1020),
.B(n_854),
.Y(n_1249)
);

INVxp33_ASAP7_75t_L g1250 ( 
.A(n_1041),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1110),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1160),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1105),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1056),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1163),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1184),
.B(n_987),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1089),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1014),
.Y(n_1258)
);

AND2x2_ASAP7_75t_SL g1259 ( 
.A(n_1169),
.B(n_733),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1168),
.B(n_856),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1165),
.B(n_858),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1014),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1074),
.B(n_860),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1016),
.B(n_817),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1166),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1016),
.B(n_850),
.Y(n_1266)
);

AND2x6_ASAP7_75t_L g1267 ( 
.A(n_1091),
.B(n_591),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1015),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1108),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1019),
.B(n_850),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1113),
.B(n_979),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1126),
.B(n_863),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1015),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1150),
.B(n_866),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_L g1275 ( 
.A(n_1164),
.B(n_959),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1089),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1161),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1025),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1028),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1043),
.A2(n_884),
.B(n_880),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1019),
.B(n_871),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1015),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1043),
.Y(n_1283)
);

NAND2x1_ASAP7_75t_L g1284 ( 
.A(n_1145),
.B(n_591),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1161),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1191),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1036),
.B(n_743),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1194),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1161),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1071),
.B(n_1061),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1194),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1066),
.B(n_743),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1194),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1144),
.A2(n_763),
.B1(n_845),
.B2(n_788),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1066),
.B(n_865),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1065),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1181),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1103),
.B(n_848),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1099),
.B(n_1128),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1059),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1099),
.B(n_835),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1155),
.B(n_874),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1022),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1124),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1078),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1078),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1134),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1181),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1119),
.B(n_736),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1022),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1137),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1159),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1181),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1046),
.B(n_838),
.Y(n_1314)
);

AND2x6_ASAP7_75t_L g1315 ( 
.A(n_1102),
.B(n_591),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1188),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1188),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1125),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1128),
.B(n_865),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1189),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1035),
.B(n_894),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1189),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1079),
.B(n_871),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1189),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1122),
.Y(n_1326)
);

CKINVDCx8_ASAP7_75t_R g1327 ( 
.A(n_1136),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1109),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1114),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1059),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1114),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1080),
.B(n_1098),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1022),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1127),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1032),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1032),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1148),
.B(n_812),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1062),
.A2(n_888),
.B(n_885),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1122),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1127),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1187),
.Y(n_1341)
);

AND2x6_ASAP7_75t_L g1342 ( 
.A(n_1107),
.B(n_600),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1187),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1109),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1123),
.B(n_1142),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1018),
.A2(n_990),
.B1(n_907),
.B2(n_764),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1010),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1029),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1062),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1192),
.B(n_910),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1072),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1072),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1047),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1051),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1216),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1216),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1241),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1300),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1216),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1283),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1283),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_1256),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1219),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1200),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_R g1366 ( 
.A(n_1332),
.B(n_1170),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1221),
.B(n_1155),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1349),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1239),
.B(n_1115),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1198),
.B(n_1162),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1229),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1261),
.A2(n_1174),
.B1(n_813),
.B2(n_815),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1253),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1248),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1254),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1219),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1349),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1219),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1351),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1257),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1276),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1227),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1227),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1351),
.Y(n_1384)
);

BUFx10_ASAP7_75t_L g1385 ( 
.A(n_1322),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1352),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1259),
.A2(n_892),
.B1(n_944),
.B2(n_896),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1352),
.Y(n_1388)
);

NAND2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1345),
.B(n_1179),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1227),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1196),
.A2(n_1132),
.B1(n_1068),
.B2(n_1082),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_SL g1392 ( 
.A(n_1304),
.B(n_1318),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1264),
.B(n_737),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1242),
.B(n_1147),
.C(n_1135),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1211),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1263),
.B(n_1112),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1290),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1208),
.B(n_1162),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1238),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1210),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1245),
.B(n_1272),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1278),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1274),
.B(n_1112),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1212),
.B(n_1112),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1230),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1279),
.B(n_1260),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1233),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1328),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1344),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1266),
.B(n_1050),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1292),
.B(n_1031),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1292),
.B(n_1031),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1217),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1203),
.B(n_1038),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1305),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1215),
.B(n_1039),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1204),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1205),
.Y(n_1419)
);

INVxp33_ASAP7_75t_L g1420 ( 
.A(n_1237),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1206),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1207),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1213),
.A2(n_1013),
.B(n_1012),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1306),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1354),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1354),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1275),
.A2(n_1044),
.B1(n_1012),
.B2(n_1013),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1287),
.B(n_1092),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1243),
.B(n_1269),
.Y(n_1429)
);

AND3x2_ASAP7_75t_L g1430 ( 
.A(n_1309),
.B(n_1058),
.C(n_828),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1294),
.B(n_1148),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1329),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1330),
.B(n_1287),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1267),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1230),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1222),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1223),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1215),
.B(n_1039),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1230),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1331),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1195),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1334),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1324),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1296),
.B(n_1178),
.Y(n_1444)
);

INVxp33_ASAP7_75t_L g1445 ( 
.A(n_1350),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1195),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1340),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1225),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1270),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1341),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1281),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1343),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1353),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1201),
.B(n_910),
.Y(n_1454)
);

NAND2xp33_ASAP7_75t_L g1455 ( 
.A(n_1271),
.B(n_960),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1347),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1251),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1228),
.A2(n_820),
.B1(n_828),
.B2(n_898),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1224),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1231),
.A2(n_820),
.B1(n_896),
.B2(n_892),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1235),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1280),
.B(n_1053),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1224),
.B(n_1178),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1199),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1249),
.B(n_1201),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1236),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1280),
.B(n_1053),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1202),
.B(n_1185),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1240),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1199),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1308),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1214),
.B(n_1060),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1251),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1308),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_SL g1476 ( 
.A(n_1314),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1319),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1288),
.B(n_1185),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1246),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1327),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1319),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1291),
.B(n_961),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1197),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1249),
.B(n_775),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1338),
.B(n_1064),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1247),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1209),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1218),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1214),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1301),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1293),
.B(n_963),
.Y(n_1491)
);

NAND2x1p5_ASAP7_75t_L g1492 ( 
.A(n_1433),
.B(n_1371),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1360),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1457),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1358),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1433),
.B(n_1326),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1428),
.A2(n_1250),
.B1(n_1064),
.B2(n_1252),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1401),
.B(n_1295),
.Y(n_1498)
);

AND2x6_ASAP7_75t_L g1499 ( 
.A(n_1361),
.B(n_1301),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1443),
.B(n_1337),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1395),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1457),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1428),
.A2(n_1255),
.B1(n_1286),
.B2(n_1265),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1368),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1376),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1377),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1401),
.B(n_1369),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1399),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1393),
.B(n_1337),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1369),
.A2(n_1302),
.B1(n_1298),
.B2(n_1299),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1376),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1411),
.B(n_1445),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1425),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1426),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1457),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1473),
.B(n_1466),
.Y(n_1516)
);

AO22x2_ASAP7_75t_L g1517 ( 
.A1(n_1458),
.A2(n_1017),
.B1(n_1104),
.B2(n_1346),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1376),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1358),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1379),
.Y(n_1520)
);

INVxp33_ASAP7_75t_L g1521 ( 
.A(n_1420),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1307),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1384),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1397),
.B(n_1320),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1386),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1383),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1373),
.A2(n_1073),
.B1(n_1314),
.B2(n_1157),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1388),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1357),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1480),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1363),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1383),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1402),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1374),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1383),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1397),
.B(n_1326),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1459),
.B(n_1311),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1484),
.B(n_1312),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1446),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1390),
.Y(n_1541)
);

INVx6_ASAP7_75t_L g1542 ( 
.A(n_1474),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1375),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1390),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1484),
.B(n_952),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1380),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1490),
.B(n_1313),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1355),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1436),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1381),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1449),
.B(n_952),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1489),
.B(n_1316),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1414),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1489),
.B(n_1317),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1418),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1362),
.B(n_1173),
.Y(n_1556)
);

BUFx8_ASAP7_75t_SL g1557 ( 
.A(n_1441),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1437),
.Y(n_1558)
);

NAND2xp33_ASAP7_75t_SL g1559 ( 
.A(n_1407),
.B(n_964),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1451),
.B(n_962),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1419),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1448),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1365),
.B(n_962),
.Y(n_1563)
);

AND2x6_ASAP7_75t_L g1564 ( 
.A(n_1412),
.B(n_1226),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1408),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1407),
.B(n_1234),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1387),
.B(n_794),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1406),
.B(n_1234),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1421),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1406),
.B(n_1234),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1400),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1422),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1416),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1366),
.B(n_1033),
.C(n_1135),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1409),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1454),
.B(n_816),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1424),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1461),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1467),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1476),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1470),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1430),
.B(n_1321),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1476),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1385),
.B(n_1069),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1430),
.B(n_1323),
.Y(n_1585)
);

INVx5_ASAP7_75t_L g1586 ( 
.A(n_1434),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_L g1587 ( 
.A(n_1479),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1486),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1432),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1578),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1507),
.B(n_1387),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1521),
.B(n_1385),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1498),
.B(n_1370),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1500),
.Y(n_1594)
);

AND2x6_ASAP7_75t_SL g1595 ( 
.A(n_1584),
.B(n_1040),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1559),
.A2(n_1415),
.B(n_1367),
.C(n_1427),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1391),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1587),
.B(n_1392),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1578),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1586),
.B(n_1434),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1567),
.A2(n_770),
.B1(n_767),
.B2(n_1458),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1524),
.B(n_1545),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1509),
.A2(n_1024),
.B1(n_1049),
.B2(n_1464),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1512),
.B(n_1415),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1561),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1494),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1510),
.B(n_1431),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1431),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1493),
.B(n_1370),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1569),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1516),
.B(n_1367),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1572),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1513),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1494),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1493),
.B(n_1440),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1579),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1579),
.B(n_1460),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1504),
.A2(n_1447),
.B1(n_1450),
.B2(n_1442),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1516),
.A2(n_1366),
.B1(n_1389),
.B2(n_1429),
.Y(n_1621)
);

NAND2x1_ASAP7_75t_L g1622 ( 
.A(n_1532),
.B(n_1355),
.Y(n_1622)
);

INVx8_ASAP7_75t_L g1623 ( 
.A(n_1494),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1556),
.A2(n_1460),
.B1(n_1394),
.B2(n_1404),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1502),
.B(n_1452),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1515),
.B(n_1464),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1514),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1501),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1539),
.B(n_1404),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_L g1630 ( 
.A(n_1574),
.B(n_1396),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1551),
.B(n_1444),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1504),
.B(n_1412),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1506),
.B(n_1413),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1506),
.B(n_1413),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1589),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1542),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1539),
.B(n_1522),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1563),
.B(n_1444),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1520),
.B(n_1410),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1492),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1396),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1520),
.B(n_1398),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1523),
.B(n_1398),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1499),
.A2(n_1403),
.B1(n_1033),
.B2(n_1469),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1523),
.B(n_1482),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1560),
.B(n_1403),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1589),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1575),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1508),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1623),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1597),
.A2(n_1499),
.B1(n_1527),
.B2(n_1517),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1642),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1591),
.B(n_1525),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1594),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1635),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1581),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1647),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

INVx4_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1629),
.Y(n_1662)
);

CKINVDCx6p67_ASAP7_75t_R g1663 ( 
.A(n_1623),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1601),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1642),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1627),
.Y(n_1666)
);

BUFx4f_ASAP7_75t_L g1667 ( 
.A(n_1601),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1599),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1608),
.Y(n_1670)
);

BUFx12f_ASAP7_75t_SL g1671 ( 
.A(n_1608),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

BUFx4f_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1616),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1610),
.B(n_1581),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1606),
.B(n_1588),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1602),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1625),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1631),
.B(n_1588),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1607),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1590),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1600),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx5_ASAP7_75t_L g1685 ( 
.A(n_1616),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1625),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1603),
.A2(n_1517),
.B1(n_1497),
.B2(n_1049),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1640),
.Y(n_1688)
);

BUFx4f_ASAP7_75t_L g1689 ( 
.A(n_1626),
.Y(n_1689)
);

AOI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1591),
.A2(n_1372),
.B(n_1491),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1612),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1655),
.B(n_1638),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1672),
.B(n_1592),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1682),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1655),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1679),
.B(n_1618),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1672),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1679),
.B(n_1626),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1668),
.B(n_1630),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1663),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1664),
.A2(n_1611),
.B(n_1423),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1653),
.A2(n_1593),
.B(n_1611),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1665),
.A2(n_1593),
.B(n_1596),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1619),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1690),
.A2(n_1624),
.B(n_1621),
.C(n_1641),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1673),
.A2(n_1649),
.B(n_1645),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1673),
.A2(n_1649),
.B(n_1645),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1667),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1652),
.B(n_1557),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1668),
.B(n_1598),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1684),
.B(n_1632),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1687),
.A2(n_1644),
.B(n_1613),
.C(n_1676),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1689),
.B(n_1620),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1667),
.B(n_1586),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1689),
.B(n_1620),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1684),
.A2(n_1633),
.B(n_1632),
.Y(n_1718)
);

BUFx10_ASAP7_75t_L g1719 ( 
.A(n_1651),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1663),
.Y(n_1720)
);

AO32x2_ASAP7_75t_L g1721 ( 
.A1(n_1686),
.A2(n_1583),
.A3(n_1580),
.B1(n_1532),
.B2(n_1535),
.Y(n_1721)
);

AND3x4_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1540),
.C(n_1530),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1659),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1657),
.B(n_1017),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1654),
.B(n_1633),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1654),
.B(n_1634),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_SL g1727 ( 
.A(n_1685),
.B(n_1634),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_SL g1728 ( 
.A1(n_1683),
.A2(n_1455),
.B(n_1491),
.C(n_1503),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1661),
.B(n_1646),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1656),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1656),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1661),
.B(n_1628),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1709),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1694),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1722),
.Y(n_1735)
);

BUFx8_ASAP7_75t_SL g1736 ( 
.A(n_1720),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1695),
.Y(n_1737)
);

CKINVDCx8_ASAP7_75t_R g1738 ( 
.A(n_1697),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1706),
.A2(n_1677),
.B(n_1680),
.C(n_1617),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1605),
.B1(n_1691),
.B2(n_1669),
.Y(n_1740)
);

BUFx2_ASAP7_75t_SL g1741 ( 
.A(n_1701),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1693),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1711),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1692),
.B(n_1104),
.Y(n_1745)
);

BUFx8_ASAP7_75t_L g1746 ( 
.A(n_1721),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1700),
.B(n_1658),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1705),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1704),
.B(n_1662),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1732),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1730),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1723),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1729),
.Y(n_1753)
);

AND2x2_ASAP7_75t_SL g1754 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1696),
.B(n_1662),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1731),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1725),
.B(n_1617),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1698),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1715),
.A2(n_1499),
.B1(n_1689),
.B2(n_1234),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1710),
.B(n_1595),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1714),
.A2(n_1528),
.B1(n_1573),
.B2(n_1571),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1705),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1725),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1726),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1713),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1726),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1717),
.A2(n_1666),
.B1(n_1678),
.B2(n_1669),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1713),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1698),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1710),
.B(n_1085),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1699),
.A2(n_1691),
.B1(n_1678),
.B2(n_1681),
.Y(n_1773)
);

OAI33xp33_ASAP7_75t_L g1774 ( 
.A1(n_1728),
.A2(n_795),
.A3(n_791),
.B1(n_798),
.B2(n_792),
.B3(n_789),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1737),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1759),
.A2(n_1708),
.B1(n_1707),
.B2(n_1674),
.Y(n_1776)
);

AO31x2_ASAP7_75t_L g1777 ( 
.A1(n_1762),
.A2(n_1727),
.A3(n_1703),
.B(n_1718),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1739),
.A2(n_1712),
.B(n_972),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1749),
.A2(n_1667),
.B(n_1674),
.Y(n_1779)
);

AOI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1762),
.A2(n_1702),
.B(n_1712),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1739),
.A2(n_808),
.B(n_972),
.C(n_906),
.Y(n_1781)
);

CKINVDCx11_ASAP7_75t_R g1782 ( 
.A(n_1738),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1734),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1742),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1764),
.B(n_891),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1770),
.B(n_893),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1745),
.A2(n_1499),
.B1(n_1668),
.B2(n_1585),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1749),
.A2(n_1570),
.B(n_1568),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1749),
.A2(n_1774),
.B(n_1748),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1737),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1765),
.B(n_895),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1772),
.A2(n_906),
.B(n_1537),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1735),
.B(n_1580),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1751),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1756),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1740),
.A2(n_821),
.B(n_819),
.C(n_814),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1774),
.A2(n_1716),
.B(n_1566),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1735),
.B(n_1583),
.Y(n_1798)
);

AO32x2_ASAP7_75t_L g1799 ( 
.A1(n_1753),
.A2(n_1688),
.A3(n_1670),
.B1(n_1651),
.B2(n_1660),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1744),
.A2(n_1668),
.B1(n_1716),
.B2(n_1685),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1733),
.Y(n_1801)
);

AO31x2_ASAP7_75t_L g1802 ( 
.A1(n_1743),
.A2(n_1681),
.A3(n_1438),
.B(n_1417),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1743),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1760),
.A2(n_944),
.B(n_991),
.C(n_808),
.Y(n_1804)
);

O2A1O1Ixp33_ASAP7_75t_L g1805 ( 
.A1(n_1757),
.A2(n_991),
.B(n_779),
.C(n_787),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1750),
.B(n_1719),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1747),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1757),
.A2(n_1685),
.B(n_1639),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1754),
.A2(n_1685),
.B(n_1639),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1747),
.A2(n_1685),
.B(n_1670),
.Y(n_1810)
);

OAI21x1_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1664),
.B(n_1438),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1755),
.A2(n_1670),
.B(n_1664),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1752),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1755),
.A2(n_1622),
.B(n_1675),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1766),
.Y(n_1815)
);

O2A1O1Ixp33_ASAP7_75t_SL g1816 ( 
.A1(n_1769),
.A2(n_1736),
.B(n_1735),
.C(n_1767),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1763),
.B(n_900),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1768),
.A2(n_908),
.B(n_902),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1750),
.B(n_909),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1761),
.A2(n_779),
.B(n_787),
.C(n_775),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1761),
.A2(n_1668),
.B1(n_1582),
.B2(n_1585),
.Y(n_1821)
);

O2A1O1Ixp33_ASAP7_75t_SL g1822 ( 
.A1(n_1741),
.A2(n_966),
.B(n_973),
.C(n_965),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1771),
.B(n_1671),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1773),
.A2(n_801),
.B(n_996),
.C(n_994),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1746),
.A2(n_1582),
.B1(n_1614),
.B2(n_1648),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1758),
.A2(n_1688),
.B1(n_1675),
.B2(n_1660),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1746),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1758),
.Y(n_1828)
);

AO31x2_ASAP7_75t_L g1829 ( 
.A1(n_1758),
.A2(n_1468),
.A3(n_1485),
.B(n_1462),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1762),
.A2(n_1485),
.B(n_1359),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1749),
.A2(n_1675),
.B(n_1528),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1739),
.A2(n_913),
.B(n_912),
.Y(n_1832)
);

A2O1A1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1739),
.A2(n_914),
.B(n_918),
.C(n_915),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1746),
.A2(n_1650),
.B1(n_1564),
.B2(n_1487),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1734),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1827),
.A2(n_1193),
.B1(n_1172),
.B2(n_1052),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1819),
.A2(n_1542),
.B1(n_998),
.B2(n_801),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1784),
.A2(n_1675),
.B1(n_1660),
.B2(n_1573),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1783),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1775),
.B(n_1675),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1781),
.A2(n_800),
.B1(n_799),
.B2(n_924),
.C(n_923),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1825),
.A2(n_1193),
.B1(n_1172),
.B2(n_1571),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1782),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1778),
.A2(n_1577),
.B1(n_1549),
.B2(n_1562),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1793),
.Y(n_1845)
);

OAI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1786),
.A2(n_1577),
.B1(n_926),
.B2(n_927),
.Y(n_1846)
);

CKINVDCx16_ASAP7_75t_R g1847 ( 
.A(n_1798),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_SL g1848 ( 
.A1(n_1816),
.A2(n_976),
.B(n_977),
.C(n_975),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1806),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1787),
.A2(n_1522),
.B1(n_1533),
.B2(n_1552),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1828),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1776),
.A2(n_1558),
.B1(n_1519),
.B2(n_1495),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1822),
.B(n_1823),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1785),
.B(n_5),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1789),
.A2(n_1535),
.B1(n_1526),
.B2(n_1511),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1835),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1790),
.B(n_1495),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1794),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1795),
.B(n_1519),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1834),
.A2(n_1564),
.B1(n_1488),
.B2(n_1483),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1811),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1801),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1815),
.Y(n_1863)
);

NAND2x1_ASAP7_75t_L g1864 ( 
.A(n_1803),
.B(n_1505),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1780),
.A2(n_1518),
.B(n_1505),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1807),
.A2(n_1564),
.B1(n_1315),
.B2(n_1342),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1813),
.A2(n_1564),
.B1(n_1315),
.B2(n_1342),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1831),
.A2(n_1548),
.B1(n_1544),
.B2(n_1518),
.Y(n_1868)
);

BUFx12f_ASAP7_75t_L g1869 ( 
.A(n_1792),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1799),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1779),
.A2(n_1511),
.B1(n_1536),
.B2(n_1526),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1821),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1791),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1799),
.B(n_1721),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1808),
.B(n_925),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1799),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1797),
.A2(n_1315),
.B1(n_1342),
.B2(n_1267),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1810),
.B(n_929),
.Y(n_1878)
);

OAI222xp33_ASAP7_75t_L g1879 ( 
.A1(n_1817),
.A2(n_1543),
.B1(n_1531),
.B2(n_1546),
.C1(n_1534),
.C2(n_1529),
.Y(n_1879)
);

OAI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1832),
.A2(n_1511),
.B1(n_1536),
.B2(n_1526),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1777),
.B(n_1721),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1845),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1861),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1870),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1839),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1849),
.B(n_1777),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1861),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1876),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1874),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1881),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1856),
.B(n_1830),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1858),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1861),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1865),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1840),
.B(n_1802),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1862),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1869),
.A2(n_1809),
.B1(n_1818),
.B2(n_1812),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1859),
.Y(n_1898)
);

AO21x2_ASAP7_75t_L g1899 ( 
.A1(n_1875),
.A2(n_1788),
.B(n_1796),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1873),
.Y(n_1900)
);

AO31x2_ASAP7_75t_L g1901 ( 
.A1(n_1868),
.A2(n_1833),
.A3(n_1814),
.B(n_1804),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1854),
.A2(n_1805),
.B(n_1824),
.C(n_1826),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1863),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1851),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1864),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1840),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1855),
.A2(n_1315),
.B1(n_1342),
.B2(n_1267),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1847),
.B(n_1802),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1844),
.A2(n_1800),
.B1(n_1820),
.B2(n_1548),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1853),
.A2(n_1544),
.B1(n_1536),
.B2(n_1541),
.Y(n_1910)
);

OAI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1890),
.A2(n_1889),
.B1(n_1884),
.B2(n_1908),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1899),
.A2(n_1908),
.B1(n_1889),
.B2(n_1890),
.Y(n_1912)
);

OA21x2_ASAP7_75t_L g1913 ( 
.A1(n_1884),
.A2(n_1878),
.B(n_1859),
.Y(n_1913)
);

OR2x6_ASAP7_75t_L g1914 ( 
.A(n_1900),
.B(n_1843),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_SL g1915 ( 
.A1(n_1899),
.A2(n_1872),
.B1(n_1852),
.B2(n_1846),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1885),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1882),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1897),
.A2(n_1836),
.B(n_1838),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1888),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1899),
.A2(n_1842),
.B1(n_1837),
.B2(n_1860),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1902),
.A2(n_1848),
.B1(n_1850),
.B2(n_1841),
.C(n_1877),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1896),
.Y(n_1922)
);

OAI211xp5_ASAP7_75t_L g1923 ( 
.A1(n_1886),
.A2(n_1843),
.B(n_1850),
.C(n_932),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1890),
.A2(n_1857),
.B1(n_1880),
.B2(n_1871),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1898),
.B(n_1857),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1900),
.A2(n_1866),
.B1(n_1277),
.B2(n_1289),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1883),
.A2(n_1879),
.B(n_1867),
.Y(n_1927)
);

OR2x6_ASAP7_75t_L g1928 ( 
.A(n_1886),
.B(n_1541),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_SL g1929 ( 
.A1(n_1895),
.A2(n_938),
.B1(n_941),
.B2(n_937),
.C(n_930),
.Y(n_1929)
);

OAI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1898),
.A2(n_945),
.B(n_946),
.C(n_942),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1888),
.A2(n_1285),
.B1(n_1325),
.B2(n_1297),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1909),
.A2(n_1550),
.B1(n_1267),
.B2(n_1338),
.Y(n_1932)
);

OAI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1910),
.A2(n_611),
.B1(n_689),
.B2(n_600),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1895),
.A2(n_1538),
.B1(n_1456),
.B2(n_1463),
.Y(n_1934)
);

NAND2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1898),
.B(n_1586),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1903),
.B(n_947),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1916),
.B(n_1885),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1925),
.B(n_1898),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1919),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1914),
.B(n_1913),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1913),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1923),
.A2(n_1887),
.B1(n_1893),
.B2(n_1883),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1914),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1914),
.B(n_1906),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1928),
.B(n_1905),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1912),
.B(n_1906),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1922),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1917),
.B(n_1904),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1915),
.B(n_1892),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1911),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1927),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1936),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1928),
.B(n_1904),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1928),
.Y(n_1954)
);

AND2x4_ASAP7_75t_SL g1955 ( 
.A(n_1934),
.B(n_1903),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1931),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1935),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1924),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1921),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1935),
.B(n_1905),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1918),
.B(n_1905),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1923),
.B(n_1892),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1920),
.B(n_1891),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1929),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1930),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1933),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1932),
.B(n_1891),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1926),
.B(n_1883),
.Y(n_1968)
);

AOI211x1_ASAP7_75t_L g1969 ( 
.A1(n_1949),
.A2(n_1921),
.B(n_956),
.C(n_957),
.Y(n_1969)
);

OR2x6_ASAP7_75t_L g1970 ( 
.A(n_1959),
.B(n_1894),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1952),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1937),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1952),
.A2(n_1883),
.B1(n_1893),
.B2(n_1887),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1944),
.B(n_1887),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1944),
.B(n_1887),
.Y(n_1975)
);

AND2x4_ASAP7_75t_SL g1976 ( 
.A(n_1943),
.B(n_1893),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1939),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1959),
.A2(n_1893),
.B1(n_1894),
.B2(n_1896),
.C(n_1907),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1964),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1937),
.Y(n_1980)
);

AOI33xp33_ASAP7_75t_L g1981 ( 
.A1(n_1958),
.A2(n_948),
.A3(n_1894),
.B1(n_8),
.B2(n_11),
.B3(n_12),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1948),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1939),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1948),
.B(n_1901),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1958),
.A2(n_1963),
.B1(n_1961),
.B2(n_1951),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1962),
.B(n_1901),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1963),
.A2(n_1961),
.B1(n_1951),
.B2(n_1965),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1965),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1938),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1955),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1971),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1982),
.B(n_1938),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1977),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1979),
.B(n_1941),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1977),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1971),
.Y(n_1996)
);

NAND2x1p5_ASAP7_75t_L g1997 ( 
.A(n_1984),
.B(n_1940),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1989),
.B(n_1940),
.Y(n_1998)
);

OR2x6_ASAP7_75t_SL g1999 ( 
.A(n_1988),
.B(n_1941),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1981),
.B(n_1950),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1972),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1974),
.B(n_1953),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1990),
.B(n_1980),
.Y(n_2003)
);

BUFx5_ASAP7_75t_L g2004 ( 
.A(n_1984),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1983),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_L g2006 ( 
.A1(n_2000),
.A2(n_1987),
.B(n_1985),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1991),
.B(n_1976),
.Y(n_2007)
);

NAND3xp33_ASAP7_75t_L g2008 ( 
.A(n_1996),
.B(n_1987),
.C(n_1981),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_2002),
.B(n_1992),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2005),
.B(n_1969),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_2003),
.B(n_1975),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2004),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1998),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1994),
.B(n_1986),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_2009),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_2006),
.B(n_1993),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_2011),
.B(n_2003),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2013),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_2014),
.B(n_2001),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2008),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2012),
.Y(n_2021)
);

OAI31xp33_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_1985),
.A3(n_2010),
.B(n_1997),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_2017),
.B(n_2007),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_2015),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_2019),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_L g2026 ( 
.A(n_2018),
.B(n_2007),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2026),
.B(n_2001),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_2023),
.B(n_2021),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2025),
.A2(n_2016),
.B1(n_2004),
.B2(n_1970),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2028),
.B(n_2024),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_2027),
.B(n_2023),
.Y(n_2031)
);

AO21x1_ASAP7_75t_L g2032 ( 
.A1(n_2030),
.A2(n_2016),
.B(n_2022),
.Y(n_2032)
);

OAI332xp33_ASAP7_75t_L g2033 ( 
.A1(n_2031),
.A2(n_1993),
.A3(n_1995),
.B1(n_2029),
.B2(n_1999),
.B3(n_1950),
.C1(n_1978),
.C2(n_2004),
.Y(n_2033)
);

OAI322xp33_ASAP7_75t_L g2034 ( 
.A1(n_2030),
.A2(n_2004),
.A3(n_1966),
.B1(n_1973),
.B2(n_1946),
.C1(n_1954),
.C2(n_1967),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_2032),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_2033),
.B(n_1976),
.Y(n_2036)
);

AOI221xp5_ASAP7_75t_SL g2037 ( 
.A1(n_2035),
.A2(n_2034),
.B1(n_2004),
.B2(n_1953),
.C(n_1966),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2035),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2036),
.A2(n_1966),
.B(n_1946),
.C(n_1960),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_2038),
.B(n_1970),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_2037),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2039),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_2038),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2041),
.B(n_1970),
.Y(n_2044)
);

NOR2x1_ASAP7_75t_L g2045 ( 
.A(n_2042),
.B(n_1538),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2043),
.B(n_2040),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_SL g2047 ( 
.A(n_2043),
.B(n_1966),
.Y(n_2047)
);

O2A1O1Ixp33_ASAP7_75t_L g2048 ( 
.A1(n_2046),
.A2(n_1496),
.B(n_1954),
.C(n_1469),
.Y(n_2048)
);

AOI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2044),
.A2(n_1966),
.B(n_1960),
.C(n_1967),
.Y(n_2049)
);

XNOR2x1_ASAP7_75t_L g2050 ( 
.A(n_2045),
.B(n_6),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2047),
.A2(n_1954),
.B1(n_1947),
.B2(n_1945),
.Y(n_2051)
);

AOI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_2044),
.A2(n_1947),
.B1(n_1956),
.B2(n_1955),
.C(n_1945),
.Y(n_2052)
);

AO21x1_ASAP7_75t_L g2053 ( 
.A1(n_2046),
.A2(n_1945),
.B(n_7),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_SL g2054 ( 
.A1(n_2044),
.A2(n_1957),
.B1(n_1968),
.B2(n_1035),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_2044),
.B(n_1942),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_2044),
.B(n_1957),
.Y(n_2056)
);

NOR2x1p5_ASAP7_75t_L g2057 ( 
.A(n_2044),
.B(n_7),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2044),
.A2(n_1968),
.B1(n_1547),
.B2(n_1554),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2044),
.A2(n_1547),
.B1(n_1554),
.B2(n_1552),
.Y(n_2059)
);

NAND2xp33_ASAP7_75t_L g2060 ( 
.A(n_2046),
.B(n_8),
.Y(n_2060)
);

A2O1A1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_2044),
.A2(n_1182),
.B(n_1176),
.C(n_1478),
.Y(n_2061)
);

NAND3xp33_ASAP7_75t_SL g2062 ( 
.A(n_2053),
.B(n_561),
.C(n_558),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_L g2063 ( 
.A(n_2060),
.B(n_1182),
.C(n_1176),
.Y(n_2063)
);

OA22x2_ASAP7_75t_L g2064 ( 
.A1(n_2055),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_2056),
.B(n_1176),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_L g2066 ( 
.A(n_2061),
.B(n_1339),
.C(n_1478),
.Y(n_2066)
);

NOR2xp67_ASAP7_75t_L g2067 ( 
.A(n_2051),
.B(n_14),
.Y(n_2067)
);

NOR3xp33_ASAP7_75t_L g2068 ( 
.A(n_2054),
.B(n_1339),
.C(n_1284),
.Y(n_2068)
);

NAND2x1p5_ASAP7_75t_L g2069 ( 
.A(n_2057),
.B(n_1356),
.Y(n_2069)
);

NOR4xp25_ASAP7_75t_L g2070 ( 
.A(n_2048),
.B(n_1471),
.C(n_1465),
.D(n_18),
.Y(n_2070)
);

NOR3xp33_ASAP7_75t_L g2071 ( 
.A(n_2052),
.B(n_1220),
.C(n_563),
.Y(n_2071)
);

NAND4xp25_ASAP7_75t_L g2072 ( 
.A(n_2049),
.B(n_19),
.C(n_15),
.D(n_16),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_2059),
.B(n_564),
.C(n_562),
.Y(n_2073)
);

AOI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_2058),
.A2(n_1182),
.B1(n_568),
.B2(n_571),
.C(n_566),
.Y(n_2074)
);

AOI21xp33_ASAP7_75t_L g2075 ( 
.A1(n_2050),
.A2(n_15),
.B(n_19),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2053),
.B(n_22),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2061),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2053),
.Y(n_2078)
);

O2A1O1Ixp33_ASAP7_75t_L g2079 ( 
.A1(n_2060),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_L g2080 ( 
.A(n_2060),
.B(n_574),
.C(n_565),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2053),
.B(n_29),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_L g2082 ( 
.A(n_2060),
.B(n_576),
.C(n_575),
.Y(n_2082)
);

NOR3xp33_ASAP7_75t_L g2083 ( 
.A(n_2060),
.B(n_581),
.C(n_579),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_L g2084 ( 
.A(n_2060),
.B(n_587),
.C(n_586),
.Y(n_2084)
);

NOR3xp33_ASAP7_75t_L g2085 ( 
.A(n_2060),
.B(n_597),
.C(n_593),
.Y(n_2085)
);

AOI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_2055),
.A2(n_602),
.B1(n_610),
.B2(n_603),
.C(n_601),
.Y(n_2086)
);

O2A1O1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_2060),
.A2(n_34),
.B(n_31),
.C(n_32),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_L g2088 ( 
.A(n_2060),
.B(n_614),
.C(n_612),
.Y(n_2088)
);

NAND4xp75_ASAP7_75t_L g2089 ( 
.A(n_2053),
.B(n_36),
.C(n_32),
.D(n_34),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_2055),
.A2(n_676),
.B1(n_723),
.B2(n_618),
.C(n_619),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2057),
.B(n_36),
.Y(n_2091)
);

NOR2x1_ASAP7_75t_L g2092 ( 
.A(n_2060),
.B(n_38),
.Y(n_2092)
);

NAND5xp2_ASAP7_75t_L g2093 ( 
.A(n_2054),
.B(n_38),
.C(n_39),
.D(n_42),
.E(n_44),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_2060),
.B(n_42),
.Y(n_2094)
);

NOR2x1_ASAP7_75t_L g2095 ( 
.A(n_2060),
.B(n_45),
.Y(n_2095)
);

NAND3xp33_ASAP7_75t_L g2096 ( 
.A(n_2060),
.B(n_624),
.C(n_621),
.Y(n_2096)
);

NOR3x1_ASAP7_75t_L g2097 ( 
.A(n_2055),
.B(n_46),
.C(n_47),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_2053),
.B(n_600),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2053),
.Y(n_2099)
);

INVxp67_ASAP7_75t_SL g2100 ( 
.A(n_2057),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2076),
.A2(n_1475),
.B1(n_1477),
.B2(n_1472),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2078),
.A2(n_2099),
.B1(n_2062),
.B2(n_2083),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2081),
.A2(n_627),
.B1(n_630),
.B2(n_625),
.Y(n_2103)
);

AOI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2100),
.A2(n_49),
.B(n_50),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2091),
.B(n_51),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_SL g2106 ( 
.A(n_2098),
.B(n_632),
.C(n_631),
.Y(n_2106)
);

XNOR2xp5_ASAP7_75t_L g2107 ( 
.A(n_2089),
.B(n_2091),
.Y(n_2107)
);

OA22x2_ASAP7_75t_L g2108 ( 
.A1(n_2077),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_2108)
);

OAI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_2086),
.A2(n_56),
.B(n_53),
.C(n_55),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2082),
.A2(n_1481),
.B1(n_640),
.B2(n_647),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2092),
.Y(n_2111)
);

NOR4xp25_ASAP7_75t_L g2112 ( 
.A(n_2090),
.B(n_57),
.C(n_55),
.D(n_56),
.Y(n_2112)
);

OAI211xp5_ASAP7_75t_SL g2113 ( 
.A1(n_2074),
.A2(n_62),
.B(n_59),
.C(n_61),
.Y(n_2113)
);

AOI31xp33_ASAP7_75t_L g2114 ( 
.A1(n_2080),
.A2(n_64),
.A3(n_59),
.B(n_62),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2094),
.Y(n_2115)
);

AOI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2075),
.A2(n_691),
.B1(n_717),
.B2(n_634),
.C(n_658),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2095),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2067),
.B(n_64),
.Y(n_2118)
);

AO22x2_ASAP7_75t_SL g2119 ( 
.A1(n_2084),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2069),
.B(n_67),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2097),
.Y(n_2121)
);

OAI211xp5_ASAP7_75t_L g2122 ( 
.A1(n_2072),
.A2(n_2087),
.B(n_2079),
.C(n_2085),
.Y(n_2122)
);

NAND3xp33_ASAP7_75t_L g2123 ( 
.A(n_2088),
.B(n_611),
.C(n_600),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2096),
.B(n_669),
.C(n_659),
.Y(n_2124)
);

OAI211xp5_ASAP7_75t_L g2125 ( 
.A1(n_2073),
.A2(n_73),
.B(n_68),
.C(n_70),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2063),
.A2(n_681),
.B(n_670),
.Y(n_2126)
);

AOI321xp33_ASAP7_75t_L g2127 ( 
.A1(n_2070),
.A2(n_68),
.A3(n_70),
.B1(n_75),
.B2(n_76),
.C(n_77),
.Y(n_2127)
);

NAND4xp25_ASAP7_75t_SL g2128 ( 
.A(n_2071),
.B(n_81),
.C(n_79),
.D(n_80),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2093),
.A2(n_699),
.B1(n_686),
.B2(n_715),
.C(n_694),
.Y(n_2129)
);

AOI311xp33_ASAP7_75t_L g2130 ( 
.A1(n_2065),
.A2(n_79),
.A3(n_81),
.B(n_82),
.C(n_84),
.Y(n_2130)
);

OAI211xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2068),
.A2(n_85),
.B(n_87),
.C(n_90),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_SL g2132 ( 
.A(n_2066),
.B(n_710),
.C(n_695),
.Y(n_2132)
);

NAND2x1p5_ASAP7_75t_L g2133 ( 
.A(n_2064),
.B(n_1356),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2076),
.A2(n_713),
.B1(n_719),
.B2(n_1541),
.Y(n_2134)
);

NAND3xp33_ASAP7_75t_SL g2135 ( 
.A(n_2078),
.B(n_87),
.C(n_90),
.Y(n_2135)
);

NAND3xp33_ASAP7_75t_SL g2136 ( 
.A(n_2078),
.B(n_92),
.C(n_93),
.Y(n_2136)
);

BUFx2_ASAP7_75t_L g2137 ( 
.A(n_2091),
.Y(n_2137)
);

AO22x2_ASAP7_75t_L g2138 ( 
.A1(n_2078),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_2138)
);

OAI211xp5_ASAP7_75t_SL g2139 ( 
.A1(n_2078),
.A2(n_97),
.B(n_1439),
.C(n_1435),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2078),
.A2(n_1434),
.B1(n_1359),
.B2(n_1439),
.Y(n_2140)
);

XNOR2x2_ASAP7_75t_L g2141 ( 
.A(n_2089),
.B(n_97),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2081),
.Y(n_2142)
);

AOI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_2078),
.A2(n_611),
.B1(n_711),
.B2(n_689),
.C(n_1405),
.Y(n_2143)
);

AOI311xp33_ASAP7_75t_L g2144 ( 
.A1(n_2078),
.A2(n_99),
.A3(n_100),
.B(n_105),
.C(n_111),
.Y(n_2144)
);

A2O1A1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_2076),
.A2(n_1382),
.B(n_1364),
.C(n_1435),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2081),
.Y(n_2146)
);

OAI222xp33_ASAP7_75t_L g2147 ( 
.A1(n_2078),
.A2(n_1434),
.B1(n_1405),
.B2(n_1382),
.C1(n_1378),
.C2(n_1364),
.Y(n_2147)
);

NAND4xp25_ASAP7_75t_L g2148 ( 
.A(n_2097),
.B(n_1378),
.C(n_1146),
.D(n_1121),
.Y(n_2148)
);

NAND3xp33_ASAP7_75t_L g2149 ( 
.A(n_2078),
.B(n_689),
.C(n_611),
.Y(n_2149)
);

NAND2xp33_ASAP7_75t_SL g2150 ( 
.A(n_2081),
.B(n_689),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2137),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2146),
.B(n_1901),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2107),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2142),
.B(n_711),
.Y(n_2154)
);

INVx1_ASAP7_75t_SL g2155 ( 
.A(n_2119),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_2111),
.B(n_711),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2141),
.Y(n_2157)
);

NOR2x1p5_ASAP7_75t_L g2158 ( 
.A(n_2135),
.B(n_711),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2138),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2115),
.B(n_1901),
.Y(n_2160)
);

OAI21xp33_ASAP7_75t_L g2161 ( 
.A1(n_2121),
.A2(n_1032),
.B(n_1232),
.Y(n_2161)
);

NAND4xp75_ASAP7_75t_L g2162 ( 
.A(n_2117),
.B(n_1086),
.C(n_1111),
.D(n_1097),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_2106),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2138),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_2105),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2122),
.A2(n_1145),
.B1(n_1175),
.B2(n_1453),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_SL g2167 ( 
.A1(n_2102),
.A2(n_1336),
.B1(n_1335),
.B2(n_1333),
.Y(n_2167)
);

NAND4xp25_ASAP7_75t_SL g2168 ( 
.A(n_2109),
.B(n_1087),
.C(n_1081),
.D(n_1070),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_2150),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2108),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2120),
.B(n_1901),
.Y(n_2171)
);

AOI221xp5_ASAP7_75t_L g2172 ( 
.A1(n_2103),
.A2(n_1034),
.B1(n_1042),
.B2(n_1057),
.C(n_1063),
.Y(n_2172)
);

AOI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_2112),
.A2(n_1034),
.B1(n_1042),
.B2(n_1057),
.C(n_1063),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2133),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2118),
.Y(n_2175)
);

NOR2x1_ASAP7_75t_SL g2176 ( 
.A(n_2136),
.B(n_1232),
.Y(n_2176)
);

NOR3xp33_ASAP7_75t_SL g2177 ( 
.A(n_2132),
.B(n_112),
.C(n_116),
.Y(n_2177)
);

AND2x4_ASAP7_75t_L g2178 ( 
.A(n_2145),
.B(n_1901),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2129),
.B(n_1145),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2110),
.A2(n_1067),
.B1(n_1335),
.B2(n_1333),
.Y(n_2180)
);

NOR3xp33_ASAP7_75t_SL g2181 ( 
.A(n_2116),
.B(n_118),
.C(n_119),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2134),
.Y(n_2182)
);

NOR3xp33_ASAP7_75t_SL g2183 ( 
.A(n_2131),
.B(n_120),
.C(n_122),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2124),
.A2(n_1175),
.B1(n_1042),
.B2(n_1057),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2113),
.A2(n_1175),
.B1(n_1034),
.B2(n_1063),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_L g2186 ( 
.A(n_2126),
.B(n_1232),
.Y(n_2186)
);

NOR2x1_ASAP7_75t_L g2187 ( 
.A(n_2123),
.B(n_1258),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2127),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_2159),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2164),
.B(n_2151),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2165),
.Y(n_2191)
);

OAI22xp5_ASAP7_75t_SL g2192 ( 
.A1(n_2157),
.A2(n_2101),
.B1(n_2149),
.B2(n_2130),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2188),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2155),
.B(n_2148),
.Y(n_2194)
);

NAND4xp25_ASAP7_75t_L g2195 ( 
.A(n_2153),
.B(n_2144),
.C(n_2104),
.D(n_2125),
.Y(n_2195)
);

NOR2x1p5_ASAP7_75t_L g2196 ( 
.A(n_2170),
.B(n_2114),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2163),
.A2(n_2139),
.B1(n_2128),
.B2(n_2140),
.Y(n_2197)
);

NOR4xp25_ASAP7_75t_L g2198 ( 
.A(n_2175),
.B(n_2143),
.C(n_2147),
.D(n_134),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_2158),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_SL g2200 ( 
.A(n_2169),
.B(n_125),
.C(n_129),
.Y(n_2200)
);

AOI22xp33_ASAP7_75t_SL g2201 ( 
.A1(n_2152),
.A2(n_1175),
.B1(n_1075),
.B2(n_1141),
.Y(n_2201)
);

NAND3xp33_ASAP7_75t_L g2202 ( 
.A(n_2163),
.B(n_1083),
.C(n_1075),
.Y(n_2202)
);

XNOR2xp5_ASAP7_75t_L g2203 ( 
.A(n_2183),
.B(n_135),
.Y(n_2203)
);

NOR2x1_ASAP7_75t_L g2204 ( 
.A(n_2174),
.B(n_1258),
.Y(n_2204)
);

NOR4xp25_ASAP7_75t_L g2205 ( 
.A(n_2154),
.B(n_137),
.C(n_144),
.D(n_148),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2176),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2160),
.B(n_149),
.Y(n_2207)
);

INVxp67_ASAP7_75t_L g2208 ( 
.A(n_2156),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2182),
.B(n_1141),
.C(n_1083),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2177),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2181),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2168),
.B(n_151),
.Y(n_2212)
);

AOI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2179),
.A2(n_1139),
.B(n_1075),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2185),
.A2(n_2186),
.B1(n_2184),
.B2(n_2178),
.Y(n_2214)
);

OAI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2173),
.A2(n_1149),
.B1(n_1084),
.B2(n_1088),
.C(n_1094),
.Y(n_2215)
);

NOR4xp25_ASAP7_75t_L g2216 ( 
.A(n_2161),
.B(n_153),
.C(n_154),
.D(n_156),
.Y(n_2216)
);

AO22x1_ASAP7_75t_L g2217 ( 
.A1(n_2180),
.A2(n_1336),
.B1(n_1335),
.B2(n_1333),
.Y(n_2217)
);

NOR3xp33_ASAP7_75t_L g2218 ( 
.A(n_2172),
.B(n_162),
.C(n_164),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_SL g2219 ( 
.A(n_2166),
.B(n_166),
.C(n_171),
.Y(n_2219)
);

OAI211xp5_ASAP7_75t_SL g2220 ( 
.A1(n_2187),
.A2(n_174),
.B(n_175),
.C(n_182),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2178),
.A2(n_1336),
.B1(n_1310),
.B2(n_1303),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_L g2222 ( 
.A(n_2167),
.B(n_1083),
.C(n_1084),
.Y(n_2222)
);

XNOR2xp5_ASAP7_75t_L g2223 ( 
.A(n_2191),
.B(n_2162),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2190),
.A2(n_2171),
.B(n_1139),
.Y(n_2224)
);

OAI22x1_ASAP7_75t_L g2225 ( 
.A1(n_2203),
.A2(n_1139),
.B1(n_185),
.B2(n_186),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2189),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_SL g2227 ( 
.A(n_2196),
.B(n_1258),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2207),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2193),
.B(n_184),
.Y(n_2229)
);

OAI22x1_ASAP7_75t_L g2230 ( 
.A1(n_2211),
.A2(n_189),
.B1(n_195),
.B2(n_200),
.Y(n_2230)
);

NAND3xp33_ASAP7_75t_L g2231 ( 
.A(n_2206),
.B(n_1141),
.C(n_1088),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2210),
.Y(n_2232)
);

NAND4xp25_ASAP7_75t_SL g2233 ( 
.A(n_2197),
.B(n_206),
.C(n_209),
.D(n_217),
.Y(n_2233)
);

HB1xp67_ASAP7_75t_L g2234 ( 
.A(n_2199),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2204),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2195),
.A2(n_1133),
.B1(n_1088),
.B2(n_1094),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2192),
.Y(n_2237)
);

XNOR2x1_ASAP7_75t_L g2238 ( 
.A(n_2194),
.B(n_218),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2200),
.B(n_1829),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2212),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_2205),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2208),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2217),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2214),
.Y(n_2244)
);

NOR2xp67_ASAP7_75t_L g2245 ( 
.A(n_2219),
.B(n_219),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2221),
.Y(n_2246)
);

NOR4xp25_ASAP7_75t_L g2247 ( 
.A(n_2215),
.B(n_228),
.C(n_229),
.D(n_232),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2201),
.B(n_234),
.Y(n_2248)
);

NAND3xp33_ASAP7_75t_SL g2249 ( 
.A(n_2226),
.B(n_2198),
.C(n_2213),
.Y(n_2249)
);

XOR2xp5_ASAP7_75t_L g2250 ( 
.A(n_2234),
.B(n_2242),
.Y(n_2250)
);

OAI221xp5_ASAP7_75t_L g2251 ( 
.A1(n_2237),
.A2(n_2216),
.B1(n_2218),
.B2(n_2220),
.C(n_2202),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2244),
.A2(n_2209),
.B(n_2222),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_2241),
.Y(n_2253)
);

NAND3x1_ASAP7_75t_L g2254 ( 
.A(n_2232),
.B(n_235),
.C(n_238),
.Y(n_2254)
);

AO211x2_ASAP7_75t_L g2255 ( 
.A1(n_2228),
.A2(n_240),
.B(n_241),
.C(n_242),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2229),
.B(n_1084),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_L g2257 ( 
.A(n_2240),
.B(n_1149),
.C(n_1096),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2238),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_L g2259 ( 
.A(n_2223),
.B(n_1149),
.C(n_1096),
.Y(n_2259)
);

OAI21xp5_ASAP7_75t_SL g2260 ( 
.A1(n_2248),
.A2(n_1094),
.B(n_1096),
.Y(n_2260)
);

XNOR2xp5_ASAP7_75t_L g2261 ( 
.A(n_2245),
.B(n_244),
.Y(n_2261)
);

AOI31xp33_ASAP7_75t_L g2262 ( 
.A1(n_2235),
.A2(n_249),
.A3(n_253),
.B(n_255),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2250),
.A2(n_2224),
.B(n_2227),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2253),
.A2(n_2243),
.B(n_2246),
.Y(n_2264)
);

XNOR2x1_ASAP7_75t_L g2265 ( 
.A(n_2261),
.B(n_2225),
.Y(n_2265)
);

INVx4_ASAP7_75t_L g2266 ( 
.A(n_2258),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2249),
.Y(n_2267)
);

OAI21x1_ASAP7_75t_SL g2268 ( 
.A1(n_2252),
.A2(n_2236),
.B(n_2247),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2254),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2255),
.A2(n_2239),
.B1(n_2233),
.B2(n_2231),
.Y(n_2270)
);

AOI221xp5_ASAP7_75t_L g2271 ( 
.A1(n_2264),
.A2(n_2251),
.B1(n_2256),
.B2(n_2260),
.C(n_2259),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2266),
.A2(n_2230),
.B1(n_2257),
.B2(n_2262),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2265),
.Y(n_2273)
);

OAI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2267),
.A2(n_1100),
.B1(n_1118),
.B2(n_1133),
.C(n_1273),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2269),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_SL g2276 ( 
.A1(n_2273),
.A2(n_2270),
.B1(n_2263),
.B2(n_2268),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2275),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2277),
.A2(n_2272),
.B1(n_2271),
.B2(n_2274),
.Y(n_2278)
);

OAI22x1_ASAP7_75t_L g2279 ( 
.A1(n_2276),
.A2(n_258),
.B1(n_259),
.B2(n_264),
.Y(n_2279)
);

OAI22x1_ASAP7_75t_L g2280 ( 
.A1(n_2278),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_2280)
);

OAI21x1_ASAP7_75t_L g2281 ( 
.A1(n_2280),
.A2(n_2279),
.B(n_278),
.Y(n_2281)
);

AOI222xp33_ASAP7_75t_L g2282 ( 
.A1(n_2281),
.A2(n_1100),
.B1(n_1118),
.B2(n_1133),
.C1(n_1273),
.C2(n_1310),
.Y(n_2282)
);

AOI22x1_ASAP7_75t_L g2283 ( 
.A1(n_2282),
.A2(n_1100),
.B1(n_1118),
.B2(n_1282),
.Y(n_2283)
);

OR2x6_ASAP7_75t_L g2284 ( 
.A(n_2283),
.B(n_1262),
.Y(n_2284)
);

AOI221xp5_ASAP7_75t_L g2285 ( 
.A1(n_2284),
.A2(n_1310),
.B1(n_1303),
.B2(n_1282),
.C(n_1273),
.Y(n_2285)
);

AOI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2285),
.A2(n_1303),
.B(n_1282),
.C(n_1268),
.Y(n_2286)
);


endmodule