module real_jpeg_25939_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_244;
wire n_167;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_1),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_1),
.A2(n_44),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_1),
.B(n_33),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_56),
.B1(n_57),
.B2(n_103),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_66),
.C(n_76),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_55),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_1),
.A2(n_63),
.B1(n_232),
.B2(n_239),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_26),
.B1(n_34),
.B2(n_37),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_26),
.B1(n_56),
.B2(n_57),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_26),
.B1(n_65),
.B2(n_66),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_34),
.B1(n_37),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_49),
.B1(n_65),
.B2(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_27),
.B1(n_44),
.B2(n_49),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_96)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_10),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_10),
.A2(n_34),
.B1(n_37),
.B2(n_117),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_117),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_117),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_34),
.B1(n_37),
.B2(n_80),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_29),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_13),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_42),
.B1(n_65),
.B2(n_66),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_34),
.B1(n_37),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_14),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_85)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_145),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_20),
.B(n_118),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_98),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_21),
.B(n_86),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_24),
.B(n_45),
.C(n_61),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_41),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_116),
.Y(n_115)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_36),
.C(n_37),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_31),
.A2(n_41),
.B(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_31),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_32),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_32),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_34),
.A2(n_38),
.B(n_102),
.C(n_104),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_34),
.B(n_103),
.CON(n_188),
.SN(n_188)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_37),
.A2(n_54),
.A3(n_57),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_40),
.B(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_58),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_48),
.B(n_55),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_50),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_50),
.A2(n_113),
.B1(n_138),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_50),
.A2(n_138),
.B1(n_155),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_51),
.B(n_59),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_51),
.A2(n_55),
.B1(n_179),
.B2(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_53),
.B(n_56),
.Y(n_189)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_57),
.B1(n_76),
.B2(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_57),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_74),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_63),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_63),
.A2(n_72),
.B(n_128),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_63),
.A2(n_89),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_63),
.A2(n_126),
.B1(n_229),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_73),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_70),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_64),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_66),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_65),
.B(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B(n_81),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_75),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_75),
.B(n_103),
.Y(n_237)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_96),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_123),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_95),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_82),
.A2(n_194),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_82),
.A2(n_95),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_82),
.A2(n_95),
.B1(n_193),
.B2(n_214),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_97),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_92),
.A2(n_108),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_98),
.A2(n_99),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.C(n_115),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_103),
.B(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_143),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_119)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_180),
.B(n_259),
.C(n_264),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_166),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_166),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_163),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_161),
.B2(n_162),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_149),
.B(n_162),
.C(n_163),
.Y(n_260)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_172),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_199),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_254),
.B(n_258),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_208),
.B(n_253),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_190),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_192),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_203),
.C(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_207),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_248),
.B(n_252),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_225),
.B(n_247),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_217),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_215),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_235),
.B(n_246),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_234),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_245),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);


endmodule