module fake_jpeg_31028_n_409 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_21;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_65),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_74),
.Y(n_131)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_9),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_84),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_7),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_19),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_106),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_36),
.B1(n_43),
.B2(n_38),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_18),
.B1(n_47),
.B2(n_45),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_32),
.B1(n_36),
.B2(n_60),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_50),
.B1(n_64),
.B2(n_46),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_61),
.B(n_38),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_54),
.B(n_42),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_22),
.B(n_42),
.C(n_32),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_18),
.B(n_78),
.C(n_37),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_119),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_34),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_36),
.C(n_43),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_75),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_146),
.Y(n_186)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_93),
.A2(n_67),
.B1(n_48),
.B2(n_58),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_150),
.Y(n_178)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_28),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_162),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_83),
.B1(n_51),
.B2(n_52),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_127),
.B(n_113),
.C(n_98),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_126),
.Y(n_180)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_44),
.B1(n_81),
.B2(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_27),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_114),
.B(n_57),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_158),
.C(n_142),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_149),
.B(n_135),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_150),
.B1(n_143),
.B2(n_145),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_196),
.B(n_206),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_155),
.B1(n_150),
.B2(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_117),
.B1(n_186),
.B2(n_98),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_168),
.B1(n_151),
.B2(n_167),
.Y(n_214)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_201),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_141),
.B(n_94),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_136),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_157),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_144),
.B1(n_91),
.B2(n_96),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_167),
.B1(n_175),
.B2(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_140),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_138),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_134),
.B(n_147),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_194),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_174),
.B1(n_176),
.B2(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_170),
.B1(n_174),
.B2(n_168),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_175),
.B(n_182),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_218),
.B1(n_223),
.B2(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_201),
.B1(n_189),
.B2(n_207),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_186),
.B1(n_100),
.B2(n_109),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_182),
.B1(n_173),
.B2(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_184),
.B1(n_153),
.B2(n_177),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_86),
.B1(n_97),
.B2(n_173),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_173),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_194),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_233),
.C(n_242),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_199),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_220),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_241),
.Y(n_249)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_225),
.B1(n_208),
.B2(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_198),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_183),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_221),
.C(n_212),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_214),
.C(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_223),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_218),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_215),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_245),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_258),
.B(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_205),
.C(n_86),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_209),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_236),
.B1(n_226),
.B2(n_177),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_215),
.B(n_211),
.C(n_194),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_236),
.B(n_231),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_271),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_230),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_278),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_236),
.B1(n_226),
.B2(n_217),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_276),
.B1(n_279),
.B2(n_284),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_169),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_177),
.B1(n_197),
.B2(n_192),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_166),
.B1(n_163),
.B2(n_139),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_259),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_266),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_187),
.C(n_169),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_286),
.C(n_254),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_249),
.B1(n_256),
.B2(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_187),
.C(n_169),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_113),
.B(n_87),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_288),
.Y(n_292)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_273),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_295),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_297),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_264),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_152),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_280),
.C(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_303),
.C(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_254),
.C(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_250),
.C(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_250),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_122),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_268),
.C(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_310),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_31),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_277),
.A2(n_266),
.B1(n_126),
.B2(n_100),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_281),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_312),
.A2(n_314),
.B1(n_132),
.B2(n_34),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_281),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_313),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_277),
.B1(n_156),
.B2(n_96),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_291),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_325),
.C(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_154),
.B(n_123),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_123),
.B(n_111),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_87),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_124),
.C(n_97),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_103),
.C(n_91),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_18),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_331),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_308),
.CI(n_289),
.CON(n_329),
.SN(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_159),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_159),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_78),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_62),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_103),
.C(n_132),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_72),
.C(n_55),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_316),
.A2(n_290),
.B(n_80),
.Y(n_335)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_340),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_322),
.A2(n_111),
.B(n_122),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_326),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_25),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_344),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_330),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_347),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_15),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_350),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_37),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_319),
.C(n_329),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.C(n_336),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_351),
.A2(n_320),
.B1(n_333),
.B2(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_341),
.B(n_315),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_358),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_318),
.C(n_325),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_37),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_334),
.B1(n_13),
.B2(n_14),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_348),
.A2(n_19),
.B1(n_35),
.B2(n_31),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_364),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_11),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_368),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_353),
.B(n_349),
.Y(n_368)
);

AOI322xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_337),
.A3(n_340),
.B1(n_342),
.B2(n_343),
.C1(n_352),
.C2(n_350),
.Y(n_371)
);

AOI211xp5_ASAP7_75t_L g382 ( 
.A1(n_371),
.A2(n_363),
.B(n_10),
.C(n_11),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_21),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_376),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_7),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_10),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_380),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_356),
.C(n_365),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_383),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_377),
.B(n_17),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_370),
.A2(n_373),
.B(n_375),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_385),
.A2(n_389),
.B(n_0),
.Y(n_394)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_369),
.A2(n_17),
.B(n_16),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_387),
.A2(n_1),
.B(n_2),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_13),
.Y(n_392)
);

NAND2x1_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_14),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_393),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_0),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_395),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_6),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_381),
.B(n_3),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_386),
.C(n_389),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_400),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_391),
.A2(n_1),
.B(n_4),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_401),
.A2(n_1),
.B(n_4),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_403),
.B(n_5),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_4),
.B(n_5),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_398),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_406),
.B(n_5),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_6),
.C(n_310),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_408),
.B(n_6),
.Y(n_409)
);


endmodule