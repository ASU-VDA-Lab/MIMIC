module fake_jpeg_10425_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_51),
.B1(n_56),
.B2(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_40),
.B1(n_47),
.B2(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_82),
.B1(n_83),
.B2(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_1),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_10),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_2),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_45),
.C(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_48),
.B1(n_44),
.B2(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_20),
.B1(n_36),
.B2(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_3),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_92),
.B(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.C(n_100),
.Y(n_102)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_99),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_91),
.B1(n_102),
.B2(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_93),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_82),
.C(n_74),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_83),
.C(n_68),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_109),
.C(n_79),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C(n_23),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_26),
.Y(n_117)
);


endmodule