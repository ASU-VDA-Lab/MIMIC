module fake_jpeg_26109_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_60),
.C(n_38),
.Y(n_80)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_55),
.Y(n_77)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_28),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_17),
.B1(n_16),
.B2(n_20),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_21),
.B1(n_23),
.B2(n_40),
.Y(n_84)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_68),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_69),
.Y(n_125)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_17),
.B1(n_39),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_84),
.B1(n_91),
.B2(n_96),
.Y(n_129)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_88),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_78),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_20),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_16),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_89),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_5),
.C(n_15),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_24),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_18),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_40),
.B1(n_17),
.B2(n_39),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_26),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_21),
.B1(n_43),
.B2(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_111),
.C(n_35),
.Y(n_146)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_38),
.C(n_44),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_95),
.Y(n_140)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_132),
.Y(n_145)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_140),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_92),
.B(n_84),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_159),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_26),
.B(n_101),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_163),
.CI(n_105),
.CON(n_182),
.SN(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_71),
.B1(n_62),
.B2(n_87),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_147),
.B1(n_162),
.B2(n_132),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_155),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_62),
.B1(n_93),
.B2(n_72),
.Y(n_147)
);

AO21x2_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_85),
.B(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_154),
.B1(n_146),
.B2(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_165),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_109),
.B1(n_111),
.B2(n_124),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_70),
.B1(n_82),
.B2(n_52),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_66),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_160),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_108),
.A2(n_103),
.B(n_31),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_73),
.B(n_1),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_52),
.B1(n_88),
.B2(n_41),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_41),
.C(n_35),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_35),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_181),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_162),
.B1(n_161),
.B2(n_73),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_195),
.B1(n_197),
.B2(n_151),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_127),
.B1(n_110),
.B2(n_114),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_210)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_121),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_194),
.B(n_137),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_113),
.B1(n_112),
.B2(n_107),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_107),
.B1(n_130),
.B2(n_41),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_130),
.B1(n_27),
.B2(n_29),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_86),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_193),
.Y(n_211)
);

AOI22x1_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_136),
.B1(n_159),
.B2(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_34),
.B1(n_33),
.B2(n_27),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_34),
.B1(n_33),
.B2(n_27),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_31),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_152),
.B(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_202),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_223),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_163),
.C(n_158),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_220),
.C(n_225),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_137),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_219),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_215),
.B(n_217),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_195),
.B1(n_178),
.B2(n_190),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_164),
.B(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_218),
.B1(n_197),
.B2(n_184),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_86),
.B(n_32),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_34),
.B1(n_33),
.B2(n_29),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_32),
.C(n_22),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_170),
.A2(n_32),
.B(n_22),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_177),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_167),
.B(n_32),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_29),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_182),
.A2(n_0),
.B(n_1),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_186),
.B1(n_185),
.B2(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_168),
.C(n_176),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_247),
.C(n_251),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_168),
.B1(n_175),
.B2(n_176),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_177),
.B1(n_182),
.B2(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_242),
.B1(n_233),
.B2(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_196),
.B1(n_179),
.B2(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_14),
.C(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_200),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_10),
.C(n_13),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_241),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_249),
.B(n_248),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_210),
.B1(n_213),
.B2(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_270),
.B1(n_243),
.B2(n_6),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_223),
.B1(n_203),
.B2(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_269),
.B1(n_243),
.B2(n_242),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_220),
.C(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_202),
.C(n_209),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_264),
.C(n_268),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_230),
.C(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_205),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_217),
.C(n_200),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_221),
.B1(n_227),
.B2(n_10),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_227),
.C(n_10),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_11),
.C(n_12),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_249),
.B(n_239),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_0),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_253),
.B(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_251),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_257),
.C(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_257),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_11),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_255),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_286),
.B(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_0),
.C(n_2),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_2),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_2),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_277),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_308),
.B(n_309),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_290),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_275),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_295),
.B1(n_288),
.B2(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_300),
.C(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_299),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_313),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_314),
.B(n_310),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_321),
.C(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_284),
.C(n_3),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_4),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_254),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_4),
.CI(n_284),
.CON(n_327),
.SN(n_327)
);


endmodule