module real_jpeg_2070_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_258, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_258;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_54),
.B1(n_61),
.B2(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_3),
.A2(n_49),
.B1(n_51),
.B2(n_113),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_61),
.B1(n_69),
.B2(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_35),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_27),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_61),
.C(n_76),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_49),
.B1(n_51),
.B2(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_55),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_65),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_4),
.B(n_74),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_35),
.B(n_162),
.Y(n_228)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_42),
.B1(n_61),
.B2(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_8),
.A2(n_61),
.B1(n_69),
.B2(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_79),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_9),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_39),
.B1(n_49),
.B2(n_51),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_9),
.A2(n_39),
.B1(n_61),
.B2(n_69),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_12),
.A2(n_37),
.B1(n_49),
.B2(n_51),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_37),
.B1(n_61),
.B2(n_69),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_49),
.B1(n_51),
.B2(n_68),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_114),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_21),
.B(n_84),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_57),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_40),
.C(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_25),
.A2(n_32),
.B1(n_36),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_25),
.A2(n_38),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_32),
.B1(n_112),
.B2(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_104),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_31),
.C(n_35),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_30),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_30),
.A2(n_33),
.B(n_103),
.C(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_35),
.B1(n_45),
.B2(n_47),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_33),
.B(n_47),
.C(n_51),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B(n_52),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_43),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_43),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_43),
.A2(n_48),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_43),
.A2(n_48),
.B1(n_147),
.B2(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_45),
.A2(n_49),
.B(n_161),
.C(n_163),
.Y(n_160)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_48),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_51),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_49),
.B(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_53),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_55),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_55),
.A2(n_108),
.B1(n_137),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_58),
.B(n_72),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_66),
.B(n_70),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_64),
.B(n_88),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_59),
.A2(n_70),
.B(n_88),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_59),
.A2(n_64),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_71),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_65),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_60),
.A2(n_87),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_60),
.A2(n_65),
.B1(n_104),
.B2(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_60),
.A2(n_65),
.B1(n_209),
.B2(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_69),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_61),
.B(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_64),
.A2(n_90),
.B(n_101),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_78),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_73),
.A2(n_93),
.B1(n_156),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_81),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_74),
.A2(n_82),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_74),
.A2(n_82),
.B1(n_195),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_158),
.Y(n_157)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_94),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_93),
.A2(n_123),
.B(n_158),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_95),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.C(n_111),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_96),
.A2(n_97),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_106),
.B(n_111),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_139),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_125),
.B2(n_126),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_138),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI321xp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_238),
.A3(n_249),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_184),
.B(n_237),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_165),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_144),
.B(n_165),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.C(n_159),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_145),
.B(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_154),
.B(n_159),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_164),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_177),
.B2(n_178),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_166),
.B(n_179),
.C(n_182),
.Y(n_250)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_168),
.B(n_172),
.C(n_176),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_232),
.B(n_236),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_222),
.B(n_231),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_203),
.B(n_221),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_215),
.B(n_220),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_210),
.B(n_214),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_213),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_241),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.C(n_248),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_243),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);


endmodule