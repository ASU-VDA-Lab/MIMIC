module fake_jpeg_1641_n_127 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_127);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_127;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_33),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_57),
.B1(n_58),
.B2(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_15),
.B(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_3),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_12),
.B(n_4),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_85),
.B1(n_92),
.B2(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_88),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_30),
.C(n_50),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_75),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_31),
.B1(n_38),
.B2(n_40),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_34),
.B(n_44),
.C(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_67),
.B1(n_68),
.B2(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_73),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_79),
.B(n_86),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_112),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_95),
.A3(n_62),
.B1(n_79),
.B2(n_75),
.C1(n_63),
.C2(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_99),
.C(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_105),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_104),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_110),
.B1(n_115),
.B2(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_119),
.B(n_107),
.Y(n_123)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.A3(n_108),
.B1(n_62),
.B2(n_64),
.C1(n_77),
.C2(n_61),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_108),
.Y(n_127)
);


endmodule