module real_aes_17273_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_0), .A2(n_69), .B1(n_327), .B2(n_346), .Y(n_345) );
INVxp33_ASAP7_75t_SL g451 ( .A(n_0), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_1), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_2), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_3), .A2(n_8), .B1(n_1275), .B2(n_1278), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_4), .A2(n_215), .B1(n_817), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_4), .A2(n_185), .B1(n_565), .B2(n_839), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_5), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_6), .A2(n_86), .B1(n_795), .B2(n_1188), .C(n_1189), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1213 ( .A1(n_6), .A2(n_133), .B1(n_334), .B2(n_510), .Y(n_1213) );
INVx1_ASAP7_75t_L g1487 ( .A(n_7), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_9), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_10), .A2(n_41), .B1(n_817), .B2(n_821), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_10), .A2(n_209), .B1(n_425), .B2(n_1574), .Y(n_1573) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_11), .A2(n_251), .B1(n_836), .B2(n_979), .C(n_981), .Y(n_978) );
INVx1_ASAP7_75t_L g1001 ( .A(n_11), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_12), .A2(n_193), .B1(n_621), .B2(n_706), .C(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g750 ( .A(n_12), .Y(n_750) );
INVx1_ASAP7_75t_L g294 ( .A(n_13), .Y(n_294) );
AND2x2_ASAP7_75t_L g407 ( .A(n_13), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g420 ( .A(n_13), .B(n_231), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_13), .B(n_304), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_14), .Y(n_1023) );
INVx1_ASAP7_75t_L g1224 ( .A(n_15), .Y(n_1224) );
OAI221xp5_ASAP7_75t_SL g1248 ( .A1(n_15), .A2(n_273), .B1(n_844), .B2(n_848), .C(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g769 ( .A(n_16), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_16), .A2(n_36), .B1(n_662), .B2(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g1271 ( .A(n_17), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_17), .B(n_110), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_17), .B(n_1277), .Y(n_1279) );
INVx1_ASAP7_75t_L g813 ( .A(n_18), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_18), .A2(n_155), .B1(n_844), .B2(n_847), .C(n_852), .Y(n_843) );
INVx1_ASAP7_75t_L g1127 ( .A(n_19), .Y(n_1127) );
OAI222xp33_ASAP7_75t_L g1175 ( .A1(n_20), .A2(n_148), .B1(n_848), .B2(n_1176), .C1(n_1177), .C2(n_1181), .Y(n_1175) );
INVx1_ASAP7_75t_L g1204 ( .A(n_20), .Y(n_1204) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_21), .A2(n_239), .B1(n_1275), .B2(n_1278), .Y(n_1304) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_22), .Y(n_1031) );
OAI21xp5_ASAP7_75t_L g1578 ( .A1(n_23), .A2(n_672), .B(n_1579), .Y(n_1578) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_24), .A2(n_268), .B1(n_296), .B2(n_1056), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_24), .A2(n_268), .B1(n_1087), .B2(n_1090), .Y(n_1086) );
INVx1_ASAP7_75t_L g1577 ( .A(n_25), .Y(n_1577) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_26), .A2(n_76), .B1(n_349), .B2(n_350), .C(n_352), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_26), .A2(n_29), .B1(n_474), .B2(n_475), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_27), .Y(n_536) );
INVx1_ASAP7_75t_L g1564 ( .A(n_28), .Y(n_1564) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_29), .A2(n_132), .B1(n_318), .B2(n_327), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_30), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_31), .A2(n_169), .B1(n_320), .B2(n_623), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_31), .A2(n_135), .B1(n_1157), .B2(n_1160), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_32), .Y(n_883) );
INVx1_ASAP7_75t_L g1193 ( .A(n_33), .Y(n_1193) );
AOI22xp5_ASAP7_75t_L g1293 ( .A1(n_34), .A2(n_272), .B1(n_1268), .B2(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g366 ( .A(n_35), .Y(n_366) );
OA222x2_ASAP7_75t_L g413 ( .A1(n_35), .A2(n_165), .B1(n_276), .B2(n_414), .C1(n_421), .C2(n_429), .Y(n_413) );
INVx1_ASAP7_75t_L g782 ( .A(n_36), .Y(n_782) );
INVx1_ASAP7_75t_L g777 ( .A(n_37), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_37), .A2(n_176), .B1(n_795), .B2(n_798), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_38), .A2(n_205), .B1(n_334), .B2(n_336), .C(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g468 ( .A(n_38), .Y(n_468) );
INVx1_ASAP7_75t_L g1133 ( .A(n_39), .Y(n_1133) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_40), .A2(n_349), .B(n_690), .C(n_694), .Y(n_689) );
INVx1_ASAP7_75t_L g742 ( .A(n_40), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g1568 ( .A1(n_41), .A2(n_123), .B1(n_649), .B2(n_856), .C(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g801 ( .A(n_42), .Y(n_801) );
INVx1_ASAP7_75t_L g985 ( .A(n_43), .Y(n_985) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_44), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_44), .A2(n_86), .B1(n_334), .B2(n_510), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_45), .A2(n_77), .B1(n_388), .B2(n_998), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_45), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_46), .A2(n_250), .B1(n_1275), .B2(n_1278), .Y(n_1297) );
AO22x1_ASAP7_75t_L g1301 ( .A1(n_47), .A2(n_58), .B1(n_1268), .B2(n_1283), .Y(n_1301) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_48), .A2(n_167), .B1(n_684), .B2(n_685), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_48), .A2(n_82), .B1(n_890), .B2(n_892), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g1512 ( .A1(n_49), .A2(n_1513), .B(n_1516), .C(n_1517), .Y(n_1512) );
INVx1_ASAP7_75t_L g1530 ( .A(n_49), .Y(n_1530) );
INVx1_ASAP7_75t_L g1180 ( .A(n_50), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_50), .A2(n_245), .B1(n_708), .B2(n_924), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_51), .A2(n_267), .B1(n_1090), .B2(n_1522), .Y(n_1521) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_51), .A2(n_126), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
AOI22xp33_ASAP7_75t_SL g1561 ( .A1(n_52), .A2(n_114), .B1(n_320), .B2(n_391), .Y(n_1561) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_52), .A2(n_81), .B1(n_442), .B2(n_650), .C(n_1154), .Y(n_1572) );
INVx1_ASAP7_75t_L g326 ( .A(n_53), .Y(n_326) );
INVx1_ASAP7_75t_L g332 ( .A(n_53), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_54), .A2(n_257), .B1(n_368), .B2(n_684), .C(n_685), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_54), .A2(n_127), .B1(n_485), .B2(n_489), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_55), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_56), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_57), .A2(n_108), .B1(n_529), .B2(n_687), .C(n_758), .Y(n_757) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_57), .Y(n_789) );
INVx1_ASAP7_75t_L g287 ( .A(n_59), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_60), .A2(n_221), .B1(n_336), .B2(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_60), .A2(n_159), .B1(n_659), .B2(n_662), .C(n_663), .Y(n_658) );
INVx2_ASAP7_75t_L g344 ( .A(n_61), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_62), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_63), .A2(n_245), .B1(n_425), .B2(n_858), .Y(n_1190) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_63), .A2(n_151), .B1(n_924), .B2(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1494 ( .A(n_64), .Y(n_1494) );
INVx1_ASAP7_75t_L g932 ( .A(n_65), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_65), .A2(n_227), .B1(n_425), .B2(n_474), .Y(n_954) );
INVxp67_ASAP7_75t_SL g968 ( .A(n_66), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g1009 ( .A1(n_66), .A2(n_368), .B(n_1010), .C(n_1011), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_67), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_68), .A2(n_181), .B1(n_1268), .B2(n_1283), .Y(n_1298) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_69), .Y(n_472) );
INVx1_ASAP7_75t_L g895 ( .A(n_70), .Y(n_895) );
INVx1_ASAP7_75t_L g1118 ( .A(n_71), .Y(n_1118) );
AO221x2_ASAP7_75t_L g1340 ( .A1(n_71), .A2(n_217), .B1(n_1275), .B2(n_1278), .C(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1491 ( .A(n_72), .Y(n_1491) );
INVx1_ASAP7_75t_L g1553 ( .A(n_73), .Y(n_1553) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_74), .A2(n_116), .B1(n_619), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_74), .A2(n_137), .B1(n_652), .B2(n_653), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_75), .A2(n_254), .B1(n_524), .B2(n_526), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_75), .A2(n_213), .B1(n_652), .B2(n_653), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_76), .A2(n_205), .B1(n_442), .B2(n_444), .C(n_447), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g1238 ( .A1(n_77), .A2(n_99), .B1(n_650), .B2(n_1162), .C(n_1239), .Y(n_1238) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_78), .Y(n_595) );
INVx1_ASAP7_75t_L g970 ( .A(n_79), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_80), .A2(n_262), .B1(n_1060), .B2(n_1063), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1107 ( .A1(n_80), .A2(n_262), .B1(n_1108), .B2(n_1110), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_81), .A2(n_230), .B1(n_1138), .B2(n_1558), .Y(n_1557) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_82), .A2(n_166), .B1(n_518), .B2(n_940), .C(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g387 ( .A(n_83), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_83), .B(n_400), .Y(n_399) );
OAI222xp33_ASAP7_75t_L g901 ( .A1(n_84), .A2(n_128), .B1(n_247), .B2(n_531), .C1(n_695), .C2(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g916 ( .A(n_84), .Y(n_916) );
INVx1_ASAP7_75t_L g780 ( .A(n_85), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_85), .A2(n_233), .B1(n_425), .B2(n_474), .Y(n_796) );
XOR2x2_ASAP7_75t_L g678 ( .A(n_87), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_88), .A2(n_94), .B1(n_1136), .B2(n_1138), .Y(n_1135) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_88), .A2(n_125), .B1(n_648), .B2(n_650), .C(n_1154), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_89), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_90), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_91), .A2(n_240), .B1(n_659), .B2(n_973), .Y(n_972) );
AOI21xp33_ASAP7_75t_L g1004 ( .A1(n_91), .A2(n_341), .B(n_1005), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_92), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_93), .A2(n_127), .B1(n_700), .B2(n_703), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_93), .A2(n_400), .B(n_716), .C(n_724), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_94), .A2(n_207), .B1(n_662), .B2(n_663), .C(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g390 ( .A(n_95), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_95), .A2(n_187), .B1(n_485), .B2(n_489), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_96), .A2(n_120), .B1(n_391), .B2(n_510), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_96), .A2(n_280), .B1(n_444), .B2(n_836), .C(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g887 ( .A(n_97), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_97), .A2(n_146), .B1(n_621), .B2(n_907), .C(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g698 ( .A(n_98), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g1232 ( .A1(n_99), .A2(n_162), .B1(n_629), .B2(n_1233), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_100), .Y(n_289) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_100), .B(n_287), .Y(n_1269) );
INVx1_ASAP7_75t_L g712 ( .A(n_101), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_102), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_103), .A2(n_156), .B1(n_350), .B2(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_103), .A2(n_104), .B1(n_475), .B2(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g548 ( .A(n_104), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g1166 ( .A1(n_105), .A2(n_672), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1227 ( .A(n_106), .Y(n_1227) );
XOR2x2_ASAP7_75t_L g802 ( .A(n_107), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g800 ( .A(n_108), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_109), .A2(n_496), .B1(n_497), .B2(n_587), .Y(n_495) );
INVx1_ASAP7_75t_L g587 ( .A(n_109), .Y(n_587) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_110), .B(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1277 ( .A(n_110), .Y(n_1277) );
INVx1_ASAP7_75t_L g710 ( .A(n_111), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g1124 ( .A(n_112), .B(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_113), .A2(n_137), .B1(n_617), .B2(n_619), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_113), .A2(n_116), .B1(n_644), .B2(n_648), .C(n_650), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_114), .A2(n_230), .B1(n_475), .B2(n_858), .Y(n_1570) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_115), .Y(n_601) );
INVx2_ASAP7_75t_L g343 ( .A(n_117), .Y(n_343) );
INVx1_ASAP7_75t_L g355 ( .A(n_117), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_117), .B(n_344), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_118), .Y(n_927) );
INVx1_ASAP7_75t_L g896 ( .A(n_119), .Y(n_896) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_119), .A2(n_153), .B1(n_684), .B2(n_685), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_120), .A2(n_270), .B1(n_839), .B2(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_121), .A2(n_147), .B1(n_501), .B2(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_122), .A2(n_211), .B1(n_1268), .B2(n_1283), .Y(n_1287) );
XNOR2xp5_ASAP7_75t_L g1480 ( .A(n_122), .B(n_1481), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1542 ( .A1(n_122), .A2(n_1543), .B1(n_1548), .B2(n_1580), .Y(n_1542) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_123), .A2(n_209), .B1(n_817), .B2(n_821), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_124), .A2(n_185), .B1(n_817), .B2(n_819), .Y(n_816) );
AOI21xp33_ASAP7_75t_L g855 ( .A1(n_124), .A2(n_836), .B(n_856), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_125), .A2(n_135), .B1(n_388), .B2(n_1138), .C(n_1143), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_126), .A2(n_179), .B1(n_1087), .B2(n_1510), .Y(n_1509) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_128), .A2(n_153), .B1(n_480), .B2(n_890), .C(n_892), .Y(n_889) );
INVx1_ASAP7_75t_L g866 ( .A(n_129), .Y(n_866) );
INVx1_ASAP7_75t_L g783 ( .A(n_130), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_130), .A2(n_189), .B1(n_652), .B2(n_653), .Y(n_799) );
INVx1_ASAP7_75t_L g1518 ( .A(n_131), .Y(n_1518) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_132), .Y(n_448) );
INVxp67_ASAP7_75t_SL g1183 ( .A(n_133), .Y(n_1183) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_134), .Y(n_805) );
OAI211xp5_ASAP7_75t_SL g1184 ( .A1(n_136), .A2(n_1185), .B(n_1186), .C(n_1191), .Y(n_1184) );
INVx1_ASAP7_75t_L g1207 ( .A(n_136), .Y(n_1207) );
INVx1_ASAP7_75t_L g1497 ( .A(n_138), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_139), .A2(n_145), .B1(n_529), .B2(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_139), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_140), .A2(n_687), .B1(n_930), .B2(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g949 ( .A(n_140), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_141), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g1554 ( .A(n_142), .Y(n_1554) );
INVx1_ASAP7_75t_L g982 ( .A(n_143), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_143), .A2(n_220), .B1(n_924), .B2(n_1007), .Y(n_1006) );
AO22x1_ASAP7_75t_L g1302 ( .A1(n_144), .A2(n_235), .B1(n_1275), .B2(n_1278), .Y(n_1302) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_145), .Y(n_720) );
INVx1_ASAP7_75t_L g873 ( .A(n_146), .Y(n_873) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_147), .A2(n_833), .B(n_834), .C(n_840), .Y(n_832) );
INVx1_ASAP7_75t_L g1203 ( .A(n_148), .Y(n_1203) );
INVx1_ASAP7_75t_L g1492 ( .A(n_149), .Y(n_1492) );
BUFx3_ASAP7_75t_L g323 ( .A(n_150), .Y(n_323) );
INVx1_ASAP7_75t_L g1179 ( .A(n_151), .Y(n_1179) );
INVx1_ASAP7_75t_L g1498 ( .A(n_152), .Y(n_1498) );
XNOR2x1_ASAP7_75t_L g1171 ( .A(n_154), .B(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g811 ( .A(n_155), .Y(n_811) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_156), .A2(n_243), .B1(n_565), .B2(n_567), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_157), .A2(n_159), .B1(n_524), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_157), .A2(n_221), .B1(n_652), .B2(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g692 ( .A(n_158), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g671 ( .A1(n_160), .A2(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g987 ( .A(n_161), .Y(n_987) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_162), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_163), .A2(n_174), .B1(n_1275), .B2(n_1278), .Y(n_1284) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_164), .Y(n_301) );
INVx1_ASAP7_75t_L g392 ( .A(n_165), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g946 ( .A1(n_166), .A2(n_947), .B(n_948), .C(n_951), .Y(n_946) );
INVx1_ASAP7_75t_L g950 ( .A(n_167), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_168), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g1155 ( .A1(n_169), .A2(n_271), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
INVx1_ASAP7_75t_L g1576 ( .A(n_170), .Y(n_1576) );
INVx1_ASAP7_75t_L g1520 ( .A(n_171), .Y(n_1520) );
OAI211xp5_ASAP7_75t_SL g1525 ( .A1(n_171), .A2(n_1072), .B(n_1526), .C(n_1527), .Y(n_1525) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_172), .A2(n_807), .B(n_1195), .Y(n_1194) );
OAI222xp33_ASAP7_75t_L g1234 ( .A1(n_173), .A2(n_212), .B1(n_246), .B2(n_594), .C1(n_597), .C2(n_672), .Y(n_1234) );
OAI211xp5_ASAP7_75t_L g1236 ( .A1(n_173), .A2(n_1185), .B(n_1237), .C(n_1243), .Y(n_1236) );
INVx1_ASAP7_75t_L g969 ( .A(n_175), .Y(n_969) );
INVx1_ASAP7_75t_L g768 ( .A(n_176), .Y(n_768) );
INVx1_ASAP7_75t_L g1563 ( .A(n_177), .Y(n_1563) );
INVx1_ASAP7_75t_L g1081 ( .A(n_178), .Y(n_1081) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_178), .A2(n_1094), .B(n_1096), .C(n_1098), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1536 ( .A1(n_179), .A2(n_267), .B1(n_296), .B2(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g514 ( .A(n_180), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_180), .A2(n_429), .B1(n_570), .B2(n_578), .C(n_579), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_182), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_183), .A2(n_253), .B1(n_1268), .B2(n_1283), .Y(n_1305) );
INVx1_ASAP7_75t_L g936 ( .A(n_184), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_184), .A2(n_190), .B1(n_474), .B2(n_568), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_186), .A2(n_256), .B1(n_826), .B2(n_830), .Y(n_825) );
INVx1_ASAP7_75t_L g841 ( .A(n_186), .Y(n_841) );
INVx1_ASAP7_75t_L g363 ( .A(n_187), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_188), .Y(n_1024) );
INVx1_ASAP7_75t_L g774 ( .A(n_189), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_190), .A2(n_227), .B1(n_351), .B2(n_924), .C(n_925), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_191), .A2(n_248), .B1(n_1268), .B2(n_1283), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_192), .Y(n_504) );
INVx1_ASAP7_75t_L g734 ( .A(n_193), .Y(n_734) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
INVx1_ASAP7_75t_L g760 ( .A(n_195), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_195), .A2(n_197), .B1(n_485), .B2(n_489), .Y(n_792) );
OAI211xp5_ASAP7_75t_L g1069 ( .A1(n_196), .A2(n_1070), .B(n_1072), .C(n_1075), .Y(n_1069) );
INVx1_ASAP7_75t_L g1106 ( .A(n_196), .Y(n_1106) );
INVx1_ASAP7_75t_L g763 ( .A(n_197), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_198), .Y(n_604) );
INVx1_ASAP7_75t_L g696 ( .A(n_199), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_200), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g1039 ( .A(n_201), .Y(n_1039) );
INVx1_ASAP7_75t_L g1495 ( .A(n_202), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_203), .Y(n_879) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_204), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_204), .A2(n_687), .B1(n_913), .B2(n_914), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_206), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1144 ( .A1(n_207), .A2(n_271), .B1(n_1136), .B2(n_1145), .Y(n_1144) );
AO22x1_ASAP7_75t_L g1267 ( .A1(n_208), .A2(n_238), .B1(n_1268), .B2(n_1272), .Y(n_1267) );
CKINVDCx16_ASAP7_75t_R g1342 ( .A(n_210), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_213), .A2(n_252), .B1(n_522), .B2(n_819), .Y(n_1231) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_214), .A2(n_991), .B(n_992), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_214), .A2(n_236), .B1(n_529), .B2(n_687), .Y(n_993) );
INVx1_ASAP7_75t_L g853 ( .A(n_215), .Y(n_853) );
OAI211xp5_ASAP7_75t_L g761 ( .A1(n_216), .A2(n_368), .B(n_394), .C(n_762), .Y(n_761) );
INVxp33_ASAP7_75t_SL g791 ( .A(n_216), .Y(n_791) );
INVx1_ASAP7_75t_L g682 ( .A(n_218), .Y(n_682) );
INVx1_ASAP7_75t_L g965 ( .A(n_219), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_220), .A2(n_264), .B1(n_425), .B2(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g1149 ( .A(n_222), .Y(n_1149) );
INVx1_ASAP7_75t_L g1131 ( .A(n_223), .Y(n_1131) );
INVx1_ASAP7_75t_L g499 ( .A(n_224), .Y(n_499) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_225), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_225), .A2(n_368), .B1(n_529), .B2(n_532), .C(n_542), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_226), .Y(n_875) );
INVx1_ASAP7_75t_L g1014 ( .A(n_228), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_229), .A2(n_265), .B1(n_1275), .B2(n_1278), .Y(n_1292) );
BUFx3_ASAP7_75t_L g304 ( .A(n_231), .Y(n_304) );
INVx1_ASAP7_75t_L g408 ( .A(n_231), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_232), .Y(n_1026) );
INVx1_ASAP7_75t_L g771 ( .A(n_233), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g1344 ( .A(n_234), .Y(n_1344) );
INVx1_ASAP7_75t_L g493 ( .A(n_235), .Y(n_493) );
INVxp33_ASAP7_75t_L g989 ( .A(n_236), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_237), .A2(n_341), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g562 ( .A(n_237), .Y(n_562) );
INVx1_ASAP7_75t_L g996 ( .A(n_240), .Y(n_996) );
XNOR2xp5_ASAP7_75t_L g1549 ( .A(n_241), .B(n_1550), .Y(n_1549) );
XOR2xp5_ASAP7_75t_L g590 ( .A(n_242), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g541 ( .A(n_243), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_244), .Y(n_511) );
INVx1_ASAP7_75t_L g898 ( .A(n_247), .Y(n_898) );
INVx2_ASAP7_75t_L g398 ( .A(n_249), .Y(n_398) );
INVx1_ASAP7_75t_L g405 ( .A(n_249), .Y(n_405) );
INVx1_ASAP7_75t_L g418 ( .A(n_249), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_251), .A2(n_264), .B1(n_352), .B2(n_629), .C(n_998), .Y(n_997) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_252), .A2(n_254), .B1(n_1154), .B2(n_1254), .C(n_1255), .Y(n_1253) );
INVx1_ASAP7_75t_L g1151 ( .A(n_255), .Y(n_1151) );
INVx1_ASAP7_75t_L g842 ( .A(n_256), .Y(n_842) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_257), .Y(n_723) );
INVx1_ASAP7_75t_L g919 ( .A(n_258), .Y(n_919) );
INVx1_ASAP7_75t_L g1226 ( .A(n_259), .Y(n_1226) );
AO22x1_ASAP7_75t_L g1274 ( .A1(n_260), .A2(n_274), .B1(n_1275), .B2(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g938 ( .A(n_261), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_263), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_266), .B(n_583), .Y(n_582) );
OAI21xp33_ASAP7_75t_SL g755 ( .A1(n_269), .A2(n_400), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_269), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_270), .A2(n_280), .B1(n_391), .B2(n_510), .Y(n_824) );
INVx1_ASAP7_75t_L g1223 ( .A(n_273), .Y(n_1223) );
XNOR2xp5_ASAP7_75t_L g1218 ( .A(n_274), .B(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1485 ( .A(n_275), .Y(n_1485) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_276), .A2(n_279), .B1(n_380), .B2(n_381), .C(n_386), .Y(n_379) );
INVx1_ASAP7_75t_L g513 ( .A(n_277), .Y(n_513) );
INVx1_ASAP7_75t_L g1192 ( .A(n_278), .Y(n_1192) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_279), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_305), .B(n_1260), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g1541 ( .A(n_284), .B(n_293), .Y(n_1541) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_286), .B(n_289), .Y(n_1547) );
INVx1_ASAP7_75t_L g1583 ( .A(n_286), .Y(n_1583) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_289), .B(n_1583), .Y(n_1585) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_293), .B(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g458 ( .A(n_294), .B(n_304), .Y(n_458) );
AND2x4_ASAP7_75t_L g664 ( .A(n_294), .B(n_303), .Y(n_664) );
AND2x4_ASAP7_75t_SL g1540 ( .A(n_295), .B(n_1541), .Y(n_1540) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_302), .Y(n_296) );
BUFx4f_ASAP7_75t_L g874 ( .A(n_297), .Y(n_874) );
INVxp67_ASAP7_75t_L g886 ( .A(n_297), .Y(n_886) );
INVx1_ASAP7_75t_L g984 ( .A(n_297), .Y(n_984) );
OR2x6_ASAP7_75t_L g1062 ( .A(n_297), .B(n_1058), .Y(n_1062) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx4f_ASAP7_75t_L g450 ( .A(n_298), .Y(n_450) );
INVx3_ASAP7_75t_L g748 ( .A(n_298), .Y(n_748) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g410 ( .A(n_300), .Y(n_410) );
INVx2_ASAP7_75t_L g428 ( .A(n_300), .Y(n_428) );
NAND2x1_ASAP7_75t_L g431 ( .A(n_300), .B(n_301), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_300), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g446 ( .A(n_300), .B(n_301), .Y(n_446) );
INVx1_ASAP7_75t_L g492 ( .A(n_300), .Y(n_492) );
INVx1_ASAP7_75t_L g411 ( .A(n_301), .Y(n_411) );
AND2x2_ASAP7_75t_L g427 ( .A(n_301), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g439 ( .A(n_301), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_301), .B(n_428), .Y(n_456) );
OR2x2_ASAP7_75t_L g467 ( .A(n_301), .B(n_410), .Y(n_467) );
BUFx2_ASAP7_75t_L g488 ( .A(n_301), .Y(n_488) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g1074 ( .A(n_303), .Y(n_1074) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_304), .Y(n_1068) );
AND2x4_ASAP7_75t_L g1080 ( .A(n_304), .B(n_491), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_1119), .B2(n_1120), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_861), .Y(n_307) );
XOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_588), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
XNOR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_495), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_493), .B(n_494), .Y(n_312) );
AND3x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_412), .C(n_440), .Y(n_313) );
AOI31xp33_ASAP7_75t_L g494 ( .A1(n_314), .A2(n_412), .A3(n_440), .B(n_493), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_395), .B(n_399), .Y(n_314) );
NAND3xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_357), .C(n_373), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_333), .B1(n_345), .B2(n_348), .Y(n_316) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g618 ( .A(n_320), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_320), .B(n_942), .Y(n_941) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_320), .Y(n_1007) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
INVx8_ASAP7_75t_L g389 ( .A(n_321), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_321), .B(n_361), .Y(n_394) );
AND2x2_ASAP7_75t_L g701 ( .A(n_321), .B(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g1558 ( .A(n_321), .Y(n_1558) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
AND2x4_ASAP7_75t_L g339 ( .A(n_322), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_323), .Y(n_329) );
AND2x4_ASAP7_75t_L g335 ( .A(n_323), .B(n_331), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_323), .B(n_332), .Y(n_385) );
OR2x2_ASAP7_75t_L g540 ( .A(n_323), .B(n_325), .Y(n_540) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g340 ( .A(n_326), .Y(n_340) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx5_ASAP7_75t_L g527 ( .A(n_328), .Y(n_527) );
AND2x4_ASAP7_75t_L g586 ( .A(n_328), .B(n_377), .Y(n_586) );
BUFx3_ASAP7_75t_L g621 ( .A(n_328), .Y(n_621) );
BUFx3_ASAP7_75t_L g623 ( .A(n_328), .Y(n_623) );
BUFx12f_ASAP7_75t_L g924 ( .A(n_328), .Y(n_924) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_329), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_329), .Y(n_1102) );
INVx1_ASAP7_75t_L g365 ( .A(n_330), .Y(n_365) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g371 ( .A(n_332), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_334), .A2(n_504), .B1(n_510), .B2(n_511), .Y(n_509) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g349 ( .A(n_335), .Y(n_349) );
BUFx2_ASAP7_75t_L g391 ( .A(n_335), .Y(n_391) );
BUFx2_ASAP7_75t_L g619 ( .A(n_335), .Y(n_619) );
BUFx2_ASAP7_75t_L g632 ( .A(n_335), .Y(n_632) );
AND2x2_ASAP7_75t_L g704 ( .A(n_335), .B(n_702), .Y(n_704) );
INVx2_ASAP7_75t_L g999 ( .A(n_335), .Y(n_999) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_335), .B(n_356), .Y(n_1097) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_337), .A2(n_1033), .B1(n_1491), .B2(n_1497), .Y(n_1503) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g347 ( .A(n_338), .Y(n_347) );
INVx3_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx5_ASAP7_75t_L g818 ( .A(n_338), .Y(n_818) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx8_ASAP7_75t_L g524 ( .A(n_339), .Y(n_524) );
INVx2_ASAP7_75t_L g531 ( .A(n_339), .Y(n_531) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_339), .Y(n_708) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_342), .B(n_461), .Y(n_1021) );
NAND2xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
AND3x4_ASAP7_75t_L g614 ( .A(n_343), .B(n_552), .C(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g693 ( .A(n_343), .B(n_615), .Y(n_693) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_343), .Y(n_1115) );
INVx3_ASAP7_75t_L g356 ( .A(n_344), .Y(n_356) );
BUFx3_ASAP7_75t_L g615 ( .A(n_344), .Y(n_615) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g908 ( .A(n_351), .Y(n_908) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_353), .A2(n_533), .B1(n_536), .B2(n_537), .C(n_541), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_353), .A2(n_535), .B1(n_710), .B2(n_711), .C(n_712), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g776 ( .A1(n_353), .A2(n_711), .B1(n_777), .B2(n_778), .C(n_780), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_353), .A2(n_535), .B1(n_711), .B2(n_875), .C(n_883), .Y(n_913) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_353), .A2(n_369), .B1(n_539), .B2(n_931), .C(n_932), .Y(n_930) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x6_ASAP7_75t_L g823 ( .A(n_354), .B(n_397), .Y(n_823) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND3x1_ASAP7_75t_L g626 ( .A(n_355), .B(n_356), .C(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g361 ( .A(n_356), .B(n_362), .Y(n_361) );
OR2x4_ASAP7_75t_L g1089 ( .A(n_356), .B(n_540), .Y(n_1089) );
INVx1_ASAP7_75t_L g1092 ( .A(n_356), .Y(n_1092) );
OR2x6_ASAP7_75t_L g1112 ( .A(n_356), .B(n_384), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_363), .B1(n_364), .B2(n_366), .C(n_367), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_358), .A2(n_364), .B1(n_513), .B2(n_514), .Y(n_512) );
INVx4_ASAP7_75t_L g684 ( .A(n_358), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_358), .A2(n_364), .B1(n_763), .B2(n_764), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_358), .A2(n_364), .B1(n_969), .B2(n_987), .Y(n_1011) );
AND2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_359), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g812 ( .A(n_359), .B(n_607), .Y(n_812) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_359), .B(n_607), .Y(n_1132) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g364 ( .A(n_361), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g372 ( .A(n_361), .Y(n_372) );
AND2x4_ASAP7_75t_L g607 ( .A(n_361), .B(n_417), .Y(n_607) );
INVx2_ASAP7_75t_L g685 ( .A(n_364), .Y(n_685) );
INVx1_ASAP7_75t_L g611 ( .A(n_365), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g905 ( .A(n_367), .B(n_906), .C(n_912), .Y(n_905) );
NOR3xp33_ASAP7_75t_L g922 ( .A(n_367), .B(n_923), .C(n_929), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_368), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g1003 ( .A(n_369), .Y(n_1003) );
INVx1_ASAP7_75t_L g1095 ( .A(n_369), .Y(n_1095) );
INVx1_ASAP7_75t_L g1515 ( .A(n_369), .Y(n_1515) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_370), .Y(n_520) );
BUFx3_ASAP7_75t_L g535 ( .A(n_370), .Y(n_535) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_371), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_379), .B1(n_392), .B2(n_393), .Y(n_373) );
INVxp67_ASAP7_75t_L g508 ( .A(n_374), .Y(n_508) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g903 ( .A(n_376), .Y(n_903) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g530 ( .A(n_377), .Y(n_530) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g600 ( .A(n_378), .B(n_461), .Y(n_600) );
INVx1_ASAP7_75t_L g702 ( .A(n_378), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_380), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_933) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g1506 ( .A(n_383), .Y(n_1506) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_384), .Y(n_1033) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g547 ( .A(n_385), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_390), .B2(n_391), .Y(n_386) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx8_ASAP7_75t_L g510 ( .A(n_389), .Y(n_510) );
INVx2_ASAP7_75t_L g629 ( .A(n_389), .Y(n_629) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_393), .A2(n_682), .B(n_683), .C(n_686), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_393), .A2(n_895), .B1(n_901), .B2(n_903), .C(n_904), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_393), .A2(n_903), .B1(n_938), .B2(n_939), .C(n_943), .Y(n_937) );
INVx2_ASAP7_75t_L g1010 ( .A(n_393), .Y(n_1010) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g501 ( .A(n_394), .B(n_502), .Y(n_501) );
OR2x6_ASAP7_75t_L g594 ( .A(n_394), .B(n_502), .Y(n_594) );
INVx1_ASAP7_75t_L g670 ( .A(n_395), .Y(n_670) );
INVx2_ASAP7_75t_L g714 ( .A(n_395), .Y(n_714) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_396), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g1013 ( .A(n_396), .Y(n_1013) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g478 ( .A(n_397), .B(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_398), .B(n_420), .Y(n_483) );
INVx2_ASAP7_75t_L g552 ( .A(n_398), .Y(n_552) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g498 ( .A1(n_401), .A2(n_435), .B1(n_499), .B2(n_500), .C1(n_504), .C2(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_401), .B(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_401), .B(n_942), .Y(n_945) );
AOI211x1_ASAP7_75t_L g964 ( .A1(n_401), .A2(n_965), .B(n_966), .C(n_990), .Y(n_964) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_406), .Y(n_401) );
AND2x4_ASAP7_75t_L g435 ( .A(n_402), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g489 ( .A(n_403), .B(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g502 ( .A(n_403), .Y(n_502) );
OR2x2_ASAP7_75t_L g892 ( .A(n_403), .B(n_490), .Y(n_892) );
INVx1_ASAP7_75t_L g1084 ( .A(n_403), .Y(n_1084) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_406), .Y(n_637) );
INVx1_ASAP7_75t_L g1245 ( .A(n_406), .Y(n_1245) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_407), .B(n_418), .Y(n_424) );
AND2x2_ASAP7_75t_L g436 ( .A(n_407), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g640 ( .A(n_407), .B(n_437), .Y(n_640) );
AND2x4_ASAP7_75t_L g642 ( .A(n_407), .B(n_568), .Y(n_642) );
AND2x4_ASAP7_75t_SL g657 ( .A(n_407), .B(n_445), .Y(n_657) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_408), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_409), .B(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
INVx3_ASAP7_75t_L g566 ( .A(n_409), .Y(n_566) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_432), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_416), .B(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g597 ( .A(n_416), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g718 ( .A(n_417), .Y(n_718) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g627 ( .A(n_418), .Y(n_627) );
INVx1_ASAP7_75t_L g719 ( .A(n_419), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_420), .B(n_491), .Y(n_490) );
AND2x6_ASAP7_75t_L g654 ( .A(n_420), .B(n_445), .Y(n_654) );
AND2x2_ASAP7_75t_L g668 ( .A(n_420), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g851 ( .A(n_420), .Y(n_851) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g503 ( .A(n_422), .Y(n_503) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_422), .A2(n_682), .B1(n_717), .B2(n_720), .C1(n_721), .C2(n_723), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g790 ( .A1(n_422), .A2(n_791), .B(n_792), .Y(n_790) );
AOI222xp33_ASAP7_75t_L g893 ( .A1(n_422), .A2(n_717), .B1(n_721), .B2(n_894), .C1(n_895), .C2(n_896), .Y(n_893) );
AOI222xp33_ASAP7_75t_L g967 ( .A1(n_422), .A2(n_580), .B1(n_581), .B2(n_968), .C1(n_969), .C2(n_970), .Y(n_967) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
AOI332xp33_ASAP7_75t_L g948 ( .A1(n_423), .A2(n_425), .A3(n_718), .B1(n_719), .B2(n_721), .B3(n_938), .C1(n_949), .C2(n_950), .Y(n_948) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g429 ( .A(n_424), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g722 ( .A(n_424), .B(n_430), .Y(n_722) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_427), .Y(n_568) );
BUFx3_ASAP7_75t_L g653 ( .A(n_427), .Y(n_653) );
BUFx3_ASAP7_75t_L g882 ( .A(n_430), .Y(n_882) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_430), .Y(n_1049) );
BUFx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_435), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_435), .B(n_789), .Y(n_788) );
NAND2xp33_ASAP7_75t_SL g915 ( .A(n_435), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g947 ( .A(n_435), .Y(n_947) );
INVx1_ASAP7_75t_L g991 ( .A(n_435), .Y(n_991) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_437), .Y(n_795) );
INVx2_ASAP7_75t_L g1165 ( .A(n_437), .Y(n_1165) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g443 ( .A(n_438), .Y(n_443) );
BUFx3_ASAP7_75t_L g649 ( .A(n_438), .Y(n_649) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_438), .B(n_1058), .Y(n_1057) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_457), .B(n_462), .C(n_484), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g661 ( .A(n_443), .Y(n_661) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g662 ( .A(n_445), .Y(n_662) );
BUFx3_ASAP7_75t_L g798 ( .A(n_445), .Y(n_798) );
INVx1_ASAP7_75t_L g980 ( .A(n_445), .Y(n_980) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_445), .B(n_1074), .Y(n_1073) );
BUFx3_ASAP7_75t_L g1154 ( .A(n_445), .Y(n_1154) );
BUFx6f_ASAP7_75t_L g1569 ( .A(n_445), .Y(n_1569) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g647 ( .A(n_446), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_451), .B2(n_452), .Y(n_447) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_450), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_452), .A2(n_1023), .B1(n_1037), .B2(n_1043), .Y(n_1042) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_452), .A2(n_1250), .B1(n_1251), .B2(n_1252), .C(n_1253), .Y(n_1249) );
INVx6_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g738 ( .A(n_454), .Y(n_738) );
INVx2_ASAP7_75t_SL g749 ( .A(n_454), .Y(n_749) );
INVx4_ASAP7_75t_L g986 ( .A(n_454), .Y(n_986) );
INVx1_ASAP7_75t_L g1053 ( .A(n_454), .Y(n_1053) );
INVx8_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_455), .B(n_1068), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_457), .Y(n_578) );
AOI332xp33_ASAP7_75t_L g793 ( .A1(n_457), .A2(n_557), .A3(n_717), .B1(n_794), .B2(n_796), .B3(n_797), .C1(n_799), .C2(n_800), .Y(n_793) );
AOI322xp5_ASAP7_75t_L g971 ( .A1(n_457), .A2(n_721), .A3(n_972), .B1(n_975), .B2(n_977), .C1(n_978), .C2(n_987), .Y(n_971) );
INVx2_ASAP7_75t_L g1050 ( .A(n_457), .Y(n_1050) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx4_ASAP7_75t_L g650 ( .A(n_458), .Y(n_650) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_458), .B(n_461), .Y(n_745) );
INVx1_ASAP7_75t_SL g837 ( .A(n_458), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_458), .B(n_459), .Y(n_955) );
INVx4_ASAP7_75t_L g1189 ( .A(n_458), .Y(n_1189) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_461), .Y(n_1117) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_476), .B(n_480), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_468), .B1(n_469), .B2(n_472), .C(n_473), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g1177 ( .A1(n_464), .A2(n_664), .B1(n_1178), .B2(n_1179), .C(n_1180), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g1493 ( .A1(n_464), .A2(n_1048), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_466), .A2(n_563), .B1(n_927), .B2(n_934), .C(n_954), .Y(n_953) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g561 ( .A(n_467), .Y(n_561) );
BUFx2_ASAP7_75t_L g573 ( .A(n_467), .Y(n_573) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g743 ( .A(n_470), .Y(n_743) );
INVx2_ASAP7_75t_L g854 ( .A(n_470), .Y(n_854) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g480 ( .A(n_471), .B(n_481), .Y(n_480) );
BUFx4f_ASAP7_75t_L g563 ( .A(n_471), .Y(n_563) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_471), .Y(n_574) );
BUFx4f_ASAP7_75t_L g733 ( .A(n_471), .Y(n_733) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_471), .Y(n_958) );
BUFx4f_ASAP7_75t_L g1178 ( .A(n_471), .Y(n_1178) );
INVx3_ASAP7_75t_L g577 ( .A(n_474), .Y(n_577) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_474), .Y(n_858) );
INVx1_ASAP7_75t_L g977 ( .A(n_476), .Y(n_977) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g558 ( .A(n_478), .Y(n_558) );
INVx2_ASAP7_75t_L g730 ( .A(n_478), .Y(n_730) );
INVx2_ASAP7_75t_L g871 ( .A(n_478), .Y(n_871) );
INVx1_ASAP7_75t_L g1041 ( .A(n_478), .Y(n_1041) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_480), .A2(n_555), .B(n_559), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_480), .Y(n_727) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2x2_ASAP7_75t_L g485 ( .A(n_482), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g580 ( .A(n_485), .Y(n_580) );
INVx2_ASAP7_75t_SL g891 ( .A(n_485), .Y(n_891) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g669 ( .A(n_488), .Y(n_669) );
INVx1_ASAP7_75t_L g850 ( .A(n_488), .Y(n_850) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_488), .B(n_1068), .Y(n_1076) );
AND2x4_ASAP7_75t_L g1529 ( .A(n_488), .B(n_1068), .Y(n_1529) );
INVx2_ASAP7_75t_SL g581 ( .A(n_489), .Y(n_581) );
AND2x4_ASAP7_75t_L g672 ( .A(n_489), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g807 ( .A(n_489), .B(n_673), .Y(n_807) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_506), .C(n_553), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_528), .B(n_549), .Y(n_506) );
OAI211xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_512), .C(n_515), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_511), .A2(n_513), .B1(n_580), .B2(n_581), .Y(n_579) );
OAI211xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_521), .C(n_525), .Y(n_515) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_516), .A2(n_536), .B1(n_571), .B2(n_574), .C(n_575), .Y(n_570) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g902 ( .A(n_519), .Y(n_902) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g673 ( .A(n_520), .B(n_600), .Y(n_673) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_520), .Y(n_767) );
INVx4_ASAP7_75t_L g779 ( .A(n_520), .Y(n_779) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_520), .A2(n_693), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_925) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_520), .Y(n_1038) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_523), .A2(n_775), .B1(n_877), .B2(n_888), .Y(n_914) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g543 ( .A(n_524), .Y(n_543) );
AND2x4_ASAP7_75t_L g677 ( .A(n_524), .B(n_676), .Y(n_677) );
INVx3_ASAP7_75t_L g691 ( .A(n_524), .Y(n_691) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g819 ( .A(n_527), .Y(n_819) );
INVx2_ASAP7_75t_R g821 ( .A(n_527), .Y(n_821) );
OR2x6_ASAP7_75t_SL g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx3_ASAP7_75t_L g911 ( .A(n_531), .Y(n_911) );
BUFx2_ASAP7_75t_L g1137 ( .A(n_531), .Y(n_1137) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_533), .A2(n_695), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_535), .A2(n_693), .B1(n_879), .B2(n_881), .C(n_910), .Y(n_909) );
BUFx6f_ASAP7_75t_L g1502 ( .A(n_535), .Y(n_1502) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx4f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g695 ( .A(n_540), .Y(n_695) );
BUFx3_ASAP7_75t_L g711 ( .A(n_540), .Y(n_711) );
INVx2_ASAP7_75t_L g773 ( .A(n_540), .Y(n_773) );
OR2x4_ASAP7_75t_L g1109 ( .A(n_540), .B(n_1092), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_548), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_544), .A2(n_560), .B1(n_562), .B2(n_563), .C(n_564), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g995 ( .A1(n_545), .A2(n_940), .B1(n_985), .B2(n_996), .C(n_997), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_545), .A2(n_1026), .B1(n_1027), .B2(n_1029), .Y(n_1025) );
CKINVDCx8_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g697 ( .A(n_546), .Y(n_697) );
INVx3_ASAP7_75t_L g775 ( .A(n_546), .Y(n_775) );
INVx3_ASAP7_75t_L g935 ( .A(n_546), .Y(n_935) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g599 ( .A(n_547), .Y(n_599) );
INVx1_ASAP7_75t_L g859 ( .A(n_549), .Y(n_859) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g1257 ( .A(n_550), .Y(n_1257) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_551), .Y(n_944) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI31xp33_ASAP7_75t_SL g756 ( .A1(n_552), .A2(n_757), .A3(n_761), .B(n_765), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_569), .C(n_582), .Y(n_553) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
OAI33xp33_ASAP7_75t_L g1483 ( .A1(n_558), .A2(n_955), .A3(n_1484), .B1(n_1490), .B2(n_1493), .B3(n_1496), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_560), .A2(n_563), .B1(n_1026), .B2(n_1031), .Y(n_1044) );
INVx1_ASAP7_75t_L g1047 ( .A(n_560), .Y(n_1047) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g741 ( .A(n_561), .Y(n_741) );
INVx2_ASAP7_75t_L g957 ( .A(n_561), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1490 ( .A1(n_563), .A2(n_571), .B1(n_1491), .B2(n_1492), .Y(n_1490) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g652 ( .A(n_566), .Y(n_652) );
INVx2_ASAP7_75t_L g976 ( .A(n_566), .Y(n_976) );
INVx2_ASAP7_75t_L g1156 ( .A(n_566), .Y(n_1156) );
INVx1_ASAP7_75t_L g1160 ( .A(n_566), .Y(n_1160) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_568), .Y(n_839) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g732 ( .A(n_572), .Y(n_732) );
INVx4_ASAP7_75t_L g878 ( .A(n_572), .Y(n_878) );
INVx4_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g1574 ( .A(n_577), .Y(n_1574) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g687 ( .A(n_586), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_751), .B1(n_752), .B2(n_860), .Y(n_588) );
INVx1_ASAP7_75t_L g860 ( .A(n_589), .Y(n_860) );
XNOR2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_678), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_633), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_596), .B2(n_601), .C(n_602), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_593), .A2(n_596), .B1(n_1127), .B2(n_1128), .C(n_1129), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_593), .B(n_1207), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1552 ( .A1(n_593), .A2(n_596), .B1(n_1553), .B2(n_1554), .C(n_1555), .Y(n_1552) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_595), .A2(n_642), .B1(n_643), .B2(n_651), .C(n_654), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g804 ( .A1(n_596), .A2(n_805), .B(n_806), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_596), .B(n_1200), .Y(n_1199) );
INVx8_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g785 ( .A(n_599), .Y(n_785) );
INVx1_ASAP7_75t_L g676 ( .A(n_600), .Y(n_676) );
INVx1_ASAP7_75t_L g829 ( .A(n_600), .Y(n_829) );
NAND3xp33_ASAP7_75t_SL g602 ( .A(n_603), .B(n_612), .C(n_630), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_603) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_604), .A2(n_608), .B1(n_656), .B2(n_658), .C1(n_665), .C2(n_666), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_605), .A2(n_1203), .B1(n_1204), .B2(n_1205), .Y(n_1202) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g609 ( .A(n_607), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g631 ( .A(n_607), .B(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_SL g1205 ( .A(n_607), .B(n_610), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_609), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_609), .A2(n_1131), .B1(n_1132), .B2(n_1133), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_609), .A2(n_1132), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1562 ( .A1(n_609), .A2(n_812), .B1(n_1563), .B2(n_1564), .Y(n_1562) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI33xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .A3(n_620), .B1(n_622), .B2(n_624), .B3(n_628), .Y(n_612) );
INVx1_ASAP7_75t_L g1143 ( .A(n_613), .Y(n_1143) );
AOI33xp33_ASAP7_75t_L g1228 ( .A1(n_613), .A2(n_1035), .A3(n_1229), .B1(n_1230), .B2(n_1231), .B3(n_1232), .Y(n_1228) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI33xp33_ASAP7_75t_L g814 ( .A1(n_614), .A2(n_815), .A3(n_816), .B1(n_820), .B2(n_822), .B3(n_824), .Y(n_814) );
AOI33xp33_ASAP7_75t_L g1208 ( .A1(n_614), .A2(n_1209), .A3(n_1210), .B1(n_1211), .B2(n_1213), .B3(n_1214), .Y(n_1208) );
AOI33xp33_ASAP7_75t_L g1556 ( .A1(n_614), .A2(n_822), .A3(n_1557), .B1(n_1559), .B2(n_1560), .B3(n_1561), .Y(n_1556) );
INVx3_ASAP7_75t_L g1101 ( .A(n_615), .Y(n_1101) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_625), .Y(n_1140) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_625), .Y(n_1214) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g1035 ( .A(n_626), .Y(n_1035) );
AND2x4_ASAP7_75t_L g675 ( .A(n_629), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_629), .B(n_676), .Y(n_1196) );
NAND3xp33_ASAP7_75t_SL g1129 ( .A(n_630), .B(n_1130), .C(n_1134), .Y(n_1129) );
INVx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_631), .B(n_809), .C(n_825), .Y(n_808) );
INVx3_ASAP7_75t_L g1215 ( .A(n_631), .Y(n_1215) );
NOR3xp33_ASAP7_75t_L g1220 ( .A(n_631), .B(n_1221), .C(n_1234), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_632), .Y(n_1233) );
AOI21xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_670), .B(n_671), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_641), .C(n_655), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_636), .A2(n_638), .B1(n_675), .B2(n_677), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_637), .A2(n_640), .B1(n_841), .B2(n_842), .Y(n_840) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_637), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_637), .A2(n_640), .B1(n_1192), .B2(n_1193), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_637), .A2(n_640), .B1(n_1576), .B2(n_1577), .Y(n_1575) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_639), .A2(n_1149), .B1(n_1150), .B2(n_1151), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g1247 ( .A(n_640), .Y(n_1247) );
INVx2_ASAP7_75t_SL g833 ( .A(n_642), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_642), .A2(n_654), .B1(n_1127), .B2(n_1153), .C(n_1155), .Y(n_1152) );
INVx3_ASAP7_75t_L g1185 ( .A(n_642), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1571 ( .A1(n_642), .A2(n_654), .B1(n_1553), .B2(n_1572), .C(n_1573), .Y(n_1571) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g974 ( .A(n_647), .Y(n_974) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g1157 ( .A(n_653), .Y(n_1157) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_654), .A2(n_835), .B(n_838), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g1186 ( .A1(n_654), .A2(n_1187), .B(n_1190), .Y(n_1186) );
AOI21xp5_ASAP7_75t_SL g1237 ( .A1(n_654), .A2(n_1238), .B(n_1242), .Y(n_1237) );
AOI222xp33_ASAP7_75t_L g1158 ( .A1(n_656), .A2(n_666), .B1(n_1131), .B2(n_1133), .C1(n_1159), .C2(n_1161), .Y(n_1158) );
AOI222xp33_ASAP7_75t_L g1567 ( .A1(n_656), .A2(n_668), .B1(n_1563), .B2(n_1564), .C1(n_1568), .C2(n_1570), .Y(n_1567) );
BUFx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g846 ( .A(n_657), .Y(n_846) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g836 ( .A(n_660), .Y(n_836) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g856 ( .A(n_664), .Y(n_856) );
INVx2_ASAP7_75t_L g1255 ( .A(n_664), .Y(n_1255) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_SL g1174 ( .A1(n_670), .A2(n_1175), .B(n_1184), .C(n_1194), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_675), .A2(n_677), .B1(n_1149), .B2(n_1151), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_675), .A2(n_677), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
INVx2_ASAP7_75t_L g830 ( .A(n_677), .Y(n_830) );
AOI211x1_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_713), .B(n_715), .C(n_726), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_688), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_699), .C(n_705), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_693), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_691), .A2(n_693), .B1(n_767), .B2(n_768), .C(n_769), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_691), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g1212 ( .A(n_691), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_692), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_695), .A2(n_1037), .B1(n_1038), .B2(n_1039), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_696), .A2(n_712), .B1(n_736), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_698), .A2(n_747), .B1(n_749), .B2(n_750), .Y(n_746) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_701), .A2(n_704), .B1(n_759), .B2(n_760), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_701), .A2(n_704), .B1(n_965), .B2(n_970), .Y(n_1008) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g928 ( .A(n_708), .Y(n_928) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_708), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g1028 ( .A(n_708), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_708), .B(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_710), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g899 ( .A1(n_714), .A2(n_900), .B(n_905), .C(n_915), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g1146 ( .A1(n_714), .A2(n_1147), .B(n_1166), .Y(n_1146) );
AOI21xp33_ASAP7_75t_L g988 ( .A1(n_717), .A2(n_727), .B(n_989), .Y(n_988) );
AND2x4_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_721), .A2(n_727), .B(n_764), .Y(n_787) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR3x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .C(n_729), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g951 ( .A(n_727), .B(n_952), .C(n_960), .Y(n_951) );
OAI33xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .A3(n_735), .B1(n_739), .B2(n_744), .B3(n_746), .Y(n_729) );
INVx1_ASAP7_75t_L g1071 ( .A(n_733), .Y(n_1071) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g1043 ( .A(n_737), .Y(n_1043) );
INVx2_ASAP7_75t_L g1250 ( .A(n_737), .Y(n_1250) );
INVx2_ASAP7_75t_SL g1486 ( .A(n_737), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_740), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_880) );
INVx4_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI33xp33_ASAP7_75t_L g870 ( .A1(n_744), .A2(n_871), .A3(n_872), .B1(n_876), .B2(n_880), .B3(n_884), .Y(n_870) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_749), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_749), .A2(n_885), .B1(n_887), .B2(n_888), .Y(n_884) );
INVx1_ASAP7_75t_L g1489 ( .A(n_749), .Y(n_1489) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_802), .Y(n_752) );
XOR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_801), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_786), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_770), .B1(n_776), .B2(n_781), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_774), .B2(n_775), .Y(n_770) );
INVx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_SL g827 ( .A(n_773), .Y(n_827) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND4xp25_ASAP7_75t_SL g786 ( .A(n_787), .B(n_788), .C(n_790), .D(n_793), .Y(n_786) );
BUFx3_ASAP7_75t_L g1254 ( .A(n_795), .Y(n_1254) );
NAND3xp33_ASAP7_75t_SL g803 ( .A(n_804), .B(n_808), .C(n_831), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
INVx2_ASAP7_75t_L g1505 ( .A(n_817), .Y(n_1505) );
INVx8_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
OR2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g1501 ( .A1(n_827), .A2(n_1485), .B1(n_1494), .B2(n_1502), .Y(n_1501) );
OAI22xp33_ASAP7_75t_L g1507 ( .A1(n_827), .A2(n_902), .B1(n_1487), .B2(n_1495), .Y(n_1507) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_829), .B(n_911), .Y(n_1197) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_843), .B(n_859), .Y(n_831) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g1176 ( .A(n_845), .Y(n_1176) );
INVx4_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
OAI211xp5_ASAP7_75t_SL g852 ( .A1(n_853), .A2(n_854), .B(n_855), .C(n_857), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_854), .A2(n_877), .B1(n_878), .B2(n_879), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g1565 ( .A1(n_859), .A2(n_1566), .B(n_1578), .Y(n_1565) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_961), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
XNOR2x1_ASAP7_75t_L g864 ( .A(n_865), .B(n_917), .Y(n_864) );
XNOR2x1_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
NOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_899), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_893), .C(n_897), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_889), .Y(n_869) );
OAI22xp5_ASAP7_75t_SL g952 ( .A1(n_871), .A2(n_953), .B1(n_955), .B2(n_956), .Y(n_952) );
BUFx2_ASAP7_75t_L g1526 ( .A(n_882), .Y(n_1526) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_910), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g940 ( .A(n_911), .Y(n_940) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
XNOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
OR2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_946), .Y(n_920) );
A2O1A1Ixp33_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_937), .B(n_944), .C(n_945), .Y(n_921) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_924), .Y(n_1145) );
OAI221xp5_ASAP7_75t_L g956 ( .A1(n_926), .A2(n_931), .B1(n_957), .B2(n_958), .C(n_959), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_963), .B1(n_1015), .B2(n_1016), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
XOR2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_1014), .Y(n_963) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_971), .C(n_988), .Y(n_966) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx2_ASAP7_75t_L g1241 ( .A(n_974), .Y(n_1241) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g1188 ( .A(n_980), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_983), .B1(n_985), .B2(n_986), .Y(n_981) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI31xp33_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .A3(n_1009), .B(n_1012), .Y(n_992) );
NAND3xp33_ASAP7_75t_L g994 ( .A(n_995), .B(n_1000), .C(n_1008), .Y(n_994) );
INVx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1138 ( .A(n_999), .Y(n_1138) );
OAI211xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B(n_1004), .C(n_1006), .Y(n_1000) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
XOR2x2_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1118), .Y(n_1016) );
AND3x1_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1054), .C(n_1085), .Y(n_1017) );
NOR2xp33_ASAP7_75t_SL g1018 ( .A(n_1019), .B(n_1040), .Y(n_1018) );
OAI33xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1022), .A3(n_1025), .B1(n_1030), .B2(n_1034), .B3(n_1036), .Y(n_1019) );
BUFx8_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
BUFx4f_ASAP7_75t_L g1500 ( .A(n_1021), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_1024), .A2(n_1039), .B1(n_1046), .B2(n_1048), .Y(n_1045) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_1029), .A2(n_1032), .B1(n_1043), .B2(n_1052), .Y(n_1051) );
OAI33xp33_ASAP7_75t_L g1499 ( .A1(n_1034), .A2(n_1500), .A3(n_1501), .B1(n_1503), .B2(n_1504), .B3(n_1507), .Y(n_1499) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
OAI33xp33_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .A3(n_1044), .B1(n_1045), .B2(n_1050), .B3(n_1051), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_1043), .A2(n_1052), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx5_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_1052), .A2(n_1486), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI31xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1059), .A3(n_1069), .B(n_1082), .Y(n_1054) );
INVx4_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
CKINVDCx16_ASAP7_75t_R g1537 ( .A(n_1057), .Y(n_1537) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
BUFx6f_ASAP7_75t_L g1533 ( .A(n_1062), .Y(n_1533) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1535 ( .A(n_1067), .Y(n_1535) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx3_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_1076), .A2(n_1077), .B1(n_1078), .B2(n_1081), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_1077), .A2(n_1099), .B1(n_1103), .B2(n_1106), .Y(n_1098) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1531 ( .A(n_1080), .Y(n_1531) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
BUFx2_ASAP7_75t_SL g1538 ( .A(n_1083), .Y(n_1538) );
OAI31xp33_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1093), .A3(n_1107), .B(n_1113), .Y(n_1085) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVxp67_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
CKINVDCx8_ASAP7_75t_R g1096 ( .A(n_1097), .Y(n_1096) );
CKINVDCx8_ASAP7_75t_R g1516 ( .A(n_1097), .Y(n_1516) );
BUFx3_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1101), .B(n_1105), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1519 ( .A(n_1101), .B(n_1102), .Y(n_1519) );
BUFx6f_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_1104), .A2(n_1518), .B1(n_1519), .B2(n_1520), .Y(n_1517) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1511 ( .A(n_1109), .Y(n_1511) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
BUFx3_ASAP7_75t_L g1522 ( .A(n_1112), .Y(n_1522) );
AND2x2_ASAP7_75t_SL g1113 ( .A(n_1114), .B(n_1116), .Y(n_1113) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_1114), .B(n_1116), .Y(n_1523) );
INVx1_ASAP7_75t_SL g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1122), .B1(n_1168), .B2(n_1169), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
NAND2xp67_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1146), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1139), .B1(n_1142), .B2(n_1144), .Y(n_1134) );
INVx2_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
NAND3xp33_ASAP7_75t_SL g1147 ( .A(n_1148), .B(n_1152), .C(n_1158), .Y(n_1147) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1216), .B1(n_1258), .B2(n_1259), .Y(n_1169) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1170), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NOR2x1p5_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1198), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_1192), .A2(n_1193), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_1196), .A2(n_1197), .B1(n_1576), .B2(n_1577), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1201), .Y(n_1198) );
AND4x1_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1206), .C(n_1208), .D(n_1215), .Y(n_1201) );
NAND3xp33_ASAP7_75t_L g1555 ( .A(n_1215), .B(n_1556), .C(n_1562), .Y(n_1555) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1216), .Y(n_1259) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1235), .Y(n_1219) );
NAND3xp33_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1225), .C(n_1228), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_1226), .A2(n_1227), .B1(n_1244), .B2(n_1246), .Y(n_1243) );
OAI21xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1248), .B(n_1256), .Y(n_1235) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
OAI221xp5_ASAP7_75t_SL g1260 ( .A1(n_1261), .A2(n_1474), .B1(n_1478), .B2(n_1539), .C(n_1542), .Y(n_1260) );
NOR3xp33_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1411), .C(n_1450), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1346), .C(n_1378), .Y(n_1262) );
AOI211xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1289), .B(n_1306), .C(n_1325), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1264), .B(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1264), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1280), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1265), .B(n_1286), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g1398 ( .A(n_1265), .B(n_1384), .C(n_1399), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1265), .B(n_1315), .Y(n_1404) );
OR2x2_ASAP7_75t_L g1422 ( .A(n_1265), .B(n_1286), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1265), .B(n_1379), .Y(n_1436) );
CKINVDCx6p67_ASAP7_75t_R g1265 ( .A(n_1266), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1266), .B(n_1286), .Y(n_1313) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1266), .B(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1266), .B(n_1315), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1266), .B(n_1286), .Y(n_1415) );
CKINVDCx5p33_ASAP7_75t_R g1438 ( .A(n_1266), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1266), .B(n_1340), .Y(n_1443) );
OR2x6_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1274), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1267), .B(n_1274), .Y(n_1427) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1268), .Y(n_1343) );
AND2x6_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1269), .B(n_1273), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1275 ( .A(n_1269), .B(n_1276), .Y(n_1275) );
AND2x6_ASAP7_75t_L g1278 ( .A(n_1269), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1269), .B(n_1273), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1269), .B(n_1273), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1271), .B(n_1277), .Y(n_1276) );
OAI21xp5_ASAP7_75t_L g1582 ( .A1(n_1273), .A2(n_1583), .B(n_1584), .Y(n_1582) );
AOI21xp33_ASAP7_75t_L g1363 ( .A1(n_1280), .A2(n_1339), .B(n_1364), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1280), .B(n_1310), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1285), .Y(n_1280) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1281), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1281), .B(n_1286), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1377 ( .A(n_1281), .B(n_1286), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1281), .B(n_1296), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1284), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1345 ( .A(n_1283), .Y(n_1345) );
HB1xp67_ASAP7_75t_L g1477 ( .A(n_1283), .Y(n_1477) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_1286), .A2(n_1307), .B1(n_1311), .B2(n_1317), .C(n_1323), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1286), .B(n_1316), .Y(n_1338) );
A2O1A1Ixp33_ASAP7_75t_L g1346 ( .A1(n_1286), .A2(n_1347), .B(n_1361), .C(n_1362), .Y(n_1346) );
INVx3_ASAP7_75t_L g1407 ( .A(n_1286), .Y(n_1407) );
O2A1O1Ixp33_ASAP7_75t_L g1451 ( .A1(n_1286), .A2(n_1452), .B(n_1453), .C(n_1454), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1286), .B(n_1296), .Y(n_1465) );
AND2x4_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
AOI21xp5_ASAP7_75t_L g1454 ( .A1(n_1290), .A2(n_1377), .B(n_1455), .Y(n_1454) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1295), .Y(n_1290) );
INVx2_ASAP7_75t_L g1308 ( .A(n_1291), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1291), .B(n_1320), .Y(n_1324) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1291), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1291), .B(n_1299), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1291), .B(n_1366), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1299), .Y(n_1295) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1296), .Y(n_1310) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1296), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1296), .B(n_1352), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1296), .B(n_1370), .Y(n_1369) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1296), .B(n_1420), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1296), .B(n_1320), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1299), .B(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1299), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1299), .B(n_1441), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1299), .B(n_1359), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1303), .Y(n_1299) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1300), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1300), .B(n_1322), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1300), .B(n_1352), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1302), .Y(n_1300) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1303), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1303), .B(n_1308), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1351 ( .A(n_1303), .B(n_1352), .Y(n_1351) );
AND3x1_ASAP7_75t_L g1355 ( .A(n_1303), .B(n_1308), .C(n_1321), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1303), .B(n_1352), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1303), .B(n_1321), .Y(n_1384) );
OAI21xp33_ASAP7_75t_L g1416 ( .A1(n_1303), .A2(n_1417), .B(n_1418), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1305), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1308), .B(n_1318), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1308), .B(n_1320), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1308), .B(n_1366), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1308), .B(n_1321), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1308), .B(n_1310), .Y(n_1441) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1310), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1310), .B(n_1366), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1310), .B(n_1373), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1310), .B(n_1370), .Y(n_1392) );
O2A1O1Ixp33_ASAP7_75t_L g1401 ( .A1(n_1310), .A2(n_1334), .B(n_1402), .C(n_1403), .Y(n_1401) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1310), .B(n_1351), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1310), .B(n_1315), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1314), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
OAI21xp33_ASAP7_75t_L g1395 ( .A1(n_1313), .A2(n_1396), .B(n_1398), .Y(n_1395) );
OAI222xp33_ASAP7_75t_L g1444 ( .A1(n_1313), .A2(n_1403), .B1(n_1445), .B2(n_1446), .C1(n_1447), .C2(n_1449), .Y(n_1444) );
OAI211xp5_ASAP7_75t_L g1347 ( .A1(n_1314), .A2(n_1348), .B(n_1353), .C(n_1356), .Y(n_1347) );
INVx2_ASAP7_75t_L g1409 ( .A(n_1314), .Y(n_1409) );
O2A1O1Ixp33_ASAP7_75t_L g1430 ( .A1(n_1314), .A2(n_1371), .B(n_1397), .C(n_1431), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1314), .B(n_1473), .Y(n_1472) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1315), .B(n_1357), .Y(n_1356) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
OAI211xp5_ASAP7_75t_SL g1421 ( .A1(n_1317), .A2(n_1379), .B(n_1422), .C(n_1423), .Y(n_1421) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1318), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1319), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1319), .B(n_1376), .Y(n_1375) );
NAND2xp5_ASAP7_75t_SL g1417 ( .A(n_1319), .B(n_1327), .Y(n_1417) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1320), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1320), .B(n_1375), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1320), .B(n_1441), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1322), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1321), .B(n_1352), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1321), .B(n_1352), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1324), .Y(n_1449) );
O2A1O1Ixp33_ASAP7_75t_SL g1325 ( .A1(n_1326), .A2(n_1328), .B(n_1332), .C(n_1339), .Y(n_1325) );
INVx2_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
OAI21xp5_ASAP7_75t_SL g1432 ( .A1(n_1327), .A2(n_1433), .B(n_1434), .Y(n_1432) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NOR2xp33_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1330), .B(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
AOI21xp33_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1336), .B(n_1337), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g1423 ( .A1(n_1336), .A2(n_1359), .B1(n_1384), .B2(n_1424), .C(n_1426), .Y(n_1423) );
AOI21xp33_ASAP7_75t_L g1431 ( .A1(n_1336), .A2(n_1337), .B(n_1402), .Y(n_1431) );
OAI21xp5_ASAP7_75t_L g1367 ( .A1(n_1338), .A2(n_1368), .B(n_1371), .Y(n_1367) );
CKINVDCx6p67_ASAP7_75t_R g1386 ( .A(n_1338), .Y(n_1386) );
INVx3_ASAP7_75t_L g1361 ( .A(n_1339), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1339), .B(n_1407), .Y(n_1406) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1340), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_1340), .Y(n_1379) );
OAI22xp5_ASAP7_75t_SL g1341 ( .A1(n_1342), .A2(n_1343), .B1(n_1344), .B2(n_1345), .Y(n_1341) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1350), .B(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1350), .Y(n_1390) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
A2O1A1Ixp33_ASAP7_75t_L g1463 ( .A1(n_1354), .A2(n_1407), .B(n_1442), .C(n_1464), .Y(n_1463) );
AND2x2_ASAP7_75t_SL g1471 ( .A(n_1355), .B(n_1376), .Y(n_1471) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1356), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1360), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1359), .B(n_1366), .Y(n_1433) );
O2A1O1Ixp33_ASAP7_75t_L g1439 ( .A1(n_1361), .A2(n_1376), .B(n_1440), .C(n_1442), .Y(n_1439) );
NAND3xp33_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1367), .C(n_1374), .Y(n_1362) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
OAI211xp5_ASAP7_75t_L g1429 ( .A1(n_1369), .A2(n_1386), .B(n_1430), .C(n_1432), .Y(n_1429) );
AOI211xp5_ASAP7_75t_L g1393 ( .A1(n_1371), .A2(n_1394), .B(n_1395), .C(n_1401), .Y(n_1393) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1373), .Y(n_1469) );
OAI21xp5_ASAP7_75t_L g1387 ( .A1(n_1376), .A2(n_1388), .B(n_1392), .Y(n_1387) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
AOI22xp5_ASAP7_75t_L g1378 ( .A1(n_1379), .A2(n_1380), .B1(n_1405), .B2(n_1408), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1387), .C(n_1393), .Y(n_1380) );
INVxp67_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
NOR2xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1385), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
AOI211xp5_ASAP7_75t_L g1457 ( .A1(n_1388), .A2(n_1407), .B(n_1458), .C(n_1460), .Y(n_1457) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1391), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1391), .B(n_1424), .Y(n_1459) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1391), .Y(n_1468) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVxp33_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1410), .Y(n_1408) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_1409), .A2(n_1453), .B(n_1471), .Y(n_1470) );
AOI221xp5_ASAP7_75t_SL g1411 ( .A1(n_1412), .A2(n_1427), .B1(n_1428), .B2(n_1435), .C(n_1437), .Y(n_1411) );
O2A1O1Ixp33_ASAP7_75t_L g1412 ( .A1(n_1413), .A2(n_1415), .B(n_1416), .C(n_1421), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVxp67_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
AOI211xp5_ASAP7_75t_L g1437 ( .A1(n_1429), .A2(n_1438), .B(n_1439), .C(n_1444), .Y(n_1437) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1433), .Y(n_1445) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
A2O1A1Ixp33_ASAP7_75t_L g1450 ( .A1(n_1438), .A2(n_1451), .B(n_1457), .C(n_1463), .Y(n_1450) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
CKINVDCx14_ASAP7_75t_R g1447 ( .A(n_1448), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1448), .B(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVxp67_ASAP7_75t_SL g1460 ( .A(n_1461), .Y(n_1460) );
OAI211xp5_ASAP7_75t_SL g1464 ( .A1(n_1465), .A2(n_1466), .B(n_1470), .C(n_1472), .Y(n_1464) );
INVxp67_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_SL g1467 ( .A(n_1468), .B(n_1469), .Y(n_1467) );
CKINVDCx20_ASAP7_75t_R g1474 ( .A(n_1475), .Y(n_1474) );
CKINVDCx20_ASAP7_75t_R g1475 ( .A(n_1476), .Y(n_1475) );
INVx4_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
BUFx2_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
NAND3xp33_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1508), .C(n_1524), .Y(n_1481) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1499), .Y(n_1482) );
OAI22xp5_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1486), .B1(n_1487), .B2(n_1488), .Y(n_1484) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
OAI22xp5_ASAP7_75t_L g1504 ( .A1(n_1492), .A2(n_1498), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
OAI31xp33_ASAP7_75t_L g1508 ( .A1(n_1509), .A2(n_1512), .A3(n_1521), .B(n_1523), .Y(n_1508) );
INVx2_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
HB1xp67_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVxp67_ASAP7_75t_SL g1514 ( .A(n_1515), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_1518), .A2(n_1528), .B1(n_1530), .B2(n_1531), .Y(n_1527) );
OAI31xp33_ASAP7_75t_L g1524 ( .A1(n_1525), .A2(n_1532), .A3(n_1536), .B(n_1538), .Y(n_1524) );
BUFx3_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
HB1xp67_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx2_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
HB1xp67_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
BUFx3_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVxp33_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
HB1xp67_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1565), .Y(n_1551) );
NAND3xp33_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1571), .C(n_1575), .Y(n_1566) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
endmodule