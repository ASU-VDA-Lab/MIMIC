module real_aes_1965_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_783, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_783;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_156;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_0), .B(n_118), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_1), .A2(n_127), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_2), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_3), .B(n_118), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_4), .B(n_134), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_5), .B(n_134), .Y(n_478) );
INVx1_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_7), .B(n_134), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_8), .Y(n_454) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_9), .B(n_136), .Y(n_533) );
AND2x2_ASAP7_75t_L g154 ( .A(n_10), .B(n_143), .Y(n_154) );
AND2x2_ASAP7_75t_L g165 ( .A(n_11), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
AOI221x1_ASAP7_75t_L g482 ( .A1(n_13), .A2(n_24), .B1(n_118), .B2(n_127), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_14), .B(n_134), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_15), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_16), .B(n_118), .Y(n_529) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_17), .A2(n_143), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_18), .B(n_138), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_19), .B(n_134), .Y(n_522) );
AO21x1_ASAP7_75t_L g473 ( .A1(n_20), .A2(n_118), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_21), .B(n_118), .Y(n_222) );
INVx1_ASAP7_75t_L g444 ( .A(n_22), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_23), .A2(n_90), .B1(n_118), .B2(n_171), .Y(n_170) );
NAND2x1_ASAP7_75t_L g493 ( .A(n_25), .B(n_134), .Y(n_493) );
NAND2x1_ASAP7_75t_L g547 ( .A(n_26), .B(n_136), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_27), .Y(n_450) );
OR2x2_ASAP7_75t_L g141 ( .A(n_28), .B(n_87), .Y(n_141) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_28), .A2(n_87), .B(n_140), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_29), .B(n_136), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_30), .B(n_134), .Y(n_532) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_31), .A2(n_166), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_32), .B(n_136), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_33), .A2(n_127), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_34), .B(n_134), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_35), .A2(n_127), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g124 ( .A(n_36), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g128 ( .A(n_36), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g179 ( .A(n_36), .Y(n_179) );
OR2x6_ASAP7_75t_L g442 ( .A(n_37), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_38), .B(n_118), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_39), .B(n_118), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_40), .B(n_134), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_41), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_42), .B(n_136), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_43), .B(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_SL g461 ( .A1(n_44), .A2(n_66), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_44), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_45), .A2(n_85), .B1(n_429), .B2(n_430), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_45), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_46), .A2(n_127), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_47), .A2(n_127), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_48), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_49), .B(n_136), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_50), .B(n_118), .Y(n_214) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_51), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g121 ( .A(n_52), .Y(n_121) );
INVx1_ASAP7_75t_L g131 ( .A(n_52), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_53), .B(n_134), .Y(n_163) );
AND2x2_ASAP7_75t_L g203 ( .A(n_54), .B(n_138), .Y(n_203) );
XOR2xp5_ASAP7_75t_L g459 ( .A(n_55), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_56), .B(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_57), .B(n_134), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_58), .B(n_136), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_59), .A2(n_127), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_60), .B(n_118), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_61), .B(n_118), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_62), .A2(n_127), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g228 ( .A(n_63), .B(n_139), .Y(n_228) );
AO21x1_ASAP7_75t_L g475 ( .A1(n_64), .A2(n_127), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_65), .B(n_118), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_66), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_67), .B(n_136), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_68), .B(n_118), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_69), .B(n_136), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_70), .A2(n_94), .B1(n_127), .B2(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_71), .B(n_134), .Y(n_225) );
AND2x2_ASAP7_75t_L g506 ( .A(n_72), .B(n_139), .Y(n_506) );
INVx1_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
INVx1_ASAP7_75t_L g129 ( .A(n_73), .Y(n_129) );
AND2x2_ASAP7_75t_L g550 ( .A(n_74), .B(n_166), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_75), .B(n_136), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_76), .A2(n_127), .B(n_207), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_77), .A2(n_127), .B(n_132), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_78), .A2(n_127), .B(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g239 ( .A(n_79), .B(n_139), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_80), .B(n_138), .Y(n_168) );
INVx1_ASAP7_75t_L g445 ( .A(n_81), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_82), .B(n_118), .Y(n_524) );
AND2x2_ASAP7_75t_L g536 ( .A(n_83), .B(n_166), .Y(n_536) );
AND2x2_ASAP7_75t_L g142 ( .A(n_84), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_85), .Y(n_429) );
AND2x2_ASAP7_75t_L g474 ( .A(n_86), .B(n_210), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_88), .A2(n_104), .B1(n_451), .B2(n_456), .C1(n_769), .C2(n_775), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_88), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_88), .B(n_105), .C(n_435), .Y(n_447) );
AND2x2_ASAP7_75t_L g496 ( .A(n_88), .B(n_166), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_89), .B(n_136), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_91), .B(n_134), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_92), .B(n_136), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_93), .A2(n_127), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_95), .A2(n_127), .B(n_224), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g426 ( .A1(n_96), .A2(n_427), .B1(n_428), .B2(n_431), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_96), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_97), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_98), .B(n_134), .Y(n_541) );
BUFx2_ASAP7_75t_L g227 ( .A(n_99), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_100), .A2(n_442), .B1(n_458), .B2(n_765), .Y(n_457) );
BUFx2_ASAP7_75t_L g455 ( .A(n_101), .Y(n_455) );
BUFx2_ASAP7_75t_SL g779 ( .A(n_101), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_102), .A2(n_127), .B(n_531), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_434), .B(n_447), .C(n_448), .Y(n_104) );
AOI22x1_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_426), .B1(n_432), .B2(n_433), .Y(n_105) );
INVx3_ASAP7_75t_L g433 ( .A(n_106), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_106), .A2(n_465), .B1(n_763), .B2(n_764), .Y(n_464) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_339), .Y(n_106) );
NOR4xp75_ASAP7_75t_L g107 ( .A(n_108), .B(n_262), .C(n_287), .D(n_314), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_198), .B(n_240), .Y(n_108) );
NOR4xp25_ASAP7_75t_L g109 ( .A(n_110), .B(n_182), .C(n_189), .D(n_193), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_155), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_145), .Y(n_113) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_114), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_114), .B(n_186), .Y(n_333) );
AND2x2_ASAP7_75t_L g358 ( .A(n_114), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_114), .B(n_167), .Y(n_383) );
AND2x2_ASAP7_75t_L g424 ( .A(n_114), .B(n_191), .Y(n_424) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_SL g195 ( .A(n_115), .B(n_188), .Y(n_195) );
AND2x2_ASAP7_75t_L g197 ( .A(n_115), .B(n_157), .Y(n_197) );
NOR2x1_ASAP7_75t_L g248 ( .A(n_115), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g259 ( .A(n_115), .Y(n_259) );
AND2x2_ASAP7_75t_L g265 ( .A(n_115), .B(n_191), .Y(n_265) );
BUFx2_ASAP7_75t_L g278 ( .A(n_115), .Y(n_278) );
AND2x4_ASAP7_75t_L g309 ( .A(n_115), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g356 ( .A(n_115), .B(n_357), .Y(n_356) );
OR2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_142), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_126), .B(n_138), .Y(n_116) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_124), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
AND2x6_ASAP7_75t_L g136 ( .A(n_120), .B(n_129), .Y(n_136) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g134 ( .A(n_122), .B(n_131), .Y(n_134) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx5_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
AND2x2_ASAP7_75t_L g130 ( .A(n_125), .B(n_131), .Y(n_130) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
AND2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
BUFx3_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
INVx2_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
AND2x4_ASAP7_75t_L g177 ( .A(n_130), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g173 ( .A(n_131), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .B(n_137), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_136), .B(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_137), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_137), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_137), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_137), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_137), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_137), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_137), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_137), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_137), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_137), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_137), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_137), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_137), .A2(n_547), .B(n_548), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_138), .Y(n_147) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_138), .A2(n_170), .B(n_176), .Y(n_169) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_138), .A2(n_482), .B(n_486), .Y(n_481) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_138), .A2(n_482), .B(n_486), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_138), .A2(n_538), .B(n_539), .Y(n_537) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g210 ( .A(n_140), .B(n_141), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_143), .A2(n_222), .B(n_223), .Y(n_221) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx1_ASAP7_75t_L g350 ( .A(n_145), .Y(n_350) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
AND2x2_ASAP7_75t_L g191 ( .A(n_146), .B(n_157), .Y(n_191) );
AOI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_154), .Y(n_146) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_147), .A2(n_544), .B(n_550), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_155), .B(n_368), .Y(n_421) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
OR2x2_ASAP7_75t_L g258 ( .A(n_156), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_167), .Y(n_156) );
INVx2_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
INVx2_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
AND2x2_ASAP7_75t_L g359 ( .A(n_157), .B(n_188), .Y(n_359) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_165), .Y(n_157) );
INVx4_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
INVx3_ASAP7_75t_L g232 ( .A(n_166), .Y(n_232) );
INVx2_ASAP7_75t_L g247 ( .A(n_167), .Y(n_247) );
BUFx3_ASAP7_75t_L g264 ( .A(n_167), .Y(n_264) );
AND2x2_ASAP7_75t_L g291 ( .A(n_167), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x4_ASAP7_75t_L g184 ( .A(n_168), .B(n_169), .Y(n_184) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_175), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2x1p5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2x1_ASAP7_75t_L g182 ( .A(n_183), .B(n_185), .Y(n_182) );
INVx2_ASAP7_75t_L g192 ( .A(n_183), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_183), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g362 ( .A(n_183), .B(n_302), .Y(n_362) );
AND2x2_ASAP7_75t_L g386 ( .A(n_183), .B(n_195), .Y(n_386) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g282 ( .A(n_184), .B(n_187), .Y(n_282) );
AND2x2_ASAP7_75t_L g364 ( .A(n_184), .B(n_357), .Y(n_364) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_SL g407 ( .A(n_186), .Y(n_407) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g292 ( .A(n_187), .Y(n_292) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
INVx2_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
INVx1_ASAP7_75t_L g310 ( .A(n_188), .Y(n_310) );
AOI222xp33_ASAP7_75t_SL g240 ( .A1(n_189), .A2(n_241), .B1(n_245), .B2(n_250), .C1(n_257), .C2(n_260), .Y(n_240) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g317 ( .A(n_191), .Y(n_317) );
BUFx2_ASAP7_75t_L g346 ( .A(n_191), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g340 ( .A1(n_192), .A2(n_341), .B(n_345), .C(n_353), .Y(n_340) );
OR2x2_ASAP7_75t_L g411 ( .A(n_192), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g419 ( .A(n_192), .B(n_324), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_195), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g394 ( .A(n_195), .B(n_282), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_195), .B(n_374), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_196), .B(n_264), .Y(n_402) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g324 ( .A(n_197), .B(n_296), .Y(n_324) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_219), .Y(n_199) );
INVx1_ASAP7_75t_L g418 ( .A(n_200), .Y(n_418) );
NOR2xp67_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g261 ( .A(n_201), .B(n_220), .Y(n_261) );
INVx1_ASAP7_75t_L g338 ( .A(n_201), .Y(n_338) );
OR2x2_ASAP7_75t_L g397 ( .A(n_201), .B(n_220), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_201), .B(n_269), .Y(n_403) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
OR2x2_ASAP7_75t_L g276 ( .A(n_202), .B(n_230), .Y(n_276) );
AND2x2_ASAP7_75t_L g285 ( .A(n_202), .B(n_212), .Y(n_285) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_202), .B(n_220), .Y(n_313) );
AND2x2_ASAP7_75t_L g360 ( .A(n_202), .B(n_255), .Y(n_360) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_210), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_210), .A2(n_214), .B(n_215), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_210), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g518 ( .A(n_210), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_210), .A2(n_529), .B(n_530), .Y(n_528) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
INVx1_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
AND2x2_ASAP7_75t_L g269 ( .A(n_212), .B(n_256), .Y(n_269) );
INVx2_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
OR2x2_ASAP7_75t_L g370 ( .A(n_212), .B(n_220), .Y(n_370) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
NOR2x1_ASAP7_75t_SL g255 ( .A(n_220), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g273 ( .A(n_220), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g286 ( .A(n_220), .B(n_230), .Y(n_286) );
BUFx2_ASAP7_75t_L g305 ( .A(n_220), .Y(n_305) );
INVx2_ASAP7_75t_SL g332 ( .A(n_220), .Y(n_332) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_228), .Y(n_220) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g242 ( .A(n_230), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g388 ( .A(n_230), .B(n_330), .Y(n_388) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_231) );
AO21x1_ASAP7_75t_SL g256 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_256) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_232), .A2(n_490), .B(n_496), .Y(n_489) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_232), .A2(n_500), .B(n_506), .Y(n_499) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_232), .A2(n_490), .B(n_496), .Y(n_511) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_232), .A2(n_500), .B(n_506), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_238), .Y(n_233) );
AOI211xp5_ASAP7_75t_L g404 ( .A1(n_241), .A2(n_265), .B(n_405), .C(n_409), .Y(n_404) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_242), .B(n_320), .Y(n_355) );
BUFx2_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
OR2x2_ASAP7_75t_L g267 ( .A(n_244), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g352 ( .A(n_244), .B(n_286), .Y(n_352) );
AND2x2_ASAP7_75t_L g373 ( .A(n_244), .B(n_329), .Y(n_373) );
INVx2_ASAP7_75t_L g380 ( .A(n_244), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_245), .A2(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g327 ( .A(n_246), .B(n_309), .Y(n_327) );
OR2x2_ASAP7_75t_L g406 ( .A(n_246), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_247), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_249), .Y(n_280) );
AND2x2_ASAP7_75t_L g357 ( .A(n_249), .B(n_304), .Y(n_357) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_SL g351 ( .A(n_252), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_252), .B(n_261), .Y(n_384) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g260 ( .A(n_253), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g379 ( .A(n_254), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g329 ( .A(n_255), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g299 ( .A(n_256), .B(n_274), .Y(n_299) );
OAI31xp33_ASAP7_75t_L g306 ( .A1(n_257), .A2(n_307), .A3(n_309), .B(n_311), .Y(n_306) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_259), .B(n_282), .Y(n_308) );
AO21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_270), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g318 ( .A(n_264), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g423 ( .A(n_264), .Y(n_423) );
INVx2_ASAP7_75t_SL g408 ( .A(n_265), .Y(n_408) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g396 ( .A(n_268), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_269), .B(n_332), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_277), .B1(n_281), .B2(n_283), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_271), .A2(n_390), .B(n_391), .Y(n_389) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g330 ( .A(n_274), .Y(n_330) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g344 ( .A(n_276), .B(n_305), .Y(n_344) );
OR2x2_ASAP7_75t_L g369 ( .A(n_276), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_278), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_278), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g368 ( .A(n_278), .Y(n_368) );
INVx2_ASAP7_75t_L g297 ( .A(n_279), .Y(n_297) );
INVx1_ASAP7_75t_L g377 ( .A(n_280), .Y(n_377) );
AND2x2_ASAP7_75t_L g300 ( .A(n_282), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g374 ( .A(n_282), .Y(n_374) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_306), .Y(n_287) );
OAI321xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_293), .A3(n_298), .B1(n_299), .B2(n_300), .C(n_305), .Y(n_288) );
AOI322xp5_ASAP7_75t_L g414 ( .A1(n_289), .A2(n_320), .A3(n_415), .B1(n_417), .B2(n_419), .C1(n_420), .C2(n_425), .Y(n_414) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g367 ( .A(n_292), .Y(n_367) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_294), .B(n_374), .Y(n_391) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g399 ( .A(n_297), .Y(n_399) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp33_ASAP7_75t_SL g331 ( .A(n_299), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_SL g398 ( .A1(n_302), .A2(n_308), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g320 ( .A(n_313), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_334), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B1(n_321), .B2(n_322), .C(n_325), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
AND2x2_ASAP7_75t_L g321 ( .A(n_319), .B(n_320), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_328), .B1(n_331), .B2(n_333), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g337 ( .A(n_329), .B(n_338), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_332), .A2(n_421), .B(n_422), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR3xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_371), .C(n_392), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_379), .B1(n_406), .B2(n_408), .Y(n_405) );
OAI21xp33_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B(n_351), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_346), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_352), .A2(n_394), .B1(n_395), .B2(n_398), .C(n_400), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B1(n_358), .B2(n_360), .C(n_361), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
INVx1_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
INVx1_ASAP7_75t_SL g410 ( .A(n_358), .Y(n_410) );
AOI31xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .A3(n_365), .B(n_369), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_362), .A2(n_372), .B1(n_374), .B2(n_375), .C(n_783), .Y(n_371) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_381), .C(n_389), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g387 ( .A(n_380), .B(n_388), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
BUFx2_ASAP7_75t_SL g425 ( .A(n_388), .Y(n_425) );
NAND3xp33_ASAP7_75t_SL g392 ( .A(n_393), .B(n_404), .C(n_414), .Y(n_392) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_403), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_413), .Y(n_409) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g432 ( .A(n_426), .Y(n_432) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_435), .B(n_446), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_437), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g774 ( .A(n_439), .Y(n_774) );
BUFx2_ASAP7_75t_L g781 ( .A(n_439), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_440), .Y(n_764) );
OR2x2_ASAP7_75t_L g768 ( .A(n_440), .B(n_442), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_SL g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx2_ASAP7_75t_L g773 ( .A(n_453), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_453), .A2(n_777), .B(n_780), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_455), .B(n_773), .Y(n_772) );
INVxp33_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_464), .Y(n_458) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_662), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_599), .C(n_622), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_551), .C(n_568), .Y(n_467) );
OAI31xp33_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_487), .A3(n_507), .B(n_514), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_469), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .Y(n_470) );
AND2x4_ASAP7_75t_L g554 ( .A(n_471), .B(n_481), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_471), .B(n_498), .Y(n_583) );
AND2x4_ASAP7_75t_L g585 ( .A(n_471), .B(n_579), .Y(n_585) );
AND2x2_ASAP7_75t_L g716 ( .A(n_471), .B(n_511), .Y(n_716) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g561 ( .A(n_472), .Y(n_561) );
OAI21x1_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_475), .B(n_479), .Y(n_472) );
INVx1_ASAP7_75t_L g480 ( .A(n_474), .Y(n_480) );
AND2x2_ASAP7_75t_L g497 ( .A(n_481), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_481), .B(n_560), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_481), .B(n_499), .Y(n_658) );
AND2x2_ASAP7_75t_L g747 ( .A(n_481), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g729 ( .A(n_487), .Y(n_729) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
BUFx2_ASAP7_75t_L g558 ( .A(n_488), .Y(n_558) );
AND2x2_ASAP7_75t_L g592 ( .A(n_488), .B(n_498), .Y(n_592) );
AND2x2_ASAP7_75t_L g641 ( .A(n_488), .B(n_499), .Y(n_641) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g598 ( .A(n_489), .B(n_499), .Y(n_598) );
INVxp67_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
BUFx3_ASAP7_75t_L g655 ( .A(n_489), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g551 ( .A1(n_497), .A2(n_552), .A3(n_557), .B(n_562), .Y(n_551) );
AND2x2_ASAP7_75t_L g559 ( .A(n_498), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g578 ( .A(n_499), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_501), .B(n_505), .Y(n_500) );
AOI322xp5_ASAP7_75t_L g752 ( .A1(n_507), .A2(n_627), .A3(n_656), .B1(n_661), .B2(n_753), .C1(n_756), .C2(n_757), .Y(n_752) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_508), .B(n_598), .Y(n_603) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_508), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g684 ( .A(n_508), .B(n_588), .Y(n_684) );
INVx1_ASAP7_75t_SL g698 ( .A(n_508), .Y(n_698) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g579 ( .A(n_509), .Y(n_579) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_509), .Y(n_722) );
AND2x2_ASAP7_75t_L g651 ( .A(n_510), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_510), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_SL g510 ( .A(n_511), .B(n_512), .Y(n_510) );
BUFx2_ASAP7_75t_L g556 ( .A(n_511), .Y(n_556) );
INVx1_ASAP7_75t_L g748 ( .A(n_511), .Y(n_748) );
OR2x2_ASAP7_75t_L g615 ( .A(n_512), .B(n_560), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_512), .B(n_585), .Y(n_649) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g588 ( .A(n_513), .B(n_560), .Y(n_588) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_534), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g644 ( .A(n_516), .Y(n_644) );
OR2x2_ASAP7_75t_L g671 ( .A(n_516), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
NOR2x1_ASAP7_75t_SL g565 ( .A(n_517), .B(n_535), .Y(n_565) );
AND2x2_ASAP7_75t_L g572 ( .A(n_517), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g744 ( .A(n_517), .B(n_606), .Y(n_744) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_518), .B(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g621 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
OR2x2_ASAP7_75t_L g566 ( .A(n_527), .B(n_567), .Y(n_566) );
BUFx3_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
INVx2_ASAP7_75t_L g606 ( .A(n_527), .Y(n_606) );
INVx1_ASAP7_75t_L g647 ( .A(n_527), .Y(n_647) );
AND2x2_ASAP7_75t_L g678 ( .A(n_527), .B(n_535), .Y(n_678) );
AND2x2_ASAP7_75t_L g709 ( .A(n_527), .B(n_636), .Y(n_709) );
AND2x2_ASAP7_75t_L g605 ( .A(n_534), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_534), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_534), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g713 ( .A(n_534), .B(n_575), .Y(n_713) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_543), .Y(n_534) );
INVx5_ASAP7_75t_L g573 ( .A(n_535), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_535), .B(n_567), .Y(n_645) );
BUFx2_ASAP7_75t_L g705 ( .A(n_535), .Y(n_705) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx4_ASAP7_75t_L g567 ( .A(n_543), .Y(n_567) );
AND2x2_ASAP7_75t_L g690 ( .A(n_543), .B(n_573), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_553), .A2(n_680), .B1(n_683), .B2(n_685), .C(n_686), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g701 ( .A(n_554), .B(n_592), .Y(n_701) );
INVx1_ASAP7_75t_SL g727 ( .A(n_554), .Y(n_727) );
AND2x2_ASAP7_75t_L g712 ( .A(n_555), .B(n_684), .Y(n_712) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_556), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g581 ( .A(n_558), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g587 ( .A(n_558), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g611 ( .A(n_559), .Y(n_611) );
AND2x2_ASAP7_75t_L g669 ( .A(n_559), .B(n_597), .Y(n_669) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g594 ( .A(n_561), .Y(n_594) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g590 ( .A(n_566), .Y(n_590) );
OR2x2_ASAP7_75t_L g758 ( .A(n_566), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g574 ( .A(n_567), .Y(n_574) );
AND2x4_ASAP7_75t_L g630 ( .A(n_567), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_567), .B(n_635), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_567), .B(n_573), .Y(n_672) );
AND2x2_ASAP7_75t_L g732 ( .A(n_567), .B(n_635), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_576), .B1(n_589), .B2(n_591), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_569), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND3x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .C(n_575), .Y(n_571) );
AND2x4_ASAP7_75t_L g589 ( .A(n_572), .B(n_590), .Y(n_589) );
INVx4_ASAP7_75t_L g629 ( .A(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_SL g762 ( .A(n_573), .B(n_630), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_574), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g674 ( .A(n_575), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g739 ( .A1(n_575), .A2(n_704), .A3(n_740), .B1(n_742), .B2(n_745), .C1(n_749), .C2(n_750), .Y(n_739) );
NAND4xp25_ASAP7_75t_SL g576 ( .A(n_577), .B(n_580), .C(n_584), .D(n_586), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_SL g706 ( .A(n_578), .B(n_594), .Y(n_706) );
BUFx2_ASAP7_75t_L g597 ( .A(n_579), .Y(n_597) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g721 ( .A(n_582), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g735 ( .A(n_583), .B(n_610), .Y(n_735) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g601 ( .A(n_585), .B(n_602), .Y(n_601) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_585), .A2(n_654), .B(n_656), .C(n_659), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_585), .B(n_592), .Y(n_711) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_587), .A2(n_669), .B1(n_670), .B2(n_673), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_588), .A2(n_624), .B1(n_628), .B2(n_632), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_588), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_588), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_588), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g755 ( .A(n_588), .Y(n_755) );
INVx1_ASAP7_75t_L g694 ( .A(n_589), .Y(n_694) );
OAI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g602 ( .A(n_592), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_592), .B(n_597), .Y(n_751) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g687 ( .A(n_594), .B(n_598), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_596), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g754 ( .A(n_597), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g728 ( .A(n_598), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B(n_604), .C(n_607), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_SL g714 ( .A1(n_602), .A2(n_633), .B1(n_680), .B2(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_606), .B(n_629), .Y(n_637) );
OR2x2_ASAP7_75t_L g666 ( .A(n_606), .B(n_667), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_612), .B(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_613), .A2(n_666), .B(n_668), .C(n_676), .Y(n_665) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp67_ASAP7_75t_SL g699 ( .A(n_618), .B(n_645), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_618), .Y(n_702) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_620), .B(n_629), .Y(n_759) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g631 ( .A(n_621), .Y(n_631) );
INVx2_ASAP7_75t_L g636 ( .A(n_621), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_638), .C(n_650), .D(n_653), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_626), .A2(n_758), .B1(n_760), .B2(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x4_ASAP7_75t_L g725 ( .A(n_629), .B(n_655), .Y(n_725) );
AND2x2_ASAP7_75t_L g646 ( .A(n_630), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g667 ( .A(n_630), .Y(n_667) );
AND2x2_ASAP7_75t_L g677 ( .A(n_630), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_636), .Y(n_691) );
INVx1_ASAP7_75t_L g681 ( .A(n_637), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .A3(n_645), .B1(n_646), .B2(n_648), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_639), .A2(n_687), .B(n_688), .Y(n_686) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_642), .A2(n_719), .B1(n_721), .B2(n_723), .C(n_726), .Y(n_718) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g703 ( .A(n_644), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g661 ( .A(n_645), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_646), .A2(n_684), .B1(n_734), .B2(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g660 ( .A(n_647), .Y(n_660) );
AND2x2_ASAP7_75t_L g738 ( .A(n_647), .B(n_691), .Y(n_738) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_654), .B(n_706), .Y(n_741) );
INVx1_ASAP7_75t_L g760 ( .A(n_654), .Y(n_760) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_663), .B(n_717), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_707), .Y(n_663) );
NOR3xp33_ASAP7_75t_SL g664 ( .A(n_665), .B(n_679), .C(n_692), .Y(n_664) );
INVx1_ASAP7_75t_L g682 ( .A(n_667), .Y(n_682) );
INVx1_ASAP7_75t_SL g693 ( .A(n_669), .Y(n_693) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g675 ( .A(n_672), .Y(n_675) );
INVx2_ASAP7_75t_L g685 ( .A(n_673), .Y(n_685) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x4_ASAP7_75t_L g731 ( .A(n_674), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g749 ( .A(n_678), .B(n_732), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g700 ( .A1(n_689), .A2(n_701), .A3(n_702), .B1(n_703), .B2(n_706), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_689), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g720 ( .A(n_691), .Y(n_720) );
OAI211xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_694), .B(n_695), .C(n_700), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g756 ( .A(n_704), .B(n_744), .Y(n_756) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_705), .B(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_707) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_718), .B(n_733), .C(n_739), .D(n_752), .Y(n_717) );
INVxp33_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_729), .C(n_730), .Y(n_726) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx3_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .Y(n_770) );
INVxp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx8_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
endmodule