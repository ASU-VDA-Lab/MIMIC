module fake_aes_687_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_7;
INVx1_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_2), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx5_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_8), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_14) );
NOR3xp33_ASAP7_75t_SL g15 ( .A(n_7), .B(n_9), .C(n_12), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_10), .B(n_3), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_11), .B(n_4), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
NAND2x1_ASAP7_75t_L g19 ( .A(n_15), .B(n_14), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
OAI211xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_16), .B(n_17), .C(n_13), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_6), .Y(n_27) );
endmodule