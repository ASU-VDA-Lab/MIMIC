module real_jpeg_13709_n_17 (n_5, n_4, n_8, n_0, n_12, n_310, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_310;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx2_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_3),
.B(n_176),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_29),
.B(n_30),
.C(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_44),
.C(n_47),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_3),
.B(n_31),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_3),
.A2(n_124),
.B(n_247),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_147),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_153),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_5),
.A2(n_44),
.B1(n_48),
.B2(n_153),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_94),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_6),
.A2(n_44),
.B1(n_48),
.B2(n_94),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_36),
.B1(n_44),
.B2(n_48),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_66),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_9),
.A2(n_44),
.B1(n_48),
.B2(n_66),
.Y(n_167)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_11),
.B(n_27),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_12),
.A2(n_44),
.B1(n_48),
.B2(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_13),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_133),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_13),
.A2(n_44),
.B1(n_48),
.B2(n_133),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_44),
.B1(n_48),
.B2(n_60),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_15),
.A2(n_39),
.B1(n_44),
.B2(n_48),
.Y(n_123)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_20),
.B(n_95),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_68),
.C(n_76),
.Y(n_20)
);

FAx1_ASAP7_75t_L g110 ( 
.A(n_21),
.B(n_68),
.CI(n_76),
.CON(n_110),
.SN(n_110)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_21)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_41),
.C(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_26),
.A2(n_32),
.B(n_147),
.Y(n_222)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_30),
.A2(n_59),
.A3(n_63),
.B1(n_149),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_31),
.B(n_173),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_33),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_38),
.A2(n_70),
.B1(n_72),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_40),
.A2(n_41),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_51),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_49),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_42),
.A2(n_49),
.B1(n_87),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_42),
.A2(n_49),
.B1(n_128),
.B2(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_42),
.B(n_159),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_42),
.A2(n_49),
.B1(n_217),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_52),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_43),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_43),
.A2(n_158),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_43),
.B(n_147),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_48),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_49),
.B(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_56),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_62),
.B(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_61),
.B(n_147),
.C(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_61),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_61),
.A2(n_62),
.B1(n_132),
.B2(n_193),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_62),
.A2(n_90),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_69),
.B(n_73),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_70),
.A2(n_72),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_70),
.A2(n_154),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_70),
.A2(n_191),
.B(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_72),
.A2(n_152),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_72),
.A2(n_130),
.B(n_172),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_74),
.A2(n_216),
.B(n_218),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_74),
.A2(n_218),
.B(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B(n_89),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_78),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_81),
.A2(n_82),
.B1(n_123),
.B2(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_81),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_81),
.A2(n_82),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_82),
.B(n_225),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_136),
.B(n_307),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_110),
.B(n_111),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_110),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_118),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_117),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_118),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_131),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_119),
.A2(n_120),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_125),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_124),
.A2(n_125),
.B1(n_167),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_124),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_125),
.A2(n_178),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_125),
.A2(n_224),
.B(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_125),
.B(n_147),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_129),
.B(n_131),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_301),
.B(n_306),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_289),
.B(n_300),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_196),
.A3(n_208),
.B1(n_287),
.B2(n_288),
.C(n_310),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_179),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_142),
.B(n_179),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_161),
.C(n_170),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_143),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_160),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_151),
.C(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_170),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_194),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_194),
.C(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_198),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_200),
.B(n_202),
.C(n_207),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_228),
.B(n_286),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_226),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_210),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_219),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_211),
.A2(n_212),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_215),
.A2(n_219),
.B1(n_220),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_221),
.B(n_223),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_279),
.B(n_285),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_267),
.B(n_278),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_248),
.B(n_266),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_265),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_254),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_260),
.B(n_264),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_269),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_274),
.C(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_299),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.C(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);


endmodule