module fake_netlist_1_6959_n_24 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_2), .B(n_10), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
AOI22xp33_ASAP7_75t_L g16 ( .A1(n_7), .A2(n_9), .B1(n_0), .B2(n_5), .Y(n_16) );
BUFx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
BUFx10_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OAI22xp5_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_16), .B1(n_13), .B2(n_15), .Y(n_21) );
OAI21xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_14), .B(n_11), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_14), .B1(n_12), .B2(n_1), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_4), .B(n_18), .Y(n_24) );
endmodule