module fake_jpeg_10873_n_382 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_55),
.B(n_88),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_60),
.A2(n_83),
.B1(n_51),
.B2(n_33),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_73),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_32),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_72),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_9),
.C(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_95),
.Y(n_107)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_26),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_23),
.B(n_3),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_32),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_104),
.Y(n_150)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_5),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_101),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_39),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_38),
.B1(n_18),
.B2(n_31),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_108),
.A2(n_125),
.B1(n_145),
.B2(n_158),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_111),
.B(n_119),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_21),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_43),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_142),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_38),
.B1(n_52),
.B2(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_21),
.B1(n_47),
.B2(n_44),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_137),
.B1(n_56),
.B2(n_67),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_68),
.B(n_51),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_33),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_75),
.A2(n_48),
.B1(n_47),
.B2(n_31),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_19),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_45),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_161),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_93),
.A2(n_48),
.B1(n_44),
.B2(n_25),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_90),
.A2(n_25),
.B1(n_28),
.B2(n_45),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_159),
.B1(n_141),
.B2(n_153),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_66),
.B(n_28),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_165),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_60),
.B1(n_105),
.B2(n_96),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_170),
.B1(n_189),
.B2(n_212),
.Y(n_240)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_62),
.B1(n_71),
.B2(n_77),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_206),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_197),
.B1(n_194),
.B2(n_184),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_129),
.A2(n_34),
.B(n_46),
.C(n_58),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_184),
.A2(n_194),
.B(n_196),
.C(n_190),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_65),
.C(n_46),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_102),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_186),
.B(n_200),
.Y(n_226)
);

FAx1_ASAP7_75t_L g187 ( 
.A(n_107),
.B(n_4),
.CI(n_5),
.CON(n_187),
.SN(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_187),
.A2(n_196),
.B(n_190),
.C(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_108),
.A2(n_5),
.B1(n_158),
.B2(n_145),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_106),
.B(n_5),
.CI(n_133),
.CON(n_192),
.SN(n_192)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_192),
.B(n_181),
.CI(n_193),
.CON(n_253),
.SN(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_147),
.B(n_125),
.C(n_151),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_134),
.B1(n_147),
.B2(n_141),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_201),
.Y(n_235)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_146),
.A2(n_140),
.B1(n_126),
.B2(n_128),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_205),
.B1(n_215),
.B2(n_172),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_120),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_117),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_123),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_152),
.C(n_126),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_140),
.A2(n_144),
.B1(n_156),
.B2(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_131),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_113),
.B(n_156),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_215),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_224),
.B1(n_234),
.B2(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_166),
.B1(n_168),
.B2(n_187),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_173),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_244),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_233),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_253),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_175),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_187),
.A2(n_189),
.B1(n_173),
.B2(n_203),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_195),
.B1(n_254),
.B2(n_250),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_SL g282 ( 
.A1(n_241),
.A2(n_249),
.B(n_256),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_212),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_169),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_167),
.Y(n_250)
);

A2O1A1O1Ixp25_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_192),
.B(n_182),
.C(n_210),
.D(n_213),
.Y(n_265)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_280),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_198),
.B1(n_204),
.B2(n_180),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_264),
.B1(n_268),
.B2(n_286),
.Y(n_288)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_180),
.B1(n_171),
.B2(n_178),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_282),
.B(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_269),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_177),
.B1(n_195),
.B2(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_270),
.B(n_273),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_278),
.B1(n_284),
.B2(n_285),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_244),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_225),
.B(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_220),
.B(n_238),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_253),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_233),
.C(n_242),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_235),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_242),
.B(n_219),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_241),
.B(n_252),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_219),
.B(n_240),
.Y(n_285)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_236),
.B1(n_252),
.B2(n_232),
.C(n_222),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_219),
.A2(n_241),
.B1(n_227),
.B2(n_230),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_295),
.B(n_262),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_296),
.B1(n_302),
.B2(n_269),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_241),
.B1(n_227),
.B2(n_237),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_258),
.A2(n_241),
.B1(n_227),
.B2(n_237),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_286),
.B1(n_259),
.B2(n_264),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_277),
.B(n_251),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_300),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_248),
.B1(n_222),
.B2(n_239),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_278),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_270),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_308),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_325),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_260),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_312),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_272),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_313),
.A2(n_293),
.B(n_290),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_317),
.B1(n_296),
.B2(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_275),
.B1(n_257),
.B2(n_261),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_318),
.B(n_323),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_267),
.C(n_291),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_268),
.B1(n_267),
.B2(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_289),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_327),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_263),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_324),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_335),
.C(n_336),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_SL g336 ( 
.A(n_316),
.B(n_289),
.C(n_291),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_303),
.B1(n_305),
.B2(n_301),
.Y(n_338)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_307),
.B(n_309),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_313),
.B(n_329),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_324),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_310),
.B1(n_314),
.B2(n_326),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_343),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_311),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_353),
.C(n_341),
.Y(n_361)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_334),
.A2(n_320),
.A3(n_326),
.B1(n_288),
.B2(n_312),
.C1(n_322),
.C2(n_316),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_345),
.B(n_346),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_327),
.Y(n_346)
);

AOI321xp33_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_324),
.A3(n_292),
.B1(n_301),
.B2(n_306),
.C(n_309),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_348),
.B(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_352),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_333),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_347),
.A2(n_351),
.B1(n_334),
.B2(n_350),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_347),
.A2(n_340),
.B1(n_339),
.B2(n_332),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_288),
.B1(n_337),
.B2(n_292),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_359),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_360),
.C(n_355),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_353),
.B(n_349),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_363),
.A2(n_366),
.B(n_348),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_344),
.C(n_331),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_367),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_357),
.B(n_359),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_365),
.B(n_266),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_354),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_372),
.B(n_373),
.C(n_368),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_358),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_287),
.C(n_281),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_SL g377 ( 
.A(n_375),
.B(n_273),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_377),
.A2(n_376),
.B(n_276),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_380),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_236),
.C(n_217),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_274),
.Y(n_382)
);


endmodule