module fake_netlist_6_2021_n_2567 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2567);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2567;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1674;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_1700;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_1815;
wire n_659;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_586;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2468;
wire n_1624;
wire n_1124;
wire n_515;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_2178;
wire n_701;
wire n_950;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_595;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_2012;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_2134;
wire n_1176;
wire n_1004;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1774;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_1475;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_527;
wire n_474;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_600;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1286;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_2181;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1397;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_1472;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_737;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1941;
wire n_1375;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_706;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1746;
wire n_1002;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_508;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1785;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1114;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1464;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_2221;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_424),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_121),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_143),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_265),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_130),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_390),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_44),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_406),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_232),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_362),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_129),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_300),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_174),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_153),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_341),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_20),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_230),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_26),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_197),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_86),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_353),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_64),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_45),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_388),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_40),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_24),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_104),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_229),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_10),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_299),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_77),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_21),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_169),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_2),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_273),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_69),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_83),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_190),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_413),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_340),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_357),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_36),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_393),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_63),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_4),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_21),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_187),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_284),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_360),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_185),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_95),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_133),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_73),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_332),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_81),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_224),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_117),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_366),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_261),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_49),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_249),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_120),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_75),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_79),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_68),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_405),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_416),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

BUFx5_ASAP7_75t_L g505 ( 
.A(n_233),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_130),
.Y(n_506)
);

INVx4_ASAP7_75t_R g507 ( 
.A(n_109),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_80),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_351),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_70),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_53),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_113),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_373),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_251),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_355),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_375),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_238),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_177),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_193),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_371),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_88),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_2),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_228),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_330),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_377),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_421),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_409),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_374),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_52),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_379),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_103),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_15),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_221),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_280),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_317),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_352),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_429),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_223),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_276),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_415),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_180),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_156),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_129),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_175),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_404),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_250),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_19),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_195),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_428),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_312),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_203),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_105),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_329),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_83),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_167),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_47),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_165),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_13),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_410),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_82),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_148),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_314),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_57),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_69),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_206),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_431),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_391),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_369),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_281),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_407),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_242),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_188),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_219),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_370),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_411),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_131),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_389),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_298),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_65),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_99),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_90),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_121),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_100),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_408),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_132),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_0),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_378),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_65),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_46),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_297),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_176),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_109),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_303),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_259),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_348),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_8),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_384),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_84),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_28),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_43),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_263),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_279),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_252),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_381),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_248),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_367),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_200),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_84),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_395),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_63),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_418),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_19),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_403),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_349),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_25),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_64),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_288),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_302),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_363),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_42),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_101),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_36),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_414),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_383),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_86),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_310),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_160),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_40),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_328),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_235),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_231),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_96),
.Y(n_633)
);

BUFx8_ASAP7_75t_SL g634 ( 
.A(n_42),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_22),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_247),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_114),
.Y(n_637)
);

CKINVDCx14_ASAP7_75t_R g638 ( 
.A(n_260),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_209),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_35),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_118),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_164),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_226),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_225),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_170),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_368),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_87),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_108),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_427),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_155),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_255),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_199),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_70),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_287),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_39),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_365),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_337),
.Y(n_657)
);

BUFx5_ASAP7_75t_L g658 ( 
.A(n_41),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_319),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_275),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_272),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_301),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_113),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_33),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_346),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_150),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_49),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_387),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_186),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_376),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_194),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_76),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_285),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_168),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_191),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_213),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_201),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_149),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_136),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_31),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_217),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_196),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_120),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_61),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_322),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_339),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_81),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_256),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_111),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_399),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_311),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_55),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_264),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_43),
.Y(n_694)
);

CKINVDCx16_ASAP7_75t_R g695 ( 
.A(n_34),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_202),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_16),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_343),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_396),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_326),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_211),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_152),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_372),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_98),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_4),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_394),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_158),
.Y(n_707)
);

BUFx2_ASAP7_75t_R g708 ( 
.A(n_432),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_106),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_382),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_335),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_134),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_204),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_91),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_422),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_107),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_364),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_124),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_82),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_24),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_132),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_392),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_400),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_106),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_30),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_98),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_100),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_320),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_430),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_11),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_61),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_91),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_262),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_53),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_291),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_307),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_77),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_111),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_417),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_59),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_283),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_12),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_44),
.Y(n_743)
);

CKINVDCx14_ASAP7_75t_R g744 ( 
.A(n_425),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_125),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_20),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_412),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_345),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_127),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_97),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_13),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_25),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_34),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_105),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_386),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_116),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_136),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_237),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_135),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_420),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_402),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_162),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_398),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_354),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_47),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_54),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_401),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_38),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_32),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_10),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_75),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_359),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_0),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_66),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_207),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_246),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_309),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_31),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_88),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_66),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_385),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_17),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_124),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_658),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_634),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_658),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_695),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_658),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_560),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_658),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_634),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_658),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_658),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_559),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_679),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_679),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_679),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_639),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_460),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_434),
.B(n_1),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_460),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_485),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_485),
.Y(n_804)
);

CKINVDCx14_ASAP7_75t_R g805 ( 
.A(n_638),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_547),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_547),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_656),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_639),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_433),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_714),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_439),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_672),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_693),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_714),
.Y(n_817)
);

CKINVDCx14_ASAP7_75t_R g818 ( 
.A(n_744),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_749),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_435),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_449),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_458),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_689),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_457),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_476),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_467),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_479),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_487),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_456),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_489),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_466),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_498),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_467),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_499),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_500),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_506),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_442),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_537),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_443),
.Y(n_840)
);

CKINVDCx16_ASAP7_75t_R g841 ( 
.A(n_612),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_510),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_767),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_484),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_511),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_554),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_505),
.Y(n_847)
);

INVxp33_ASAP7_75t_SL g848 ( 
.A(n_464),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_556),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_580),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_493),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_581),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_587),
.Y(n_853)
);

INVxp33_ASAP7_75t_SL g854 ( 
.A(n_464),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_589),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_593),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_610),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_613),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_616),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_621),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_445),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_637),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_663),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_667),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_680),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_683),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_684),
.Y(n_867)
);

BUFx2_ASAP7_75t_SL g868 ( 
.A(n_447),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_448),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_452),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_456),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_726),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_664),
.Y(n_874)
);

CKINVDCx14_ASAP7_75t_R g875 ( 
.A(n_450),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_505),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_509),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_552),
.Y(n_878)
);

INVxp33_ASAP7_75t_L g879 ( 
.A(n_731),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_745),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_751),
.B(n_1),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_756),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_757),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_454),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_509),
.Y(n_885)
);

CKINVDCx14_ASAP7_75t_R g886 ( 
.A(n_450),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_766),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_770),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_773),
.Y(n_889)
);

INVxp33_ASAP7_75t_SL g890 ( 
.A(n_465),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_518),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_778),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_783),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_518),
.Y(n_894)
);

BUFx2_ASAP7_75t_SL g895 ( 
.A(n_447),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_576),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_576),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_461),
.Y(n_898)
);

CKINVDCx14_ASAP7_75t_R g899 ( 
.A(n_450),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_664),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_646),
.Y(n_901)
);

CKINVDCx16_ASAP7_75t_R g902 ( 
.A(n_645),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_646),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_696),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_696),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_698),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_698),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_664),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_747),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_747),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_493),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_463),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_761),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_481),
.Y(n_914)
);

INVxp33_ASAP7_75t_SL g915 ( 
.A(n_465),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_761),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_639),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_438),
.Y(n_918)
);

INVxp33_ASAP7_75t_SL g919 ( 
.A(n_470),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_441),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_446),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_488),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_468),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_436),
.Y(n_925)
);

INVxp33_ASAP7_75t_SL g926 ( 
.A(n_470),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_471),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_472),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_734),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_490),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_639),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_552),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_475),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_483),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_582),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_491),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_492),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_582),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_734),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_505),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_504),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_520),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_497),
.B(n_3),
.Y(n_943)
);

INVxp33_ASAP7_75t_SL g944 ( 
.A(n_478),
.Y(n_944)
);

INVxp33_ASAP7_75t_SL g945 ( 
.A(n_478),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_740),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_523),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_494),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_533),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_534),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_544),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_740),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_550),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_617),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_553),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_562),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_563),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_569),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_588),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_602),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_740),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_604),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_505),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_495),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_614),
.Y(n_965)
);

INVxp33_ASAP7_75t_L g966 ( 
.A(n_541),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_505),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_615),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_502),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_541),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_619),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_769),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_624),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_631),
.Y(n_974)
);

CKINVDCx14_ASAP7_75t_R g975 ( 
.A(n_546),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_769),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_642),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_649),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_782),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_660),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_617),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_666),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_669),
.Y(n_983)
);

CKINVDCx16_ASAP7_75t_R g984 ( 
.A(n_699),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_715),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_670),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_690),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_691),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_546),
.Y(n_989)
);

INVxp33_ASAP7_75t_L g990 ( 
.A(n_715),
.Y(n_990)
);

CKINVDCx16_ASAP7_75t_R g991 ( 
.A(n_514),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_700),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_729),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_733),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_503),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_739),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_741),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_748),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_758),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_760),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_763),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_764),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_772),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_777),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_514),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_735),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_623),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_735),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_776),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_776),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_497),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_525),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_771),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_525),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_568),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_568),
.Y(n_1016)
);

CKINVDCx14_ASAP7_75t_R g1017 ( 
.A(n_546),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_608),
.Y(n_1018)
);

INVxp67_ASAP7_75t_SL g1019 ( 
.A(n_705),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_746),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_623),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_608),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_620),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_620),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_651),
.Y(n_1025)
);

CKINVDCx14_ASAP7_75t_R g1026 ( 
.A(n_591),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_771),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_513),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_651),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_774),
.Y(n_1030)
);

INVxp33_ASAP7_75t_L g1031 ( 
.A(n_507),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_657),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_657),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_591),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_774),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_591),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_629),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_728),
.Y(n_1038)
);

INVxp33_ASAP7_75t_SL g1039 ( 
.A(n_779),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_629),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_469),
.B(n_3),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_437),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_782),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_440),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_759),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_444),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_728),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_451),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_517),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_779),
.Y(n_1050)
);

CKINVDCx14_ASAP7_75t_R g1051 ( 
.A(n_728),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_515),
.Y(n_1052)
);

CKINVDCx16_ASAP7_75t_R g1053 ( 
.A(n_515),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_453),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_519),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_455),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_524),
.Y(n_1057)
);

INVxp33_ASAP7_75t_SL g1058 ( 
.A(n_780),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_574),
.B(n_5),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_526),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_459),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_647),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_482),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_462),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_647),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_736),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_811),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_785),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_989),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_813),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_799),
.Y(n_1071)
);

BUFx8_ASAP7_75t_SL g1072 ( 
.A(n_826),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_816),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_972),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_894),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_817),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_799),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_791),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_799),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_953),
.B(n_473),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_809),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1013),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_809),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_809),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_796),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_991),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_797),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_809),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_917),
.Y(n_1089)
);

BUFx8_ASAP7_75t_L g1090 ( 
.A(n_1036),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_993),
.B(n_473),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_917),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_989),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_810),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_917),
.Y(n_1095)
);

INVx6_ASAP7_75t_L g1096 ( 
.A(n_1018),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_931),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_931),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1034),
.B(n_650),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_896),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_788),
.A2(n_528),
.B(n_527),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_970),
.A2(n_477),
.B(n_474),
.Y(n_1102)
);

BUFx8_ASAP7_75t_SL g1103 ( 
.A(n_826),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_798),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_966),
.B(n_474),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_931),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_879),
.A2(n_727),
.B1(n_743),
.B2(n_721),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_788),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_851),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_784),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_1018),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_972),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_789),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_851),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_812),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_786),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1018),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1018),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_838),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_970),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_879),
.B(n_736),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1034),
.B(n_579),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_985),
.A2(n_775),
.B(n_477),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_985),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_840),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_805),
.B(n_736),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_966),
.B(n_775),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_790),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_805),
.B(n_762),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_918),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_861),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_990),
.B(n_781),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_792),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_869),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_793),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_794),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_820),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_847),
.A2(n_535),
.B(n_530),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_871),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_821),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_818),
.B(n_762),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1047),
.B(n_877),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_822),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_884),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_814),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_825),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_819),
.A2(n_727),
.B1(n_743),
.B2(n_721),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_827),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_828),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_847),
.A2(n_538),
.B(n_536),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_920),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_823),
.Y(n_1152)
);

BUFx8_ASAP7_75t_SL g1153 ( 
.A(n_833),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_990),
.B(n_781),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_897),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_898),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1041),
.A2(n_754),
.B1(n_521),
.B2(n_597),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1063),
.B(n_605),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1027),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_921),
.B(n_539),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_912),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_830),
.Y(n_1162)
);

BUFx8_ASAP7_75t_SL g1163 ( 
.A(n_833),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_923),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_876),
.B(n_665),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_1005),
.B(n_708),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1035),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1047),
.B(n_668),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_927),
.Y(n_1169)
);

BUFx8_ASAP7_75t_SL g1170 ( 
.A(n_878),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_928),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_832),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_834),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_914),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_922),
.Y(n_1175)
);

INVx6_ASAP7_75t_L g1176 ( 
.A(n_881),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_835),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_976),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_885),
.B(n_540),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_930),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_836),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1042),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_948),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_842),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_878),
.A2(n_754),
.B1(n_954),
.B2(n_932),
.Y(n_1185)
);

INVx6_ASAP7_75t_L g1186 ( 
.A(n_824),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_845),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_933),
.Y(n_1188)
);

CKINVDCx6p67_ASAP7_75t_R g1189 ( 
.A(n_787),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_846),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1036),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_934),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_964),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_969),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_849),
.Y(n_1195)
);

BUFx8_ASAP7_75t_SL g1196 ( 
.A(n_932),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_936),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_901),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_850),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1059),
.A2(n_516),
.B1(n_567),
.B2(n_566),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_937),
.B(n_542),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_852),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_995),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_941),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_942),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1028),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_947),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_853),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_949),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1055),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_855),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_950),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1057),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_940),
.A2(n_548),
.B(n_545),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_856),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_858),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_891),
.B(n_549),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_951),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1060),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_955),
.B(n_551),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_979),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_859),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_956),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_954),
.A2(n_780),
.B1(n_611),
.B2(n_641),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_860),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_818),
.B(n_762),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_943),
.B(n_486),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1006),
.A2(n_557),
.B(n_555),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_957),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_875),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_958),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_862),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1059),
.A2(n_516),
.B1(n_567),
.B2(n_566),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_959),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_905),
.B(n_561),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_L g1237 ( 
.A(n_1044),
.B(n_592),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_1038),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_960),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_863),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_864),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1030),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1108),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1117),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1117),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1237),
.A2(n_857),
.B1(n_844),
.B2(n_808),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1122),
.B(n_1031),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1158),
.B(n_925),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1130),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1071),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1110),
.Y(n_1251)
);

AND2x6_ASAP7_75t_L g1252 ( 
.A(n_1126),
.B(n_943),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1121),
.B(n_1031),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1128),
.A2(n_1009),
.B(n_1008),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1010),
.B(n_965),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1200),
.A2(n_1007),
.B1(n_1021),
.B2(n_981),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1113),
.B(n_875),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1120),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1151),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1113),
.B(n_886),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1133),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1133),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1164),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1071),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1133),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1135),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1145),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_L g1269 ( 
.A(n_1165),
.B(n_592),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1145),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1152),
.B(n_886),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1169),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1135),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1171),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1188),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1135),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1152),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

AND2x6_ASAP7_75t_L g1279 ( 
.A(n_1129),
.B(n_1066),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1192),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1136),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1197),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1105),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1136),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1204),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1071),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1067),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1077),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1205),
.Y(n_1289)
);

AND2x6_ASAP7_75t_L g1290 ( 
.A(n_1141),
.B(n_1066),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1105),
.B(n_899),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1207),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1210),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1158),
.B(n_899),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1079),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1081),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1081),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1213),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1083),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1228),
.A2(n_815),
.B1(n_843),
.B2(n_795),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1186),
.B(n_868),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1081),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1228),
.B(n_848),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1219),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1224),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1097),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1230),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1084),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1084),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1127),
.B(n_975),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1127),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1232),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1235),
.Y(n_1313)
);

XNOR2xp5_ASAP7_75t_L g1314 ( 
.A(n_1200),
.B(n_981),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1239),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1074),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1089),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1074),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1096),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1106),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1089),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1096),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1096),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1165),
.B(n_975),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1085),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1150),
.A2(n_968),
.B(n_962),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1132),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1087),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1089),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1104),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1112),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1165),
.B(n_1142),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1137),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1137),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1070),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1092),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1122),
.B(n_831),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1073),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1140),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1076),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1165),
.B(n_1017),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1132),
.B(n_1154),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1092),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1092),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1098),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1098),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1168),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1140),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1098),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1176),
.A2(n_841),
.B1(n_902),
.B2(n_839),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1170),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1140),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1146),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1088),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1154),
.B(n_1017),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1178),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1111),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1088),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1111),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1146),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1178),
.B(n_1026),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1146),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1148),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1222),
.B(n_1026),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1142),
.B(n_800),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1101),
.A2(n_967),
.B(n_963),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1111),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1148),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1069),
.B(n_802),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1148),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1182),
.B(n_1051),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1149),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1118),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1118),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1149),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1149),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1179),
.B(n_1051),
.Y(n_1378)
);

XNOR2xp5_ASAP7_75t_L g1379 ( 
.A(n_1234),
.B(n_1007),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1118),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1215),
.A2(n_973),
.B(n_971),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1179),
.B(n_974),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1162),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1095),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1075),
.B(n_1011),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1168),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1222),
.B(n_984),
.Y(n_1387)
);

XOR2xp5_ASAP7_75t_L g1388 ( 
.A(n_1086),
.B(n_1052),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1093),
.B(n_803),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1072),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1218),
.B(n_977),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1162),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1242),
.B(n_1043),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1102),
.B(n_1123),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1112),
.B(n_1062),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1095),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1242),
.B(n_1227),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1162),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1090),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1218),
.B(n_978),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1143),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1255),
.Y(n_1402)
);

AND2x6_ASAP7_75t_L g1403 ( 
.A(n_1343),
.B(n_1099),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1332),
.A2(n_1201),
.B(n_1160),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1268),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1249),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1255),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1260),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1264),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1303),
.B(n_1234),
.C(n_1091),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1243),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1272),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1277),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1243),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1303),
.A2(n_1157),
.B1(n_1229),
.B2(n_1225),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1283),
.B(n_1099),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1270),
.B(n_1254),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1274),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1275),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1283),
.B(n_1236),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1257),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1352),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1280),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1262),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1311),
.B(n_1236),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1259),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1311),
.B(n_1080),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1282),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1285),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1352),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1252),
.A2(n_1157),
.B1(n_1229),
.B2(n_1225),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1289),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1292),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1327),
.B(n_1080),
.Y(n_1436)
);

INVxp33_ASAP7_75t_L g1437 ( 
.A(n_1270),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1293),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1298),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1385),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1385),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1259),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1288),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.B(n_1348),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1304),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1288),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1386),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1327),
.B(n_1156),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1295),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1305),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1366),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1307),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1252),
.B(n_1091),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1344),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1295),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1299),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1370),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1312),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1299),
.Y(n_1459)
);

NOR2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1294),
.B(n_1231),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1306),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_L g1462 ( 
.A(n_1337),
.B(n_1053),
.C(n_1107),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1306),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1320),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1313),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1315),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1397),
.B(n_1394),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1366),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1252),
.A2(n_1167),
.B1(n_1082),
.B2(n_1176),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1401),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_SL g1471 ( 
.A(n_1301),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1401),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1248),
.B(n_1082),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1325),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1320),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1300),
.B(n_1167),
.C(n_1048),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1252),
.B(n_1160),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1279),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1251),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1251),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1358),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1394),
.B(n_1180),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1250),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1253),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1328),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1279),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1253),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1330),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1355),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1355),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1388),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1291),
.B(n_1183),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1359),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1247),
.B(n_1094),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1359),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1324),
.B(n_606),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1396),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1396),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1335),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1287),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1287),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1335),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1338),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1338),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1310),
.B(n_1203),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1341),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1252),
.B(n_1201),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1370),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1341),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1279),
.B(n_1221),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1344),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1389),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1279),
.B(n_1221),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1389),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1279),
.B(n_1094),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1244),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1384),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1262),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1245),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1301),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1384),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1346),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1263),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_1316),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1269),
.A2(n_1176),
.B1(n_1214),
.B2(n_618),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1266),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1269),
.B(n_1054),
.C(n_1046),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1319),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1400),
.A2(n_1147),
.B1(n_1159),
.B2(n_1144),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1326),
.A2(n_829),
.B1(n_872),
.B2(n_1102),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1322),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1266),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_L g1534 ( 
.A(n_1290),
.B(n_606),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1382),
.A2(n_801),
.B(n_1012),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1267),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1314),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1290),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1342),
.B(n_618),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1356),
.B(n_1134),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1323),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1346),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1391),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1247),
.B(n_1134),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1267),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1350),
.Y(n_1546)
);

INVxp33_ASAP7_75t_SL g1547 ( 
.A(n_1351),
.Y(n_1547)
);

INVxp33_ASAP7_75t_SL g1548 ( 
.A(n_1258),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1350),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1273),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1273),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1412),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1405),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1429),
.B(n_1261),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1443),
.Y(n_1555)
);

BUFx4f_ASAP7_75t_L g1556 ( 
.A(n_1414),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1412),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1473),
.B(n_895),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1426),
.B(n_1301),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1415),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1410),
.A2(n_1378),
.B1(n_1357),
.B2(n_1246),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1436),
.B(n_1473),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1415),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1418),
.B(n_1393),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1403),
.A2(n_1290),
.B1(n_1337),
.B2(n_1387),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1451),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1428),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1428),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1442),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1437),
.B(n_1357),
.Y(n_1570)
);

BUFx10_ASAP7_75t_L g1571 ( 
.A(n_1471),
.Y(n_1571)
);

INVx5_ASAP7_75t_L g1572 ( 
.A(n_1481),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1451),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1468),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1468),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1443),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1481),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1437),
.B(n_1271),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1290),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1481),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1551),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1448),
.B(n_1115),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1421),
.B(n_1290),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1479),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1403),
.B(n_1144),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1448),
.B(n_1119),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1454),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1446),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1480),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1480),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1481),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1484),
.Y(n_1594)
);

OAI22x1_ASAP7_75t_SL g1595 ( 
.A1(n_1422),
.A2(n_1021),
.B1(n_1040),
.B2(n_1037),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1484),
.Y(n_1596)
);

INVx4_ASAP7_75t_SL g1597 ( 
.A(n_1471),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1487),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1426),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1525),
.B(n_1362),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1454),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1457),
.B(n_1399),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1487),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1440),
.B(n_1333),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1525),
.B(n_1125),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1500),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1489),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1446),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1489),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1548),
.B(n_1494),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1444),
.B(n_1365),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1490),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1490),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1441),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1548),
.B(n_1131),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1423),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1449),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1493),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1511),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1455),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1513),
.B(n_1318),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1547),
.A2(n_1166),
.B1(n_1185),
.B2(n_1107),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1447),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1441),
.B(n_1339),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1508),
.B(n_1331),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1432),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1529),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1455),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1512),
.B(n_1340),
.Y(n_1630)
);

BUFx4f_ASAP7_75t_L g1631 ( 
.A(n_1403),
.Y(n_1631)
);

AO22x2_ASAP7_75t_L g1632 ( 
.A1(n_1462),
.A2(n_1379),
.B1(n_1185),
.B2(n_874),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1515),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_L g1634 ( 
.A(n_1403),
.B(n_1516),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1403),
.B(n_1161),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1417),
.B(n_1161),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1526),
.B(n_1331),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1456),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1416),
.A2(n_1147),
.B1(n_1020),
.B2(n_1045),
.C(n_1019),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1532),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1521),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1456),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1494),
.B(n_1175),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1493),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1483),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_1544),
.Y(n_1646)
);

AND2x6_ASAP7_75t_L g1647 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1417),
.B(n_1175),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1495),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1506),
.B(n_1194),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1478),
.Y(n_1651)
);

NOR2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1476),
.B(n_1189),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1495),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1544),
.B(n_1139),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1491),
.Y(n_1655)
);

NAND2x1p5_ASAP7_75t_L g1656 ( 
.A(n_1478),
.B(n_1194),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1483),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1486),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1406),
.B(n_1349),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1496),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1459),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1496),
.Y(n_1662)
);

AND2x6_ASAP7_75t_SL g1663 ( 
.A(n_1583),
.B(n_1072),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1610),
.B(n_1453),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1645),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1578),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1553),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1646),
.B(n_1477),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1607),
.Y(n_1669)
);

INVx8_ASAP7_75t_L g1670 ( 
.A(n_1572),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1607),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1609),
.Y(n_1672)
);

AND2x2_ASAP7_75t_SL g1673 ( 
.A(n_1654),
.B(n_1534),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1646),
.B(n_1507),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1558),
.B(n_1040),
.C(n_1037),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1562),
.B(n_1416),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1564),
.B(n_1427),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1554),
.B(n_1427),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1609),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1613),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1637),
.B(n_1530),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1613),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1636),
.B(n_1433),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1634),
.A2(n_1534),
.B(n_1483),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1639),
.A2(n_1433),
.B1(n_1531),
.B2(n_1467),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1559),
.B(n_1408),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1570),
.B(n_1492),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1587),
.B(n_1469),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1627),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1612),
.B(n_1159),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1616),
.B(n_1492),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1614),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1614),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1619),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1619),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1648),
.B(n_1409),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1561),
.A2(n_1539),
.B1(n_1540),
.B2(n_1505),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1413),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1580),
.B(n_1510),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1647),
.B(n_1419),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1647),
.B(n_1420),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1623),
.A2(n_1531),
.B1(n_1467),
.B2(n_1404),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1565),
.A2(n_1539),
.B1(n_1540),
.B2(n_1643),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1556),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1584),
.A2(n_1528),
.B(n_1514),
.C(n_1424),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1622),
.B(n_1505),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1631),
.B(n_1482),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1605),
.B(n_1211),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1660),
.A2(n_1482),
.B1(n_1404),
.B2(n_1431),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1578),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1647),
.B(n_1430),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1647),
.B(n_1434),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1631),
.A2(n_1538),
.B1(n_1486),
.B2(n_1438),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1556),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_SL g1716 ( 
.A1(n_1574),
.A2(n_1509),
.B(n_1506),
.C(n_1502),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_SL g1717 ( 
.A(n_1617),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1599),
.B(n_1206),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1579),
.B(n_1435),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1644),
.Y(n_1720)
);

AND2x6_ASAP7_75t_L g1721 ( 
.A(n_1651),
.B(n_1538),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1626),
.B(n_1439),
.Y(n_1722)
);

NOR2xp67_ASAP7_75t_SL g1723 ( 
.A(n_1572),
.B(n_1174),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1600),
.B(n_1445),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1599),
.B(n_1206),
.Y(n_1725)
);

AO22x1_ASAP7_75t_L g1726 ( 
.A1(n_1559),
.A2(n_929),
.B1(n_961),
.B2(n_900),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1659),
.B(n_1450),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1624),
.B(n_1220),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1572),
.B(n_1509),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1682),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1687),
.B(n_1662),
.Y(n_1731)
);

AND2x6_ASAP7_75t_L g1732 ( 
.A(n_1665),
.B(n_1651),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1692),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1693),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1670),
.Y(n_1735)
);

BUFx4f_ASAP7_75t_L g1736 ( 
.A(n_1670),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1670),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1694),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1691),
.B(n_1566),
.Y(n_1739)
);

BUFx12f_ASAP7_75t_L g1740 ( 
.A(n_1689),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1676),
.B(n_1683),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1669),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1721),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1667),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1728),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1687),
.B(n_1599),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1691),
.B(n_1566),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1681),
.B(n_1677),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1671),
.Y(n_1749)
);

AND2x4_ASAP7_75t_SL g1750 ( 
.A(n_1686),
.B(n_1571),
.Y(n_1750)
);

INVx3_ASAP7_75t_SL g1751 ( 
.A(n_1717),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1672),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1679),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1663),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1680),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1695),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1686),
.B(n_1651),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1696),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1705),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1720),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1727),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1709),
.B(n_1566),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1681),
.B(n_1615),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1721),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1666),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1709),
.B(n_1065),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1719),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1721),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1711),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1690),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1701),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1673),
.A2(n_1632),
.B1(n_1422),
.B2(n_1628),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1537),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1745),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1748),
.A2(n_1664),
.B(n_1684),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1730),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1774),
.A2(n_1673),
.B1(n_1685),
.B2(n_1707),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1772),
.B(n_1707),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1769),
.A2(n_1664),
.B(n_1685),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1764),
.B(n_1632),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1769),
.A2(n_1708),
.B(n_1688),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1731),
.B(n_1724),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1768),
.B(n_1678),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1741),
.B(n_1722),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_SL g1787 ( 
.A1(n_1755),
.A2(n_1723),
.B(n_1698),
.C(n_1704),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1739),
.A2(n_1675),
.B(n_1535),
.C(n_1674),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1749),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1655),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1769),
.A2(n_1708),
.B(n_1706),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1747),
.A2(n_1635),
.B(n_1586),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1746),
.A2(n_1700),
.B(n_1697),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1763),
.A2(n_1710),
.B(n_1703),
.C(n_1699),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1773),
.A2(n_1703),
.B(n_1668),
.C(n_1674),
.Y(n_1797)
);

XOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1754),
.B(n_1491),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1741),
.B(n_1726),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1773),
.A2(n_1700),
.B(n_1668),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_SL g1801 ( 
.A1(n_1755),
.A2(n_1714),
.B(n_1712),
.C(n_1713),
.Y(n_1801)
);

BUFx4f_ASAP7_75t_L g1802 ( 
.A(n_1751),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1751),
.B(n_1615),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1755),
.A2(n_1716),
.B(n_1657),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1736),
.A2(n_1715),
.B1(n_1640),
.B2(n_1656),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1744),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_SL g1807 ( 
.A(n_1740),
.B(n_1390),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1736),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1765),
.A2(n_1716),
.B(n_1657),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1742),
.A2(n_1038),
.B(n_1725),
.C(n_1718),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1740),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1752),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1733),
.A2(n_1702),
.B(n_1652),
.C(n_1458),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1735),
.B(n_1602),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1765),
.A2(n_1645),
.B(n_1729),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1759),
.A2(n_1367),
.B(n_1567),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1733),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_SL g1818 ( 
.A1(n_1765),
.A2(n_1665),
.B(n_1061),
.C(n_1064),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1758),
.B(n_1633),
.Y(n_1819)
);

INVx8_ASAP7_75t_L g1820 ( 
.A(n_1732),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1808),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1802),
.Y(n_1822)
);

BUFx12f_ASAP7_75t_L g1823 ( 
.A(n_1811),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1793),
.B(n_1766),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1766),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1802),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1771),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1817),
.Y(n_1828)
);

OR2x6_ASAP7_75t_L g1829 ( 
.A(n_1820),
.B(n_1770),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1778),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1800),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1808),
.B(n_1814),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1808),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1779),
.A2(n_1065),
.B1(n_1738),
.B2(n_1734),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1775),
.B(n_1537),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1784),
.B(n_1771),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1797),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1820),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1806),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1776),
.Y(n_1842)
);

AOI21x1_ASAP7_75t_L g1843 ( 
.A1(n_1804),
.A2(n_1738),
.B(n_1729),
.Y(n_1843)
);

OAI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1796),
.A2(n_1759),
.B(n_1756),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1820),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1790),
.B(n_1758),
.Y(n_1846)
);

INVx8_ASAP7_75t_L g1847 ( 
.A(n_1780),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1791),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1785),
.B(n_1752),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1799),
.B(n_1753),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1819),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1812),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1781),
.A2(n_1103),
.B1(n_1163),
.B2(n_1153),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1813),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1803),
.B(n_1761),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1783),
.B(n_1615),
.Y(n_1856)
);

INVx4_ASAP7_75t_L g1857 ( 
.A(n_1807),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1816),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1815),
.B(n_1758),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1807),
.A2(n_1595),
.B1(n_1754),
.B2(n_1193),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1798),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1805),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1777),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1795),
.A2(n_1103),
.B1(n_1163),
.B2(n_1153),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1787),
.B(n_1757),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1788),
.B(n_1757),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1792),
.B(n_1732),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1816),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1810),
.B(n_1573),
.Y(n_1869)
);

INVx5_ASAP7_75t_L g1870 ( 
.A(n_1818),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1794),
.A2(n_1196),
.B1(n_915),
.B2(n_648),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1809),
.A2(n_1196),
.B1(n_915),
.B2(n_753),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1801),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1842),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1871),
.A2(n_837),
.B(n_1014),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1830),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1825),
.B(n_1750),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1836),
.B(n_1641),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1850),
.Y(n_1879)
);

AO31x2_ASAP7_75t_L g1880 ( 
.A1(n_1858),
.A2(n_1402),
.A3(n_1411),
.B(n_1407),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1822),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_SL g1882 ( 
.A1(n_1835),
.A2(n_625),
.B(n_654),
.C(n_630),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1871),
.A2(n_625),
.B(n_654),
.C(n_630),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1828),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1872),
.A2(n_1191),
.B(n_1090),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1863),
.A2(n_1736),
.B(n_1743),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1848),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1835),
.A2(n_1186),
.B1(n_755),
.B2(n_1743),
.Y(n_1888)
);

NOR2xp67_ASAP7_75t_L g1889 ( 
.A(n_1857),
.B(n_1209),
.Y(n_1889)
);

AOI21x1_ASAP7_75t_L g1890 ( 
.A1(n_1856),
.A2(n_904),
.B(n_903),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1837),
.B(n_480),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1872),
.A2(n_1016),
.B(n_1015),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1822),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1837),
.B(n_1123),
.Y(n_1894)
);

OAI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1857),
.A2(n_1743),
.B1(n_1770),
.B2(n_908),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1853),
.A2(n_755),
.B(n_1023),
.C(n_1022),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1838),
.A2(n_872),
.B(n_829),
.C(n_1024),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_SL g1898 ( 
.A(n_1823),
.B(n_1735),
.Y(n_1898)
);

AO32x2_ASAP7_75t_L g1899 ( 
.A1(n_1862),
.A2(n_1402),
.A3(n_1737),
.B1(n_1735),
.B2(n_919),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1863),
.A2(n_1743),
.B(n_1770),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1840),
.B(n_911),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1822),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1831),
.A2(n_1770),
.B(n_1519),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1831),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1840),
.B(n_854),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1832),
.Y(n_1906)
);

O2A1O1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1838),
.A2(n_1029),
.B(n_1032),
.C(n_1025),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1843),
.A2(n_1569),
.B(n_1568),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1852),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1861),
.B(n_1760),
.Y(n_1910)
);

AO32x2_ASAP7_75t_L g1911 ( 
.A1(n_1841),
.A2(n_1402),
.A3(n_1737),
.B1(n_944),
.B2(n_945),
.Y(n_1911)
);

AO32x2_ASAP7_75t_L g1912 ( 
.A1(n_1826),
.A2(n_1737),
.A3(n_1039),
.B1(n_1058),
.B2(n_926),
.Y(n_1912)
);

A2O1A1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1853),
.A2(n_1033),
.B(n_1460),
.C(n_1750),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1867),
.A2(n_1770),
.B(n_1425),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1854),
.A2(n_939),
.B(n_924),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1864),
.A2(n_907),
.B(n_909),
.C(n_906),
.Y(n_1916)
);

BUFx12f_ASAP7_75t_L g1917 ( 
.A(n_1833),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1851),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1867),
.A2(n_1411),
.B(n_1578),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1849),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1864),
.A2(n_1860),
.B1(n_952),
.B2(n_946),
.C(n_1844),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1847),
.B(n_1760),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1866),
.B(n_890),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1849),
.B(n_496),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1869),
.A2(n_1593),
.B(n_1581),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1855),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1824),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1846),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1846),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1847),
.A2(n_1602),
.B1(n_1575),
.B2(n_1576),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1824),
.B(n_911),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1865),
.A2(n_1050),
.B(n_938),
.C(n_935),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1833),
.B(n_1573),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1827),
.B(n_935),
.Y(n_1934)
);

AO31x2_ASAP7_75t_L g1935 ( 
.A1(n_1868),
.A2(n_1653),
.A3(n_1649),
.B(n_1557),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1847),
.A2(n_1191),
.B1(n_1238),
.B2(n_1186),
.Y(n_1936)
);

AO32x2_ASAP7_75t_L g1937 ( 
.A1(n_1873),
.A2(n_7),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1827),
.Y(n_1938)
);

AO31x2_ASAP7_75t_L g1939 ( 
.A1(n_1869),
.A2(n_1870),
.A3(n_1873),
.B(n_1653),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1859),
.Y(n_1940)
);

AO21x1_ASAP7_75t_L g1941 ( 
.A1(n_1859),
.A2(n_913),
.B(n_910),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1839),
.B(n_1829),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1821),
.Y(n_1943)
);

NOR2xp67_ASAP7_75t_L g1944 ( 
.A(n_1821),
.B(n_804),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1870),
.A2(n_1503),
.B(n_1499),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1904),
.B(n_1873),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1940),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1884),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1888),
.A2(n_1829),
.B1(n_1870),
.B2(n_1834),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1885),
.A2(n_1870),
.B1(n_1845),
.B2(n_1238),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1879),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1876),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1882),
.A2(n_512),
.B1(n_522),
.B2(n_508),
.C(n_501),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1906),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1921),
.A2(n_1845),
.B1(n_1834),
.B2(n_1829),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1927),
.Y(n_1956)
);

INVx6_ASAP7_75t_L g1957 ( 
.A(n_1917),
.Y(n_1957)
);

BUFx2_ASAP7_75t_R g1958 ( 
.A(n_1887),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1920),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1909),
.Y(n_1960)
);

OAI22xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1923),
.A2(n_531),
.B1(n_532),
.B2(n_529),
.Y(n_1961)
);

OAI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1918),
.A2(n_1845),
.B1(n_1575),
.B2(n_1576),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1903),
.A2(n_1504),
.B(n_1604),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1915),
.A2(n_1918),
.B1(n_1941),
.B2(n_1878),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1880),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1931),
.A2(n_866),
.B1(n_867),
.B2(n_865),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1934),
.A2(n_873),
.B1(n_880),
.B2(n_870),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1926),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1938),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_SL g1970 ( 
.A1(n_1898),
.A2(n_1945),
.B1(n_1875),
.B2(n_1891),
.Y(n_1970)
);

OAI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1883),
.A2(n_558),
.B(n_564),
.C(n_543),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1939),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1935),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1910),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1942),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1880),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1935),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1899),
.B(n_882),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1943),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1905),
.A2(n_887),
.B1(n_888),
.B2(n_883),
.Y(n_1980)
);

A2O1A1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1896),
.A2(n_577),
.B(n_583),
.C(n_565),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1939),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1895),
.A2(n_892),
.B1(n_893),
.B2(n_889),
.Y(n_1983)
);

CKINVDCx8_ASAP7_75t_R g1984 ( 
.A(n_1922),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1901),
.B(n_938),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1874),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1894),
.B(n_980),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1935),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1939),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1908),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1937),
.A2(n_1732),
.B1(n_1068),
.B2(n_586),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1937),
.Y(n_1992)
);

INVx4_ASAP7_75t_L g1993 ( 
.A(n_1881),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1899),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1924),
.B(n_982),
.Y(n_1995)
);

OAI221xp5_ASAP7_75t_L g1996 ( 
.A1(n_1913),
.A2(n_599),
.B1(n_600),
.B2(n_590),
.C(n_584),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1982),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1947),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1951),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1947),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1948),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1959),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1954),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1959),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1960),
.Y(n_2005)
);

OAI21x1_ASAP7_75t_L g2006 ( 
.A1(n_1982),
.A2(n_1919),
.B(n_1900),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1968),
.B(n_1886),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1965),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1956),
.B(n_1899),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1956),
.B(n_1877),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1952),
.Y(n_2012)
);

INVx5_ASAP7_75t_L g2013 ( 
.A(n_1982),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1979),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1994),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1979),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1946),
.B(n_1969),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_SL g2018 ( 
.A1(n_1991),
.A2(n_1970),
.B1(n_1964),
.B2(n_1986),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_R g2019 ( 
.A(n_1957),
.B(n_1078),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1965),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1994),
.B(n_1928),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_SL g2022 ( 
.A1(n_1949),
.A2(n_1937),
.B1(n_1892),
.B2(n_1902),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1985),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1976),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1984),
.B(n_1889),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1973),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_2022),
.A2(n_1981),
.B(n_1978),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2001),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2011),
.B(n_1975),
.Y(n_2029)
);

NOR4xp25_ASAP7_75t_L g2030 ( 
.A(n_2023),
.B(n_1981),
.C(n_1971),
.D(n_1932),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_2008),
.A2(n_1984),
.B1(n_1992),
.B2(n_1996),
.Y(n_2031)
);

OAI21xp33_ASAP7_75t_SL g2032 ( 
.A1(n_1998),
.A2(n_1978),
.B(n_1946),
.Y(n_2032)
);

O2A1O1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_2018),
.A2(n_1961),
.B(n_1995),
.C(n_1953),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_2018),
.A2(n_1950),
.B1(n_1955),
.B2(n_1957),
.Y(n_2034)
);

AOI21x1_ASAP7_75t_L g2035 ( 
.A1(n_2015),
.A2(n_2000),
.B(n_1972),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_2025),
.A2(n_1957),
.B1(n_1975),
.B2(n_1987),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1998),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1999),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_2010),
.A2(n_1957),
.B1(n_1975),
.B2(n_1963),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_2021),
.Y(n_2040)
);

OAI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2017),
.A2(n_1986),
.B1(n_1974),
.B2(n_1972),
.Y(n_2041)
);

OAI21xp33_ASAP7_75t_L g2042 ( 
.A1(n_2010),
.A2(n_1980),
.B(n_2021),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2012),
.A2(n_1983),
.B1(n_1936),
.B2(n_1967),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2001),
.Y(n_2044)
);

OAI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_2012),
.A2(n_1897),
.B(n_1966),
.C(n_609),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2003),
.B(n_1979),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_2003),
.A2(n_1974),
.B(n_1907),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_2011),
.Y(n_2048)
);

AOI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_2005),
.A2(n_626),
.B1(n_633),
.B2(n_622),
.C(n_601),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2005),
.A2(n_640),
.B1(n_653),
.B2(n_635),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2015),
.Y(n_2051)
);

OAI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_2006),
.A2(n_1944),
.B(n_1914),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2044),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2035),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2040),
.B(n_2002),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_L g2057 ( 
.A(n_2037),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2029),
.B(n_2002),
.Y(n_2058)
);

INVx5_ASAP7_75t_SL g2059 ( 
.A(n_2037),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_2037),
.B(n_2013),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2051),
.Y(n_2061)
);

INVx4_ASAP7_75t_L g2062 ( 
.A(n_2038),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2042),
.B(n_2026),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2046),
.B(n_2039),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2027),
.A2(n_1929),
.B1(n_1930),
.B2(n_687),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2048),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2047),
.B(n_2004),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2032),
.B(n_2002),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2036),
.B(n_2004),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_2033),
.B(n_2019),
.Y(n_2070)
);

INVx2_ASAP7_75t_R g2071 ( 
.A(n_2031),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2052),
.B(n_2007),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2034),
.B(n_2007),
.Y(n_2073)
);

INVx3_ASAP7_75t_L g2074 ( 
.A(n_2041),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2031),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2041),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2030),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2050),
.Y(n_2078)
);

NOR4xp25_ASAP7_75t_SL g2079 ( 
.A(n_2049),
.B(n_2026),
.C(n_1958),
.D(n_2019),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2050),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2043),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2043),
.B(n_2007),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2045),
.B(n_2014),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_2038),
.Y(n_2084)
);

OAI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2077),
.A2(n_1997),
.B1(n_1916),
.B2(n_1893),
.C(n_694),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2071),
.A2(n_1993),
.B1(n_2006),
.B2(n_1989),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2071),
.A2(n_1993),
.B1(n_1989),
.B2(n_1990),
.Y(n_2087)
);

AOI322xp5_ASAP7_75t_L g2088 ( 
.A1(n_2070),
.A2(n_704),
.A3(n_692),
.B1(n_709),
.B2(n_712),
.C1(n_697),
.C2(n_655),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2057),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2073),
.B(n_2014),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2079),
.A2(n_1989),
.B1(n_2013),
.B2(n_2016),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2054),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_2070),
.A2(n_1912),
.B1(n_2013),
.B2(n_1911),
.Y(n_2093)
);

OAI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_2075),
.A2(n_2013),
.B1(n_2016),
.B2(n_1993),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_2084),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_2081),
.A2(n_1990),
.B1(n_2013),
.B2(n_1988),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2074),
.A2(n_2013),
.B1(n_1962),
.B2(n_1997),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2062),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_2066),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_L g2100 ( 
.A(n_2076),
.B(n_718),
.C(n_716),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2073),
.B(n_1912),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2083),
.B(n_1997),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2074),
.A2(n_1997),
.B1(n_1977),
.B2(n_1933),
.Y(n_2103)
);

OAI221xp5_ASAP7_75t_L g2104 ( 
.A1(n_2074),
.A2(n_725),
.B1(n_730),
.B2(n_724),
.C(n_720),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_2078),
.A2(n_2080),
.B1(n_2076),
.B2(n_2065),
.C(n_2067),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2064),
.A2(n_1977),
.B1(n_1925),
.B2(n_2024),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2098),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_2099),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2095),
.B(n_2059),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2095),
.B(n_2082),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2098),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2092),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_2089),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2090),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2102),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2105),
.B(n_2101),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2093),
.B(n_2062),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2100),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2104),
.A2(n_2065),
.B1(n_2082),
.B2(n_2062),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2106),
.B(n_2059),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2087),
.B(n_2059),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2094),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2111),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2107),
.Y(n_2124)
);

NAND3xp33_ASAP7_75t_L g2125 ( 
.A(n_2119),
.B(n_2088),
.C(n_2093),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2116),
.A2(n_2119),
.B1(n_2117),
.B2(n_2108),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2107),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2108),
.Y(n_2128)
);

OAI31xp33_ASAP7_75t_SL g2129 ( 
.A1(n_2120),
.A2(n_2097),
.A3(n_2091),
.B(n_2103),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2110),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_2113),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2130),
.B(n_2114),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2124),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2127),
.Y(n_2134)
);

NAND2x1_ASAP7_75t_L g2135 ( 
.A(n_2131),
.B(n_2109),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2128),
.B(n_2115),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2123),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2125),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2132),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2136),
.B(n_2126),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2133),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2138),
.B(n_2109),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2137),
.B(n_2113),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2142),
.B(n_2140),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_2139),
.B(n_2129),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2143),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_2146),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2144),
.B(n_2135),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_2148),
.B(n_2145),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2147),
.B(n_2134),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2147),
.B(n_2141),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2151),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2149),
.B(n_2125),
.Y(n_2153)
);

OAI321xp33_ASAP7_75t_L g2154 ( 
.A1(n_2153),
.A2(n_2150),
.A3(n_2122),
.B1(n_2113),
.B2(n_2112),
.C(n_2121),
.Y(n_2154)
);

OAI221xp5_ASAP7_75t_L g2155 ( 
.A1(n_2152),
.A2(n_2122),
.B1(n_2118),
.B2(n_2113),
.C(n_2086),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2152),
.B(n_2120),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_2155),
.A2(n_2121),
.B(n_2055),
.C(n_2060),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_2156),
.Y(n_2158)
);

AOI21xp33_ASAP7_75t_L g2159 ( 
.A1(n_2154),
.A2(n_2085),
.B(n_1056),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2156),
.B(n_2055),
.Y(n_2160)
);

NOR2x1_ASAP7_75t_L g2161 ( 
.A(n_2160),
.B(n_806),
.Y(n_2161)
);

NOR3x1_ASAP7_75t_L g2162 ( 
.A(n_2159),
.B(n_1597),
.C(n_1571),
.Y(n_2162)
);

NAND4xp25_ASAP7_75t_L g2163 ( 
.A(n_2158),
.B(n_1597),
.C(n_2096),
.D(n_1177),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_2157),
.A2(n_807),
.B(n_737),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2162),
.B(n_2164),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_2161),
.Y(n_2166)
);

AO22x2_ASAP7_75t_L g2167 ( 
.A1(n_2163),
.A2(n_2053),
.B1(n_2060),
.B2(n_2063),
.Y(n_2167)
);

O2A1O1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2164),
.A2(n_1212),
.B(n_1172),
.C(n_1195),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2162),
.B(n_2057),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2161),
.Y(n_2170)
);

AOI21xp33_ASAP7_75t_L g2171 ( 
.A1(n_2161),
.A2(n_738),
.B(n_732),
.Y(n_2171)
);

NOR3xp33_ASAP7_75t_L g2172 ( 
.A(n_2164),
.B(n_1226),
.C(n_1216),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2161),
.Y(n_2173)
);

A2O1A1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_2164),
.A2(n_2060),
.B(n_2057),
.C(n_2053),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2164),
.A2(n_750),
.B(n_742),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2164),
.A2(n_768),
.B(n_752),
.C(n_1233),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2161),
.B(n_1212),
.Y(n_2177)
);

AOI211x1_ASAP7_75t_L g2178 ( 
.A1(n_2164),
.A2(n_2069),
.B(n_2072),
.C(n_2061),
.Y(n_2178)
);

NOR3xp33_ASAP7_75t_L g2179 ( 
.A(n_2176),
.B(n_2165),
.C(n_2171),
.Y(n_2179)
);

NOR3x1_ASAP7_75t_L g2180 ( 
.A(n_2169),
.B(n_986),
.C(n_983),
.Y(n_2180)
);

NAND3xp33_ASAP7_75t_L g2181 ( 
.A(n_2170),
.B(n_1240),
.C(n_1181),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2175),
.A2(n_988),
.B(n_987),
.Y(n_2182)
);

NAND4xp75_ASAP7_75t_L g2183 ( 
.A(n_2177),
.B(n_1452),
.C(n_1466),
.D(n_1465),
.Y(n_2183)
);

AND5x1_ASAP7_75t_L g2184 ( 
.A(n_2174),
.B(n_1912),
.C(n_2057),
.D(n_9),
.E(n_6),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2167),
.B(n_2072),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2167),
.B(n_2053),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2166),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2173),
.B(n_2068),
.Y(n_2188)
);

AND2x2_ASAP7_75t_SL g2189 ( 
.A(n_2172),
.B(n_1573),
.Y(n_2189)
);

NAND5xp2_ASAP7_75t_L g2190 ( 
.A(n_2168),
.B(n_2178),
.C(n_1485),
.D(n_1488),
.E(n_1474),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_2169),
.B(n_7),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2167),
.B(n_2068),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2167),
.Y(n_2193)
);

NOR2xp67_ASAP7_75t_L g2194 ( 
.A(n_2169),
.B(n_9),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2169),
.B(n_11),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2167),
.B(n_2056),
.Y(n_2196)
);

NOR3x1_ASAP7_75t_L g2197 ( 
.A(n_2169),
.B(n_994),
.C(n_992),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2167),
.Y(n_2198)
);

NOR2x1_ASAP7_75t_L g2199 ( 
.A(n_2177),
.B(n_1100),
.Y(n_2199)
);

NAND2x1_ASAP7_75t_SL g2200 ( 
.A(n_2177),
.B(n_916),
.Y(n_2200)
);

NOR2xp67_ASAP7_75t_L g2201 ( 
.A(n_2169),
.B(n_12),
.Y(n_2201)
);

INVx2_ASAP7_75t_SL g2202 ( 
.A(n_2169),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2169),
.B(n_1173),
.Y(n_2203)
);

NAND4xp25_ASAP7_75t_L g2204 ( 
.A(n_2169),
.B(n_1198),
.C(n_1155),
.D(n_997),
.Y(n_2204)
);

OAI21xp33_ASAP7_75t_L g2205 ( 
.A1(n_2169),
.A2(n_2056),
.B(n_2058),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2169),
.B(n_2058),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2167),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2167),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2167),
.B(n_996),
.Y(n_2209)
);

NOR2x1_ASAP7_75t_L g2210 ( 
.A(n_2177),
.B(n_1109),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2167),
.Y(n_2211)
);

NAND3xp33_ASAP7_75t_SL g2212 ( 
.A(n_2170),
.B(n_571),
.C(n_570),
.Y(n_2212)
);

NAND3xp33_ASAP7_75t_L g2213 ( 
.A(n_2170),
.B(n_1181),
.C(n_1173),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_2169),
.B(n_1173),
.Y(n_2214)
);

NAND4xp25_ASAP7_75t_L g2215 ( 
.A(n_2169),
.B(n_999),
.C(n_1000),
.D(n_998),
.Y(n_2215)
);

NOR2x1_ASAP7_75t_L g2216 ( 
.A(n_2177),
.B(n_1109),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2169),
.B(n_14),
.Y(n_2217)
);

NAND3xp33_ASAP7_75t_L g2218 ( 
.A(n_2170),
.B(n_1184),
.C(n_1181),
.Y(n_2218)
);

XNOR2xp5_ASAP7_75t_L g2219 ( 
.A(n_2169),
.B(n_14),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_SL g2220 ( 
.A(n_2176),
.B(n_1002),
.C(n_1001),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2169),
.B(n_1184),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2167),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_SL g2223 ( 
.A(n_2170),
.B(n_573),
.C(n_572),
.Y(n_2223)
);

NAND4xp25_ASAP7_75t_L g2224 ( 
.A(n_2191),
.B(n_1004),
.C(n_1003),
.D(n_1114),
.Y(n_2224)
);

OA22x2_ASAP7_75t_L g2225 ( 
.A1(n_2219),
.A2(n_1541),
.B1(n_1114),
.B2(n_1630),
.Y(n_2225)
);

AOI21xp33_ASAP7_75t_L g2226 ( 
.A1(n_2193),
.A2(n_1187),
.B(n_1184),
.Y(n_2226)
);

NOR2x1_ASAP7_75t_L g2227 ( 
.A(n_2194),
.B(n_1187),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2188),
.A2(n_1190),
.B1(n_1199),
.B2(n_1187),
.Y(n_2228)
);

NAND4xp75_ASAP7_75t_L g2229 ( 
.A(n_2201),
.B(n_17),
.C(n_15),
.D(n_16),
.Y(n_2229)
);

OAI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2184),
.A2(n_1576),
.B1(n_1575),
.B2(n_1202),
.C(n_1208),
.Y(n_2230)
);

AOI211x1_ASAP7_75t_L g2231 ( 
.A1(n_2186),
.A2(n_1890),
.B(n_23),
.C(n_18),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2192),
.A2(n_1199),
.B1(n_1202),
.B2(n_1190),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_2185),
.B(n_2206),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2196),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2217),
.A2(n_1199),
.B1(n_1202),
.B2(n_1190),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2195),
.A2(n_1217),
.B1(n_1223),
.B2(n_1208),
.Y(n_2236)
);

AOI322xp5_ASAP7_75t_L g2237 ( 
.A1(n_2187),
.A2(n_2024),
.A3(n_2020),
.B1(n_2009),
.B2(n_26),
.C1(n_27),
.C2(n_28),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2198),
.Y(n_2238)
);

NOR3x1_ASAP7_75t_L g2239 ( 
.A(n_2202),
.B(n_18),
.C(n_22),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2205),
.A2(n_1217),
.B1(n_1223),
.B2(n_1208),
.Y(n_2240)
);

OAI211xp5_ASAP7_75t_L g2241 ( 
.A1(n_2207),
.A2(n_1223),
.B(n_1241),
.C(n_1217),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2208),
.A2(n_1241),
.B1(n_2020),
.B2(n_2009),
.Y(n_2242)
);

AOI211xp5_ASAP7_75t_L g2243 ( 
.A1(n_2211),
.A2(n_1241),
.B(n_29),
.C(n_23),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2200),
.Y(n_2244)
);

AOI211xp5_ASAP7_75t_SL g2245 ( 
.A1(n_2222),
.A2(n_1630),
.B(n_1659),
.C(n_30),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2179),
.A2(n_2189),
.B1(n_2223),
.B2(n_2212),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2190),
.B(n_27),
.Y(n_2247)
);

AOI322xp5_ASAP7_75t_L g2248 ( 
.A1(n_2199),
.A2(n_2024),
.A3(n_2020),
.B1(n_2009),
.B2(n_35),
.C1(n_37),
.C2(n_38),
.Y(n_2248)
);

INVxp33_ASAP7_75t_SL g2249 ( 
.A(n_2210),
.Y(n_2249)
);

NAND4xp25_ASAP7_75t_L g2250 ( 
.A(n_2180),
.B(n_33),
.C(n_29),
.D(n_32),
.Y(n_2250)
);

OAI21xp33_ASAP7_75t_L g2251 ( 
.A1(n_2209),
.A2(n_578),
.B(n_575),
.Y(n_2251)
);

OAI221xp5_ASAP7_75t_L g2252 ( 
.A1(n_2216),
.A2(n_595),
.B1(n_596),
.B2(n_594),
.C(n_585),
.Y(n_2252)
);

OAI211xp5_ASAP7_75t_L g2253 ( 
.A1(n_2203),
.A2(n_41),
.B(n_37),
.C(n_39),
.Y(n_2253)
);

CKINVDCx16_ASAP7_75t_R g2254 ( 
.A(n_2197),
.Y(n_2254)
);

OAI211xp5_ASAP7_75t_L g2255 ( 
.A1(n_2214),
.A2(n_48),
.B(n_45),
.C(n_46),
.Y(n_2255)
);

AOI31xp33_ASAP7_75t_L g2256 ( 
.A1(n_2213),
.A2(n_603),
.A3(n_607),
.B(n_598),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_2220),
.Y(n_2257)
);

AOI21xp33_ASAP7_75t_L g2258 ( 
.A1(n_2181),
.A2(n_2221),
.B(n_2218),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2182),
.B(n_48),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2183),
.Y(n_2260)
);

NOR3xp33_ASAP7_75t_L g2261 ( 
.A(n_2204),
.B(n_1354),
.C(n_1353),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2215),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2192),
.B(n_1911),
.Y(n_2263)
);

AO22x2_ASAP7_75t_L g2264 ( 
.A1(n_2193),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2264)
);

AOI221xp5_ASAP7_75t_L g2265 ( 
.A1(n_2193),
.A2(n_632),
.B1(n_636),
.B2(n_628),
.C(n_627),
.Y(n_2265)
);

OAI221xp5_ASAP7_75t_SL g2266 ( 
.A1(n_2188),
.A2(n_54),
.B1(n_50),
.B2(n_51),
.C(n_55),
.Y(n_2266)
);

AOI221x1_ASAP7_75t_L g2267 ( 
.A1(n_2193),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_2267)
);

OAI221xp5_ASAP7_75t_L g2268 ( 
.A1(n_2184),
.A2(n_652),
.B1(n_659),
.B2(n_644),
.C(n_643),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2186),
.Y(n_2269)
);

AO22x2_ASAP7_75t_L g2270 ( 
.A1(n_2193),
.A2(n_60),
.B1(n_56),
.B2(n_58),
.Y(n_2270)
);

NOR3xp33_ASAP7_75t_L g2271 ( 
.A(n_2191),
.B(n_1363),
.C(n_1361),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_2194),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2188),
.B(n_60),
.Y(n_2273)
);

A2O1A1Ixp33_ASAP7_75t_L g2274 ( 
.A1(n_2191),
.A2(n_68),
.B(n_62),
.C(n_67),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2194),
.B(n_62),
.Y(n_2275)
);

OAI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2186),
.A2(n_1658),
.B1(n_662),
.B2(n_671),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2193),
.A2(n_673),
.B(n_661),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2186),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2194),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2186),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_2194),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2186),
.Y(n_2282)
);

NAND4xp75_ASAP7_75t_L g2283 ( 
.A(n_2194),
.B(n_72),
.C(n_67),
.D(n_71),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2191),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2186),
.Y(n_2285)
);

OAI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2194),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_2286)
);

O2A1O1Ixp33_ASAP7_75t_L g2287 ( 
.A1(n_2193),
.A2(n_78),
.B(n_74),
.C(n_76),
.Y(n_2287)
);

AOI211xp5_ASAP7_75t_L g2288 ( 
.A1(n_2194),
.A2(n_79),
.B(n_74),
.C(n_78),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2192),
.A2(n_675),
.B1(n_676),
.B2(n_674),
.Y(n_2289)
);

OA22x2_ASAP7_75t_L g2290 ( 
.A1(n_2219),
.A2(n_87),
.B1(n_80),
.B2(n_85),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2193),
.A2(n_678),
.B(n_677),
.Y(n_2291)
);

AOI211xp5_ASAP7_75t_L g2292 ( 
.A1(n_2194),
.A2(n_90),
.B(n_85),
.C(n_89),
.Y(n_2292)
);

AOI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2193),
.A2(n_685),
.B1(n_686),
.B2(n_682),
.C(n_681),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2192),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.C1(n_94),
.C2(n_95),
.Y(n_2294)
);

OAI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2188),
.A2(n_701),
.B1(n_702),
.B2(n_688),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2193),
.A2(n_707),
.B1(n_710),
.B2(n_706),
.C(n_703),
.Y(n_2296)
);

AOI211xp5_ASAP7_75t_L g2297 ( 
.A1(n_2194),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2285),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2275),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2290),
.Y(n_2300)
);

NOR2x1_ASAP7_75t_L g2301 ( 
.A(n_2229),
.B(n_96),
.Y(n_2301)
);

NOR2x1p5_ASAP7_75t_L g2302 ( 
.A(n_2283),
.B(n_711),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2238),
.A2(n_717),
.B(n_713),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_2239),
.Y(n_2304)
);

NOR3xp33_ASAP7_75t_L g2305 ( 
.A(n_2234),
.B(n_1369),
.C(n_1364),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2273),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_SL g2307 ( 
.A(n_2294),
.B(n_723),
.C(n_722),
.Y(n_2307)
);

NOR3x1_ASAP7_75t_L g2308 ( 
.A(n_2286),
.B(n_97),
.C(n_99),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2269),
.B(n_1373),
.C(n_1371),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2266),
.A2(n_1520),
.B1(n_1517),
.B2(n_1377),
.Y(n_2310)
);

NAND2x1_ASAP7_75t_SL g2311 ( 
.A(n_2275),
.B(n_101),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2250),
.B(n_102),
.Y(n_2312)
);

OAI21xp33_ASAP7_75t_SL g2313 ( 
.A1(n_2227),
.A2(n_102),
.B(n_103),
.Y(n_2313)
);

NOR2x1_ASAP7_75t_L g2314 ( 
.A(n_2230),
.B(n_104),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2233),
.A2(n_1611),
.B1(n_1625),
.B2(n_1604),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2264),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2264),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2272),
.B(n_107),
.Y(n_2318)
);

NAND3xp33_ASAP7_75t_SL g2319 ( 
.A(n_2288),
.B(n_108),
.C(n_110),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2270),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2292),
.B(n_1376),
.Y(n_2321)
);

A2O1A1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2287),
.A2(n_114),
.B(n_110),
.C(n_112),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2279),
.B(n_2281),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2278),
.A2(n_1625),
.B1(n_1611),
.B2(n_1392),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2253),
.A2(n_116),
.B(n_112),
.C(n_115),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2280),
.A2(n_1398),
.B1(n_1383),
.B2(n_1470),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2282),
.A2(n_967),
.B(n_963),
.Y(n_2327)
);

NAND4xp75_ASAP7_75t_L g2328 ( 
.A(n_2267),
.B(n_118),
.C(n_115),
.D(n_117),
.Y(n_2328)
);

NOR3xp33_ASAP7_75t_SL g2329 ( 
.A(n_2254),
.B(n_119),
.C(n_122),
.Y(n_2329)
);

NAND4xp75_ASAP7_75t_L g2330 ( 
.A(n_2260),
.B(n_123),
.C(n_119),
.D(n_122),
.Y(n_2330)
);

NOR4xp75_ASAP7_75t_L g2331 ( 
.A(n_2259),
.B(n_126),
.C(n_123),
.D(n_125),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2270),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2247),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2297),
.B(n_126),
.Y(n_2334)
);

OAI21xp33_ASAP7_75t_L g2335 ( 
.A1(n_2262),
.A2(n_127),
.B(n_128),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2284),
.B(n_128),
.Y(n_2336)
);

NAND4xp75_ASAP7_75t_L g2337 ( 
.A(n_2289),
.B(n_134),
.C(n_131),
.D(n_133),
.Y(n_2337)
);

NAND3xp33_ASAP7_75t_L g2338 ( 
.A(n_2243),
.B(n_135),
.C(n_137),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2225),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2274),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2255),
.B(n_137),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2244),
.B(n_138),
.Y(n_2342)
);

NOR3xp33_ASAP7_75t_L g2343 ( 
.A(n_2251),
.B(n_138),
.C(n_139),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2261),
.B(n_2271),
.C(n_2246),
.Y(n_2344)
);

NOR4xp75_ASAP7_75t_L g2345 ( 
.A(n_2295),
.B(n_141),
.C(n_139),
.D(n_140),
.Y(n_2345)
);

AND4x2_ASAP7_75t_L g2346 ( 
.A(n_2277),
.B(n_142),
.C(n_140),
.D(n_141),
.Y(n_2346)
);

CKINVDCx12_ASAP7_75t_R g2347 ( 
.A(n_2257),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2237),
.B(n_2248),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2245),
.Y(n_2349)
);

NAND4xp25_ASAP7_75t_L g2350 ( 
.A(n_2231),
.B(n_144),
.C(n_142),
.D(n_143),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_SL g2351 ( 
.A(n_2249),
.B(n_144),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2263),
.A2(n_1658),
.B1(n_1472),
.B2(n_1593),
.Y(n_2352)
);

NOR3xp33_ASAP7_75t_L g2353 ( 
.A(n_2252),
.B(n_1374),
.C(n_1368),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2291),
.A2(n_1381),
.B(n_1326),
.Y(n_2354)
);

NOR3xp33_ASAP7_75t_SL g2355 ( 
.A(n_2276),
.B(n_145),
.C(n_146),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2224),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2311),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_SL g2358 ( 
.A(n_2319),
.B(n_2241),
.C(n_2235),
.Y(n_2358)
);

NOR3xp33_ASAP7_75t_L g2359 ( 
.A(n_2298),
.B(n_2293),
.C(n_2265),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2298),
.B(n_2258),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2328),
.Y(n_2361)
);

AOI22x1_ASAP7_75t_L g2362 ( 
.A1(n_2316),
.A2(n_2256),
.B1(n_2226),
.B2(n_2232),
.Y(n_2362)
);

XNOR2xp5_ASAP7_75t_L g2363 ( 
.A(n_2331),
.B(n_2236),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2299),
.B(n_2240),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2304),
.B(n_2306),
.C(n_2344),
.Y(n_2365)
);

INVx4_ASAP7_75t_L g2366 ( 
.A(n_2323),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2317),
.B(n_2296),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2318),
.Y(n_2368)
);

AO22x2_ASAP7_75t_L g2369 ( 
.A1(n_2320),
.A2(n_2228),
.B1(n_2242),
.B2(n_2268),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2332),
.B(n_147),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2318),
.Y(n_2371)
);

AO22x2_ASAP7_75t_L g2372 ( 
.A1(n_2300),
.A2(n_1546),
.B1(n_1501),
.B2(n_1500),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2336),
.Y(n_2373)
);

A2O1A1Ixp33_ASAP7_75t_L g2374 ( 
.A1(n_2312),
.A2(n_1374),
.B(n_1380),
.C(n_1368),
.Y(n_2374)
);

AOI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2348),
.A2(n_1381),
.B(n_1326),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2335),
.B(n_151),
.Y(n_2376)
);

OA22x2_ASAP7_75t_L g2377 ( 
.A1(n_2334),
.A2(n_1501),
.B1(n_1522),
.B2(n_1518),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2350),
.B(n_154),
.Y(n_2378)
);

NAND4xp75_ASAP7_75t_L g2379 ( 
.A(n_2301),
.B(n_1381),
.C(n_1256),
.D(n_1518),
.Y(n_2379)
);

NOR3xp33_ASAP7_75t_L g2380 ( 
.A(n_2340),
.B(n_1380),
.C(n_1278),
.Y(n_2380)
);

AOI221xp5_ASAP7_75t_L g2381 ( 
.A1(n_2341),
.A2(n_1581),
.B1(n_1593),
.B2(n_1375),
.C(n_1360),
.Y(n_2381)
);

AO22x1_ASAP7_75t_L g2382 ( 
.A1(n_2308),
.A2(n_1732),
.B1(n_1658),
.B2(n_1522),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2323),
.A2(n_1581),
.B1(n_1732),
.B2(n_1527),
.Y(n_2383)
);

AOI221xp5_ASAP7_75t_SL g2384 ( 
.A1(n_2313),
.A2(n_1358),
.B1(n_1375),
.B2(n_1360),
.C(n_1598),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_2329),
.B(n_1911),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2325),
.B(n_1358),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2351),
.B(n_157),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2342),
.B(n_159),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2346),
.Y(n_2389)
);

NAND4xp25_ASAP7_75t_L g2390 ( 
.A(n_2338),
.B(n_1302),
.C(n_1309),
.D(n_1296),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2347),
.Y(n_2391)
);

NAND4xp25_ASAP7_75t_L g2392 ( 
.A(n_2322),
.B(n_1302),
.C(n_1309),
.D(n_1296),
.Y(n_2392)
);

AO221x1_ASAP7_75t_L g2393 ( 
.A1(n_2333),
.A2(n_1588),
.B1(n_1574),
.B2(n_1582),
.C(n_1601),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2330),
.B(n_161),
.Y(n_2394)
);

NAND3xp33_ASAP7_75t_L g2395 ( 
.A(n_2343),
.B(n_1360),
.C(n_1358),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2345),
.Y(n_2396)
);

NAND4xp75_ASAP7_75t_L g2397 ( 
.A(n_2314),
.B(n_2321),
.C(n_2303),
.D(n_2355),
.Y(n_2397)
);

NAND4xp25_ASAP7_75t_L g2398 ( 
.A(n_2307),
.B(n_1321),
.C(n_1347),
.D(n_1317),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2349),
.Y(n_2399)
);

AOI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2352),
.A2(n_1375),
.B1(n_1360),
.B2(n_1347),
.C(n_1317),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2302),
.A2(n_1375),
.B1(n_1732),
.B2(n_1284),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2336),
.Y(n_2402)
);

O2A1O1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_2356),
.A2(n_1284),
.B(n_1276),
.C(n_1281),
.Y(n_2403)
);

NAND5xp2_ASAP7_75t_L g2404 ( 
.A(n_2305),
.B(n_163),
.C(n_166),
.D(n_171),
.E(n_172),
.Y(n_2404)
);

NOR2x1p5_ASAP7_75t_L g2405 ( 
.A(n_2337),
.B(n_1276),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2315),
.B(n_173),
.Y(n_2406)
);

NAND5xp2_ASAP7_75t_L g2407 ( 
.A(n_2309),
.B(n_178),
.C(n_179),
.D(n_181),
.E(n_182),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2366),
.Y(n_2408)
);

NOR2x1_ASAP7_75t_L g2409 ( 
.A(n_2357),
.B(n_2339),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2378),
.Y(n_2410)
);

AOI22xp5_ASAP7_75t_L g2411 ( 
.A1(n_2391),
.A2(n_2353),
.B1(n_2324),
.B2(n_2326),
.Y(n_2411)
);

O2A1O1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2389),
.A2(n_2327),
.B(n_2310),
.C(n_2354),
.Y(n_2412)
);

OAI211xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2399),
.A2(n_1281),
.B(n_1278),
.C(n_1321),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2360),
.A2(n_1588),
.B1(n_1620),
.B2(n_1601),
.Y(n_2414)
);

NAND5xp2_ASAP7_75t_L g2415 ( 
.A(n_2365),
.B(n_183),
.C(n_184),
.D(n_189),
.E(n_192),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2370),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2361),
.A2(n_1620),
.B1(n_1582),
.B2(n_1524),
.Y(n_2417)
);

AND3x2_ASAP7_75t_L g2418 ( 
.A(n_2368),
.B(n_1533),
.C(n_1527),
.Y(n_2418)
);

AOI211xp5_ASAP7_75t_L g2419 ( 
.A1(n_2396),
.A2(n_2394),
.B(n_2402),
.C(n_2376),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_SL g2420 ( 
.A1(n_2371),
.A2(n_1256),
.B1(n_1545),
.B2(n_1536),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2388),
.Y(n_2421)
);

AOI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2373),
.A2(n_1533),
.B1(n_1536),
.B2(n_1550),
.Y(n_2422)
);

INVxp33_ASAP7_75t_SL g2423 ( 
.A(n_2363),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2387),
.A2(n_2397),
.B1(n_2364),
.B2(n_2359),
.Y(n_2424)
);

OAI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2401),
.A2(n_1256),
.B1(n_1606),
.B2(n_1603),
.C(n_1596),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_SL g2426 ( 
.A1(n_2405),
.A2(n_198),
.B(n_205),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2377),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2382),
.B(n_208),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2385),
.B(n_210),
.Y(n_2429)
);

AND2x2_ASAP7_75t_SL g2430 ( 
.A(n_2364),
.B(n_1545),
.Y(n_2430)
);

OAI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2367),
.A2(n_1550),
.B1(n_1590),
.B2(n_1585),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2384),
.B(n_212),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2381),
.B(n_214),
.Y(n_2433)
);

AND2x4_ASAP7_75t_L g2434 ( 
.A(n_2358),
.B(n_215),
.Y(n_2434)
);

OA22x2_ASAP7_75t_L g2435 ( 
.A1(n_2406),
.A2(n_1591),
.B1(n_1592),
.B2(n_1594),
.Y(n_2435)
);

HB1xp67_ASAP7_75t_L g2436 ( 
.A(n_2379),
.Y(n_2436)
);

XNOR2x1_ASAP7_75t_L g2437 ( 
.A(n_2369),
.B(n_216),
.Y(n_2437)
);

OAI211xp5_ASAP7_75t_L g2438 ( 
.A1(n_2362),
.A2(n_218),
.B(n_220),
.C(n_222),
.Y(n_2438)
);

XOR2xp5_ASAP7_75t_L g2439 ( 
.A(n_2369),
.B(n_2392),
.Y(n_2439)
);

AO22x2_ASAP7_75t_L g2440 ( 
.A1(n_2386),
.A2(n_227),
.B1(n_234),
.B2(n_236),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2374),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2393),
.B(n_239),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2390),
.Y(n_2443)
);

OAI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2375),
.A2(n_1498),
.B(n_1497),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2395),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2380),
.A2(n_1649),
.B1(n_1560),
.B2(n_1557),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2372),
.Y(n_2447)
);

INVx4_ASAP7_75t_L g2448 ( 
.A(n_2372),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2383),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2398),
.B(n_240),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2403),
.B(n_241),
.Y(n_2451)
);

CKINVDCx20_ASAP7_75t_R g2452 ( 
.A(n_2404),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2400),
.B(n_243),
.Y(n_2453)
);

NOR4xp25_ASAP7_75t_L g2454 ( 
.A(n_2407),
.B(n_1549),
.C(n_1542),
.D(n_1523),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_L g2455 ( 
.A1(n_2366),
.A2(n_1563),
.B1(n_1560),
.B2(n_1552),
.C(n_1549),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2408),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2429),
.B(n_244),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2434),
.B(n_245),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2454),
.B(n_253),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_2448),
.Y(n_2460)
);

NOR3xp33_ASAP7_75t_L g2461 ( 
.A(n_2409),
.B(n_254),
.C(n_257),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2437),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2442),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2423),
.A2(n_1577),
.B1(n_1555),
.B2(n_1661),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_2416),
.A2(n_1297),
.B1(n_1308),
.B2(n_1250),
.Y(n_2465)
);

OAI211xp5_ASAP7_75t_SL g2466 ( 
.A1(n_2419),
.A2(n_258),
.B(n_266),
.C(n_267),
.Y(n_2466)
);

XNOR2x1_ASAP7_75t_L g2467 ( 
.A(n_2424),
.B(n_2410),
.Y(n_2467)
);

INVxp67_ASAP7_75t_L g2468 ( 
.A(n_2432),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2452),
.Y(n_2469)
);

NAND4xp25_ASAP7_75t_L g2470 ( 
.A(n_2426),
.B(n_2415),
.C(n_2428),
.D(n_2411),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2421),
.B(n_268),
.Y(n_2471)
);

NAND2x1_ASAP7_75t_L g2472 ( 
.A(n_2440),
.B(n_1250),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2443),
.A2(n_1297),
.B1(n_1308),
.B2(n_1250),
.Y(n_2473)
);

XNOR2xp5_ASAP7_75t_L g2474 ( 
.A(n_2439),
.B(n_270),
.Y(n_2474)
);

OAI221xp5_ASAP7_75t_L g2475 ( 
.A1(n_2438),
.A2(n_1542),
.B1(n_1523),
.B2(n_1511),
.C(n_278),
.Y(n_2475)
);

INVx1_ASAP7_75t_SL g2476 ( 
.A(n_2450),
.Y(n_2476)
);

NOR4xp25_ASAP7_75t_L g2477 ( 
.A(n_2412),
.B(n_271),
.C(n_274),
.D(n_277),
.Y(n_2477)
);

NOR3x1_ASAP7_75t_L g2478 ( 
.A(n_2433),
.B(n_282),
.C(n_286),
.Y(n_2478)
);

NAND4xp75_ASAP7_75t_L g2479 ( 
.A(n_2445),
.B(n_289),
.C(n_290),
.D(n_292),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2441),
.B(n_293),
.C(n_294),
.Y(n_2480)
);

NOR2x2_ASAP7_75t_L g2481 ( 
.A(n_2427),
.B(n_295),
.Y(n_2481)
);

AOI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_2436),
.A2(n_1336),
.B(n_1265),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2449),
.B(n_296),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2453),
.A2(n_1608),
.B1(n_1589),
.B2(n_1642),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2430),
.B(n_304),
.Y(n_2485)
);

INVx1_ASAP7_75t_SL g2486 ( 
.A(n_2451),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2414),
.B(n_305),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2456),
.A2(n_2440),
.B1(n_2435),
.B2(n_2417),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2457),
.Y(n_2489)
);

XNOR2xp5_ASAP7_75t_L g2490 ( 
.A(n_2467),
.B(n_2418),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2458),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2472),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2481),
.Y(n_2493)
);

OAI22xp5_ASAP7_75t_SL g2494 ( 
.A1(n_2469),
.A2(n_2447),
.B1(n_2455),
.B2(n_2431),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2471),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2459),
.Y(n_2496)
);

OAI22x1_ASAP7_75t_L g2497 ( 
.A1(n_2474),
.A2(n_2422),
.B1(n_2446),
.B2(n_2413),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2485),
.Y(n_2498)
);

XNOR2x1_ASAP7_75t_L g2499 ( 
.A(n_2462),
.B(n_2444),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2478),
.Y(n_2500)
);

OAI22x1_ASAP7_75t_L g2501 ( 
.A1(n_2460),
.A2(n_2425),
.B1(n_2420),
.B2(n_313),
.Y(n_2501)
);

XNOR2xp5_ASAP7_75t_L g2502 ( 
.A(n_2470),
.B(n_306),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2460),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2483),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2479),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2487),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2463),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2468),
.Y(n_2508)
);

OAI222xp33_ASAP7_75t_L g2509 ( 
.A1(n_2503),
.A2(n_2502),
.B1(n_2507),
.B2(n_2475),
.C1(n_2508),
.C2(n_2505),
.Y(n_2509)
);

AO22x2_ASAP7_75t_L g2510 ( 
.A1(n_2495),
.A2(n_2486),
.B1(n_2476),
.B2(n_2461),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_SL g2511 ( 
.A1(n_2498),
.A2(n_2482),
.B1(n_2484),
.B2(n_2466),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2493),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_L g2513 ( 
.A(n_2494),
.B(n_2480),
.C(n_2464),
.Y(n_2513)
);

XNOR2xp5_ASAP7_75t_L g2514 ( 
.A(n_2490),
.B(n_2477),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2492),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2500),
.Y(n_2516)
);

OAI221xp5_ASAP7_75t_L g2517 ( 
.A1(n_2488),
.A2(n_2473),
.B1(n_2465),
.B2(n_316),
.C(n_318),
.Y(n_2517)
);

OAI222xp33_ASAP7_75t_L g2518 ( 
.A1(n_2504),
.A2(n_2496),
.B1(n_2491),
.B2(n_2489),
.C1(n_2506),
.C2(n_2497),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2499),
.Y(n_2519)
);

OAI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2501),
.A2(n_1497),
.B1(n_1498),
.B2(n_1621),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2503),
.Y(n_2521)
);

OAI221xp5_ASAP7_75t_SL g2522 ( 
.A1(n_2503),
.A2(n_308),
.B1(n_315),
.B2(n_321),
.C(n_323),
.Y(n_2522)
);

OAI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2503),
.A2(n_1638),
.B1(n_1629),
.B2(n_1618),
.Y(n_2523)
);

OAI221xp5_ASAP7_75t_L g2524 ( 
.A1(n_2503),
.A2(n_324),
.B1(n_325),
.B2(n_327),
.C(n_331),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2503),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2521),
.A2(n_2525),
.B1(n_2515),
.B2(n_2519),
.Y(n_2526)
);

OAI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_2512),
.A2(n_1345),
.B1(n_1286),
.B2(n_1297),
.Y(n_2527)
);

INVxp67_ASAP7_75t_L g2528 ( 
.A(n_2515),
.Y(n_2528)
);

HB1xp67_ASAP7_75t_L g2529 ( 
.A(n_2514),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2510),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2516),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2511),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2513),
.A2(n_1336),
.B1(n_1286),
.B2(n_1297),
.Y(n_2533)
);

AO22x2_ASAP7_75t_L g2534 ( 
.A1(n_2520),
.A2(n_1475),
.B1(n_1464),
.B2(n_1463),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2517),
.Y(n_2535)
);

XNOR2xp5_ASAP7_75t_L g2536 ( 
.A(n_2518),
.B(n_2524),
.Y(n_2536)
);

AO22x2_ASAP7_75t_L g2537 ( 
.A1(n_2509),
.A2(n_1475),
.B1(n_1464),
.B2(n_1463),
.Y(n_2537)
);

CKINVDCx20_ASAP7_75t_R g2538 ( 
.A(n_2523),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2537),
.Y(n_2539)
);

XNOR2xp5_ASAP7_75t_L g2540 ( 
.A(n_2529),
.B(n_2522),
.Y(n_2540)
);

INVx4_ASAP7_75t_L g2541 ( 
.A(n_2530),
.Y(n_2541)
);

AND2x2_ASAP7_75t_SL g2542 ( 
.A(n_2526),
.B(n_1265),
.Y(n_2542)
);

XNOR2xp5_ASAP7_75t_L g2543 ( 
.A(n_2536),
.B(n_338),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2531),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2528),
.B(n_342),
.Y(n_2545)
);

NAND4xp75_ASAP7_75t_L g2546 ( 
.A(n_2535),
.B(n_1461),
.C(n_1459),
.D(n_350),
.Y(n_2546)
);

AOI21xp33_ASAP7_75t_SL g2547 ( 
.A1(n_2544),
.A2(n_2527),
.B(n_2533),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2540),
.A2(n_2538),
.B(n_2534),
.Y(n_2548)
);

XNOR2xp5_ASAP7_75t_L g2549 ( 
.A(n_2543),
.B(n_2532),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2541),
.A2(n_1124),
.B(n_1345),
.Y(n_2550)
);

AO21x1_ASAP7_75t_L g2551 ( 
.A1(n_2545),
.A2(n_1461),
.B(n_347),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2542),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2549),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2551),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2552),
.Y(n_2555)
);

XNOR2xp5_ASAP7_75t_L g2556 ( 
.A(n_2548),
.B(n_2539),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2547),
.Y(n_2557)
);

OAI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2555),
.A2(n_2550),
.B(n_2546),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2557),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2554),
.B(n_344),
.Y(n_2560)
);

AO22x2_ASAP7_75t_L g2561 ( 
.A1(n_2559),
.A2(n_2553),
.B1(n_2556),
.B2(n_361),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2558),
.B(n_356),
.Y(n_2562)
);

AOI221xp5_ASAP7_75t_L g2563 ( 
.A1(n_2561),
.A2(n_2560),
.B1(n_1345),
.B2(n_1336),
.C(n_1329),
.Y(n_2563)
);

OR2x6_ASAP7_75t_L g2564 ( 
.A(n_2562),
.B(n_1345),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2562),
.B(n_358),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2564),
.A2(n_2563),
.B(n_2565),
.Y(n_2566)
);

AOI211xp5_ASAP7_75t_L g2567 ( 
.A1(n_2566),
.A2(n_1329),
.B(n_1286),
.C(n_1308),
.Y(n_2567)
);


endmodule