module fake_jpeg_32184_n_418 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

HAxp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_0),
.CON(n_49),
.SN(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_49),
.A2(n_65),
.B(n_33),
.C(n_1),
.Y(n_119)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_0),
.B(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_84),
.Y(n_90)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_92),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_40),
.B1(n_26),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_89),
.A2(n_93),
.B1(n_97),
.B2(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_45),
.B(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_40),
.B1(n_29),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_44),
.A2(n_66),
.B1(n_78),
.B2(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_30),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_29),
.B1(n_39),
.B2(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_75),
.B1(n_29),
.B2(n_74),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_26),
.B1(n_39),
.B2(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_41),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_121),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_33),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_74),
.B(n_34),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_19),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_145),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_127),
.Y(n_141)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_153),
.B1(n_161),
.B2(n_163),
.Y(n_182)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_156),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_76),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_155),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_29),
.B1(n_20),
.B2(n_30),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_60),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_115),
.C(n_94),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_29),
.B1(n_130),
.B2(n_114),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_164)
);

OR2x4_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_21),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_93),
.A2(n_55),
.B1(n_79),
.B2(n_29),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_168),
.Y(n_177)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_145),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_105),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_140),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_188),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_201),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_138),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_167),
.B1(n_161),
.B2(n_137),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_212),
.B1(n_178),
.B2(n_177),
.Y(n_216)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_211),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_209),
.C(n_210),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_184),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_140),
.B1(n_164),
.B2(n_101),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_178),
.B1(n_150),
.B2(n_162),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_152),
.B(n_141),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_178),
.B(n_184),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_171),
.B(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_154),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_166),
.B1(n_89),
.B2(n_162),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_220),
.B(n_212),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_177),
.B1(n_182),
.B2(n_181),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_222),
.B1(n_227),
.B2(n_231),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_181),
.B1(n_187),
.B2(n_178),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_201),
.B1(n_209),
.B2(n_199),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_232),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_208),
.B(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_176),
.B1(n_175),
.B2(n_183),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_150),
.C(n_147),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.C(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_172),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_200),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_176),
.B1(n_175),
.B2(n_183),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_172),
.C(n_174),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_235),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_232),
.C(n_213),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_230),
.B1(n_231),
.B2(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_221),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_197),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_244),
.B(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_216),
.A2(n_203),
.B1(n_196),
.B2(n_211),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_243),
.B(n_228),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_212),
.B1(n_194),
.B2(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_247),
.B1(n_250),
.B2(n_219),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_252),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_222),
.A2(n_175),
.B1(n_172),
.B2(n_204),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_202),
.B(n_189),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_139),
.B1(n_204),
.B2(n_190),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_224),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_220),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_217),
.C(n_233),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_267),
.C(n_238),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_240),
.B1(n_246),
.B2(n_252),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_218),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_256),
.B(n_257),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_272),
.C(n_251),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_269),
.B1(n_271),
.B2(n_273),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_240),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_233),
.B(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_231),
.B1(n_227),
.B2(n_222),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_225),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_215),
.B1(n_219),
.B2(n_223),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_228),
.C(n_191),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_224),
.B1(n_180),
.B2(n_136),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_243),
.B(n_247),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_248),
.B(n_242),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_280),
.B(n_266),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_237),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_276),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_292),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_240),
.B(n_244),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_259),
.C(n_257),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_295),
.C(n_155),
.Y(n_304)
);

NAND2x1_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_296),
.B1(n_141),
.B2(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_185),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_269),
.B1(n_260),
.B2(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_180),
.C(n_185),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_265),
.A2(n_88),
.B1(n_168),
.B2(n_165),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_266),
.B1(n_273),
.B2(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_297),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_318),
.C(n_320),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_319),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_264),
.B1(n_88),
.B2(n_111),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_111),
.B1(n_94),
.B2(n_143),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_308),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_160),
.B1(n_173),
.B2(n_135),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_156),
.B1(n_169),
.B2(n_146),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_99),
.B1(n_117),
.B2(n_131),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_307),
.A2(n_313),
.B1(n_296),
.B2(n_290),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_149),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_159),
.B1(n_148),
.B2(n_157),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_315),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_144),
.C(n_85),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_170),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_85),
.C(n_103),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_294),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_329),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_125),
.B1(n_2),
.B2(n_3),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_310),
.A2(n_285),
.B1(n_294),
.B2(n_275),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_327),
.A2(n_339),
.B1(n_22),
.B2(n_36),
.Y(n_357)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_303),
.A2(n_289),
.B1(n_280),
.B2(n_287),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_295),
.C(n_287),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_332),
.C(n_334),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_132),
.B1(n_96),
.B2(n_106),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_108),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_86),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_118),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_320),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_102),
.B1(n_112),
.B2(n_86),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_98),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_125),
.C(n_112),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_309),
.B(n_297),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_347),
.B(n_2),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_337),
.B(n_317),
.CI(n_309),
.CON(n_344),
.SN(n_344)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_349),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_355),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_335),
.A2(n_318),
.B(n_307),
.Y(n_347)
);

INVx11_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_337),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_353),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_330),
.A2(n_301),
.B1(n_98),
.B2(n_32),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_357),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_358),
.A2(n_321),
.B1(n_36),
.B2(n_338),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_350),
.C(n_322),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_363),
.C(n_369),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_364),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_322),
.C(n_321),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_334),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_374),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_332),
.Y(n_368)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_2),
.C(n_5),
.Y(n_369)
);

INVx11_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_345),
.Y(n_378)
);

INVx11_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_377),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_344),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_378),
.B(n_358),
.Y(n_390)
);

NOR3xp33_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_345),
.C(n_351),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_382),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_365),
.B(n_360),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_359),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_356),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_355),
.B(n_351),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_386),
.A2(n_369),
.B(n_348),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_388),
.B(n_390),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_367),
.B(n_362),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_389),
.A2(n_381),
.B(n_6),
.Y(n_400)
);

OAI21x1_ASAP7_75t_SL g392 ( 
.A1(n_375),
.A2(n_367),
.B(n_372),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_392),
.A2(n_383),
.B(n_379),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_352),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_SL g405 ( 
.A(n_398),
.B(n_401),
.C(n_399),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_400),
.B(n_402),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_394),
.A2(n_5),
.B(n_6),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_5),
.C(n_6),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_390),
.B1(n_8),
.B2(n_9),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_9),
.C(n_10),
.Y(n_409)
);

OAI311xp33_ASAP7_75t_L g410 ( 
.A1(n_405),
.A2(n_397),
.A3(n_12),
.B1(n_13),
.C1(n_14),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_7),
.B(n_8),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_408),
.B(n_11),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_409),
.A2(n_11),
.B(n_12),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_406),
.B(n_13),
.C(n_14),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_412),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_413),
.B(n_11),
.Y(n_415)
);

A2O1A1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_415),
.A2(n_414),
.B(n_15),
.C(n_16),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_11),
.C(n_16),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_417),
.A2(n_16),
.B(n_404),
.Y(n_418)
);


endmodule