module real_jpeg_21558_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_0),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_0),
.A2(n_29),
.B1(n_33),
.B2(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_29),
.B1(n_33),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_49),
.B1(n_52),
.B2(n_64),
.Y(n_139)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_24),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_3),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_25),
.B(n_106),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_33),
.B(n_58),
.C(n_66),
.D(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_28),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_47),
.B(n_140),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_24),
.B(n_38),
.C(n_71),
.D(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_46),
.B1(n_50),
.B2(n_53),
.Y(n_45)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_50),
.B(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_6),
.A2(n_46),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_37),
.B1(n_49),
.B2(n_52),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_37),
.B1(n_92),
.B2(n_97),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_26),
.B1(n_49),
.B2(n_52),
.Y(n_146)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_77),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_77),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_56),
.C(n_69),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_20),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_55),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_41),
.C(n_45),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_23),
.A2(n_27),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_28),
.B(n_30),
.C(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_27),
.B(n_36),
.Y(n_169)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_29),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_33),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_42),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_44),
.B(n_92),
.C(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_92),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_44),
.A2(n_92),
.B(n_96),
.C(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_47),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

NAND2x1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_49),
.A2(n_60),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_52),
.B(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_52),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_56),
.B(n_69),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_65),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_83),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_82),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_67),
.B(n_96),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_70),
.B(n_74),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_76),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_101),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_95),
.B(n_98),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_146),
.B(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_175),
.B(n_179),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_162),
.B(n_174),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_142),
.B(n_161),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_136),
.C(n_138),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_139),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_150),
.B(n_160),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_148),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_155),
.B(n_159),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_R g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_164),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_173),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_171),
.C(n_173),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_177),
.Y(n_179)
);


endmodule