module fake_ariane_2721_n_1095 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1095);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1095;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_940;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_989;
wire n_242;
wire n_645;
wire n_858;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_894;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_192;
wire n_887;
wire n_729;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_991;
wire n_750;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_SL g189 ( 
.A(n_109),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_3),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_30),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_26),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_64),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_58),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_77),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_76),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_137),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_70),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_14),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_120),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_41),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_95),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_56),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_117),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_127),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_29),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_25),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_108),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_28),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_104),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_31),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_143),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_14),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_110),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_51),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_101),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_179),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_144),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_83),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_191),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_216),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_206),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_195),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_228),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_246),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_196),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_198),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_208),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_200),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_202),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_204),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_218),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_218),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_269),
.A2(n_222),
.B1(n_250),
.B2(n_226),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_201),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_189),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

OAI22x1_ASAP7_75t_SL g317 ( 
.A1(n_269),
.A2(n_207),
.B1(n_240),
.B2(n_226),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_266),
.A2(n_268),
.B1(n_287),
.B2(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_286),
.A2(n_222),
.B1(n_250),
.B2(n_212),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_209),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_214),
.B(n_211),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_239),
.Y(n_335)
);

BUFx8_ASAP7_75t_SL g336 ( 
.A(n_286),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_275),
.A2(n_225),
.B(n_239),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_217),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_220),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_239),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_281),
.A2(n_224),
.B(n_223),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_279),
.A2(n_242),
.B1(n_260),
.B2(n_259),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_282),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_280),
.A2(n_238),
.B1(n_258),
.B2(n_257),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_248),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_288),
.Y(n_358)
);

CKINVDCx6p67_ASAP7_75t_R g359 ( 
.A(n_273),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_267),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_302),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_312),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_R g374 ( 
.A(n_359),
.B(n_304),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_336),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_359),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_323),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_R g380 ( 
.A(n_350),
.B(n_306),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_R g381 ( 
.A(n_341),
.B(n_306),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_324),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_326),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_352),
.B(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_341),
.B(n_308),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_341),
.B(n_229),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_353),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_314),
.B(n_248),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_337),
.A2(n_234),
.B(n_230),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_330),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g412 ( 
.A(n_351),
.B(n_235),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_313),
.A2(n_245),
.B1(n_256),
.B2(n_249),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_338),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_317),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_343),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_340),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_318),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_344),
.B(n_236),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_357),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_357),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_358),
.Y(n_424)
);

BUFx10_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_358),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_339),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_339),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_339),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_339),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_347),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_361),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_371),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_374),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_356),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_354),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_351),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_351),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_332),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_378),
.B(n_419),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_416),
.B(n_329),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_379),
.B(n_332),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_381),
.B(n_400),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_372),
.B(n_329),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_380),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_426),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_381),
.B(n_362),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_425),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_421),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_375),
.B(n_321),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_373),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_386),
.B(n_334),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_400),
.B(n_362),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_375),
.B(n_364),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_438),
.B(n_345),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_404),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_423),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_383),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_406),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_413),
.A2(n_332),
.B1(n_346),
.B2(n_345),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_439),
.A2(n_346),
.B1(n_345),
.B2(n_362),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_366),
.B(n_345),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_406),
.B(n_335),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_390),
.B(n_346),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_380),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_401),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_410),
.B(n_346),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_377),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_327),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_436),
.B(n_327),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_367),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_453),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_414),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_460),
.B(n_420),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_488),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_376),
.C(n_415),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_469),
.A2(n_408),
.B1(n_412),
.B2(n_407),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_474),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_480),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_441),
.Y(n_539)
);

OR2x2_ASAP7_75t_SL g540 ( 
.A(n_513),
.B(n_407),
.Y(n_540)
);

OR2x2_ASAP7_75t_SL g541 ( 
.A(n_464),
.B(n_524),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_433),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_495),
.B(n_452),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_469),
.A2(n_431),
.B1(n_362),
.B2(n_327),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_453),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_445),
.A2(n_446),
.B1(n_485),
.B2(n_492),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_477),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_476),
.B(n_362),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_524),
.A2(n_412),
.B1(n_1),
.B2(n_2),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_488),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_444),
.B(n_327),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_476),
.B(n_327),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

OR2x6_ASAP7_75t_SL g560 ( 
.A(n_449),
.B(n_237),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_478),
.B(n_337),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_497),
.B(n_316),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_466),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_457),
.A2(n_319),
.B1(n_316),
.B2(n_225),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_501),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_490),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_466),
.B(n_470),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_488),
.B(n_473),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_490),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

AND2x6_ASAP7_75t_SL g572 ( 
.A(n_473),
.B(n_0),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_465),
.Y(n_573)
);

NAND3x1_ASAP7_75t_L g574 ( 
.A(n_465),
.B(n_319),
.C(n_316),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_495),
.B(n_319),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_456),
.B(n_485),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_525),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_492),
.B(n_4),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_482),
.B(n_320),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_455),
.A2(n_225),
.B1(n_320),
.B2(n_322),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_455),
.B(n_5),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_496),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_5),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_519),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_SL g588 ( 
.A(n_449),
.B(n_6),
.C(n_7),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_482),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_6),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_525),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_543),
.B(n_472),
.Y(n_593)
);

AOI21x1_ASAP7_75t_L g594 ( 
.A1(n_577),
.A2(n_459),
.B(n_521),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_558),
.B(n_481),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_561),
.A2(n_577),
.B(n_542),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_531),
.A2(n_506),
.B(n_515),
.C(n_516),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_481),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_561),
.A2(n_506),
.B(n_489),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_563),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_556),
.A2(n_479),
.B(n_447),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_546),
.A2(n_505),
.B1(n_484),
.B2(n_481),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_527),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_556),
.A2(n_521),
.B(n_512),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_546),
.A2(n_515),
.B(n_516),
.C(n_522),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_551),
.A2(n_522),
.B(n_511),
.C(n_512),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_579),
.B(n_484),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_447),
.B(n_443),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_536),
.B(n_475),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_537),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_575),
.A2(n_493),
.B(n_486),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_558),
.B(n_467),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_573),
.B(n_464),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_530),
.B(n_484),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_559),
.A2(n_511),
.B(n_509),
.C(n_508),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_569),
.B(n_505),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_567),
.A2(n_447),
.B(n_443),
.Y(n_619)
);

CKINVDCx6p67_ASAP7_75t_R g620 ( 
.A(n_529),
.Y(n_620)
);

AOI33xp33_ASAP7_75t_L g621 ( 
.A1(n_528),
.A2(n_548),
.A3(n_550),
.B1(n_549),
.B2(n_535),
.B3(n_566),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_505),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_450),
.B(n_443),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_571),
.A2(n_454),
.B(n_450),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_563),
.B(n_500),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_591),
.B(n_464),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_582),
.A2(n_508),
.B1(n_487),
.B2(n_475),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_584),
.A2(n_454),
.B(n_450),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_585),
.B(n_511),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_530),
.B(n_520),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_565),
.B(n_510),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_564),
.A2(n_517),
.B(n_586),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_590),
.A2(n_454),
.B(n_468),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_557),
.A2(n_468),
.B(n_517),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_539),
.B(n_510),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_588),
.B(n_523),
.C(n_519),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_562),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_555),
.B(n_510),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_564),
.A2(n_493),
.B(n_486),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_576),
.B(n_520),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_578),
.A2(n_592),
.B1(n_508),
.B2(n_487),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

BUFx12f_ASAP7_75t_L g643 ( 
.A(n_587),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_576),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_547),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_552),
.A2(n_468),
.B(n_463),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_576),
.B(n_523),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_581),
.A2(n_463),
.B(n_487),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_589),
.B(n_510),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_589),
.B(n_510),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_599),
.B(n_589),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_593),
.B(n_534),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_603),
.B(n_608),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_560),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_629),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_614),
.B(n_553),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_597),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_611),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_637),
.B(n_553),
.Y(n_659)
);

NOR2x1_ASAP7_75t_R g660 ( 
.A(n_643),
.B(n_538),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_606),
.A2(n_545),
.B(n_533),
.C(n_568),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_647),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_630),
.A2(n_534),
.B1(n_544),
.B2(n_592),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_620),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_600),
.A2(n_574),
.B(n_581),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_604),
.A2(n_578),
.B1(n_541),
.B2(n_529),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_622),
.A2(n_503),
.B1(n_562),
.B2(n_540),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_641),
.A2(n_494),
.B1(n_514),
.B2(n_507),
.Y(n_669)
);

INVx3_ASAP7_75t_SL g670 ( 
.A(n_601),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_605),
.A2(n_471),
.B(n_467),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_607),
.A2(n_494),
.B1(n_507),
.B2(n_514),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_618),
.B(n_572),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_621),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_644),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_642),
.B(n_580),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_617),
.B(n_631),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_601),
.B(n_580),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_601),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_610),
.B(n_520),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_612),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_599),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_625),
.B(n_467),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_615),
.A2(n_483),
.B1(n_467),
.B2(n_504),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_605),
.A2(n_467),
.B(n_483),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_645),
.B(n_8),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_640),
.B(n_483),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_635),
.B(n_572),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_649),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_650),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_617),
.B(n_461),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_627),
.B(n_483),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_638),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_636),
.B(n_483),
.Y(n_695)
);

O2A1O1Ixp5_ASAP7_75t_L g696 ( 
.A1(n_632),
.A2(n_462),
.B(n_461),
.C(n_458),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_SL g697 ( 
.A(n_598),
.B(n_616),
.C(n_595),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_595),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_639),
.A2(n_462),
.B(n_458),
.C(n_448),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_613),
.B(n_448),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_648),
.B(n_322),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_594),
.A2(n_510),
.B(n_225),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_609),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_633),
.B(n_225),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_619),
.B(n_10),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_634),
.A2(n_261),
.B(n_248),
.Y(n_706)
);

AOI222xp33_ASAP7_75t_L g707 ( 
.A1(n_623),
.A2(n_261),
.B1(n_248),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_707)
);

CKINVDCx8_ASAP7_75t_R g708 ( 
.A(n_624),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_657),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_682),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_658),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_670),
.Y(n_712)
);

BUFx2_ASAP7_75t_SL g713 ( 
.A(n_675),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_679),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_684),
.B(n_628),
.Y(n_715)
);

BUFx2_ASAP7_75t_SL g716 ( 
.A(n_665),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_663),
.Y(n_717)
);

INVx6_ASAP7_75t_L g718 ( 
.A(n_679),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_674),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_673),
.B(n_10),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_690),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_659),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_654),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_691),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_694),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_656),
.B(n_646),
.Y(n_726)
);

BUFx12f_ASAP7_75t_L g727 ( 
.A(n_679),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_651),
.Y(n_728)
);

BUFx4_ASAP7_75t_SL g729 ( 
.A(n_660),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_676),
.B(n_11),
.Y(n_730)
);

BUFx4_ASAP7_75t_SL g731 ( 
.A(n_661),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_651),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_708),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_662),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_689),
.B(n_11),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_677),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_688),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_667),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_678),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_687),
.B(n_12),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_667),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_652),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_664),
.B(n_13),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_652),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_677),
.Y(n_749)
);

BUFx4_ASAP7_75t_SL g750 ( 
.A(n_680),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_683),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_701),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_705),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_655),
.Y(n_755)
);

BUFx4_ASAP7_75t_SL g756 ( 
.A(n_695),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_701),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_653),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_666),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_655),
.B(n_15),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_669),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_700),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_693),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_707),
.B(n_16),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_668),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_668),
.B(n_16),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_685),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_702),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_755),
.B(n_738),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_SL g771 ( 
.A(n_733),
.B(n_671),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_767),
.A2(n_669),
.B1(n_672),
.B2(n_685),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_738),
.B(n_681),
.Y(n_773)
);

AOI21x1_ASAP7_75t_L g774 ( 
.A1(n_760),
.A2(n_704),
.B(n_706),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_712),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_722),
.B(n_686),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_769),
.A2(n_704),
.B(n_696),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_733),
.Y(n_778)
);

AOI222xp33_ASAP7_75t_L g779 ( 
.A1(n_765),
.A2(n_672),
.B1(n_697),
.B2(n_261),
.C1(n_699),
.C2(n_21),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_722),
.B(n_17),
.Y(n_780)
);

AO21x2_ASAP7_75t_L g781 ( 
.A1(n_719),
.A2(n_725),
.B(n_743),
.Y(n_781)
);

BUFx8_ASAP7_75t_L g782 ( 
.A(n_712),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_720),
.A2(n_602),
.B(n_18),
.C(n_19),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_758),
.B(n_737),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_712),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_766),
.A2(n_225),
.B1(n_261),
.B2(n_19),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_769),
.A2(n_34),
.B(n_33),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_721),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_740),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_735),
.A2(n_36),
.B(n_35),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_740),
.B(n_20),
.Y(n_792)
);

AOI22x1_ASAP7_75t_L g793 ( 
.A1(n_713),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_SL g794 ( 
.A1(n_761),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_744),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_749),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_709),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_744),
.B(n_27),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_726),
.A2(n_128),
.B(n_185),
.Y(n_799)
);

OA21x2_ASAP7_75t_L g800 ( 
.A1(n_759),
.A2(n_28),
.B(n_29),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_754),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_762),
.B(n_37),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_714),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_714),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_754),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_746),
.B(n_38),
.Y(n_806)
);

CKINVDCx11_ASAP7_75t_R g807 ( 
.A(n_723),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_711),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_734),
.B(n_40),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_747),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_724),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_728),
.A2(n_47),
.B(n_48),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_768),
.A2(n_49),
.B(n_52),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_763),
.A2(n_54),
.B(n_55),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_728),
.A2(n_57),
.B(n_59),
.Y(n_815)
);

INVx5_ASAP7_75t_L g816 ( 
.A(n_754),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_764),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_714),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_730),
.A2(n_60),
.B(n_63),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_717),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_736),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_764),
.B(n_68),
.Y(n_822)
);

OAI21xp33_ASAP7_75t_SL g823 ( 
.A1(n_739),
.A2(n_71),
.B(n_72),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_763),
.A2(n_74),
.B(n_75),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_731),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_817),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_781),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_781),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_801),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_797),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_808),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_796),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_811),
.Y(n_834)
);

AO21x2_ASAP7_75t_L g835 ( 
.A1(n_773),
.A2(n_715),
.B(n_742),
.Y(n_835)
);

CKINVDCx11_ASAP7_75t_R g836 ( 
.A(n_807),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_803),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_770),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_804),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_770),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_826),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_773),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_776),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_776),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_774),
.A2(n_732),
.B(n_756),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_801),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_788),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_821),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_805),
.Y(n_850)
);

BUFx8_ASAP7_75t_L g851 ( 
.A(n_821),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_805),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_816),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_786),
.A2(n_751),
.B1(n_748),
.B2(n_745),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_798),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_778),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_800),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_814),
.A2(n_757),
.B(n_753),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_778),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_818),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_800),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_816),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_814),
.A2(n_757),
.B(n_753),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_784),
.B(n_739),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_816),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_779),
.A2(n_741),
.B1(n_710),
.B2(n_752),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_816),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_790),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_771),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_833),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_SL g871 ( 
.A1(n_854),
.A2(n_795),
.B(n_789),
.C(n_825),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_854),
.A2(n_789),
.B1(n_795),
.B2(n_786),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_866),
.A2(n_772),
.B1(n_793),
.B2(n_784),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_833),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_827),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_857),
.A2(n_783),
.B(n_813),
.C(n_772),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_855),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_837),
.B(n_785),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_837),
.B(n_807),
.Y(n_879)
);

INVxp67_ASAP7_75t_R g880 ( 
.A(n_864),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_838),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_856),
.B(n_821),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_838),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_857),
.A2(n_783),
.B(n_825),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_863),
.A2(n_822),
.B(n_813),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_841),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_840),
.B(n_775),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_861),
.A2(n_855),
.B1(n_846),
.B2(n_835),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_836),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_841),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_845),
.B(n_791),
.Y(n_891)
);

OR2x2_ASAP7_75t_SL g892 ( 
.A(n_846),
.B(n_780),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_869),
.A2(n_820),
.B(n_823),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_840),
.Y(n_894)
);

INVxp33_ASAP7_75t_L g895 ( 
.A(n_867),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_R g896 ( 
.A(n_846),
.B(n_806),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_860),
.B(n_716),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_860),
.B(n_802),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_851),
.B(n_782),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_891),
.B(n_845),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_881),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_891),
.B(n_845),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_877),
.B(n_835),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_894),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_880),
.B(n_845),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_870),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_889),
.B(n_782),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_878),
.B(n_859),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_879),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_897),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_882),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_892),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_883),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_874),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_887),
.B(n_864),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_886),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_890),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_875),
.B(n_835),
.Y(n_918)
);

AOI221xp5_ASAP7_75t_L g919 ( 
.A1(n_871),
.A2(n_861),
.B1(n_794),
.B2(n_820),
.C(n_843),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_895),
.B(n_835),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_895),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_885),
.B(n_869),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_909),
.Y(n_923)
);

AO31x2_ASAP7_75t_L g924 ( 
.A1(n_913),
.A2(n_876),
.A3(n_828),
.B(n_829),
.Y(n_924)
);

AO21x2_ASAP7_75t_L g925 ( 
.A1(n_922),
.A2(n_884),
.B(n_876),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_901),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_919),
.A2(n_872),
.B1(n_873),
.B2(n_893),
.Y(n_927)
);

NOR2x1_ASAP7_75t_SL g928 ( 
.A(n_903),
.B(n_898),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_920),
.A2(n_829),
.B(n_828),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_911),
.B(n_888),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_911),
.A2(n_871),
.B(n_872),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_852),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_912),
.A2(n_873),
.B1(n_844),
.B2(n_847),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_901),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_903),
.B(n_844),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_922),
.B(n_896),
.C(n_852),
.Y(n_937)
);

AOI221xp5_ASAP7_75t_SL g938 ( 
.A1(n_921),
.A2(n_810),
.B1(n_839),
.B2(n_865),
.C(n_862),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_925),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_923),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_931),
.B(n_930),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_930),
.B(n_909),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_927),
.A2(n_937),
.B1(n_912),
.B2(n_933),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_926),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_935),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_932),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_932),
.B(n_846),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_925),
.A2(n_896),
.B1(n_922),
.B2(n_917),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_932),
.B(n_908),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_934),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_907),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_940),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_944),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_950),
.B(n_927),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_942),
.B(n_945),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_946),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_949),
.B(n_910),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_946),
.B(n_910),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_954),
.B(n_943),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_953),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_955),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_915),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_954),
.B(n_939),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_952),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_952),
.B(n_939),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_956),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_959),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_962),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_961),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_965),
.B(n_943),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_963),
.A2(n_948),
.B1(n_947),
.B2(n_951),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_963),
.B(n_729),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_966),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_964),
.B(n_958),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_962),
.B(n_915),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_L g978 ( 
.A(n_976),
.B(n_899),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_967),
.B(n_938),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_970),
.Y(n_980)
);

OAI211xp5_ASAP7_75t_L g981 ( 
.A1(n_971),
.A2(n_899),
.B(n_791),
.C(n_794),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_921),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_973),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_968),
.B(n_922),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_974),
.B(n_918),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_980),
.B(n_969),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_982),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_986),
.Y(n_989)
);

AOI211xp5_ASAP7_75t_SL g990 ( 
.A1(n_983),
.A2(n_975),
.B(n_977),
.C(n_972),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_978),
.Y(n_991)
);

OAI22xp33_ASAP7_75t_L g992 ( 
.A1(n_979),
.A2(n_947),
.B1(n_975),
.B2(n_936),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_981),
.A2(n_984),
.B1(n_985),
.B2(n_947),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_980),
.B(n_928),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_986),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_989),
.B(n_904),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_995),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_L g998 ( 
.A(n_987),
.B(n_904),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_936),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_991),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_990),
.B(n_924),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_992),
.B(n_924),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

NOR2x1_ASAP7_75t_L g1004 ( 
.A(n_993),
.B(n_710),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_924),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_914),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_914),
.B1(n_916),
.B2(n_906),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_996),
.B(n_908),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_998),
.B(n_1004),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_1002),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1001),
.B(n_924),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1000),
.B(n_916),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1000),
.B(n_913),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_1010),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.Y(n_1016)
);

NAND4xp25_ASAP7_75t_L g1017 ( 
.A(n_1014),
.B(n_905),
.C(n_902),
.D(n_900),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1005),
.Y(n_1018)
);

AOI222xp33_ASAP7_75t_L g1019 ( 
.A1(n_1012),
.A2(n_929),
.B1(n_810),
.B2(n_822),
.C1(n_868),
.C2(n_710),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_1007),
.B(n_917),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_1011),
.B(n_819),
.C(n_812),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_1013),
.B(n_900),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_SL g1023 ( 
.A1(n_1016),
.A2(n_1009),
.B1(n_1008),
.B2(n_920),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_1018),
.A2(n_929),
.B(n_790),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_SL g1025 ( 
.A1(n_1015),
.A2(n_1020),
.B1(n_1022),
.B2(n_1017),
.C(n_1021),
.Y(n_1025)
);

OAI211xp5_ASAP7_75t_L g1026 ( 
.A1(n_1019),
.A2(n_905),
.B(n_787),
.C(n_821),
.Y(n_1026)
);

OAI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1015),
.A2(n_815),
.B(n_824),
.C(n_839),
.Y(n_1027)
);

OAI211xp5_ASAP7_75t_SL g1028 ( 
.A1(n_1015),
.A2(n_839),
.B(n_830),
.C(n_847),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1015),
.A2(n_900),
.B(n_902),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1025),
.A2(n_868),
.B1(n_829),
.B2(n_809),
.C(n_830),
.Y(n_1030)
);

AND4x1_ASAP7_75t_L g1031 ( 
.A(n_1029),
.B(n_750),
.C(n_809),
.D(n_865),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_1023),
.A2(n_1026),
.B1(n_1024),
.B2(n_1028),
.C(n_1027),
.Y(n_1032)
);

NAND4xp75_ASAP7_75t_L g1033 ( 
.A(n_1025),
.B(n_862),
.C(n_850),
.D(n_853),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_868),
.B1(n_850),
.B2(n_902),
.C(n_900),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1023),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_1025),
.Y(n_1036)
);

AOI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1025),
.A2(n_902),
.B1(n_848),
.B2(n_843),
.C(n_741),
.Y(n_1037)
);

AOI222xp33_ASAP7_75t_L g1038 ( 
.A1(n_1026),
.A2(n_799),
.B1(n_848),
.B2(n_843),
.C1(n_741),
.C2(n_832),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_1025),
.A2(n_831),
.B1(n_832),
.B2(n_834),
.C(n_842),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_849),
.Y(n_1040)
);

AOI322xp5_ASAP7_75t_L g1041 ( 
.A1(n_1035),
.A2(n_853),
.A3(n_831),
.B1(n_832),
.B2(n_834),
.C1(n_842),
.C2(n_736),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_1033),
.Y(n_1042)
);

AOI311xp33_ASAP7_75t_L g1043 ( 
.A1(n_1032),
.A2(n_849),
.A3(n_851),
.B(n_718),
.C(n_85),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_718),
.Y(n_1044)
);

OAI211xp5_ASAP7_75t_L g1045 ( 
.A1(n_1034),
.A2(n_736),
.B(n_745),
.C(n_851),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1030),
.A2(n_853),
.B1(n_734),
.B2(n_831),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_1037),
.A2(n_842),
.B(n_82),
.C(n_84),
.Y(n_1047)
);

AOI32xp33_ASAP7_75t_L g1048 ( 
.A1(n_1038),
.A2(n_863),
.A3(n_858),
.B1(n_834),
.B2(n_849),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_863),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_1042),
.B(n_81),
.C(n_86),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1040),
.B(n_849),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1044),
.A2(n_87),
.B(n_88),
.C(n_89),
.Y(n_1052)
);

NAND4xp75_ASAP7_75t_L g1053 ( 
.A(n_1043),
.B(n_90),
.C(n_91),
.D(n_92),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1045),
.B(n_94),
.C(n_96),
.Y(n_1054)
);

NOR3x2_ASAP7_75t_L g1055 ( 
.A(n_1047),
.B(n_851),
.C(n_98),
.Y(n_1055)
);

INVx6_ASAP7_75t_L g1056 ( 
.A(n_1041),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_SL g1057 ( 
.A(n_1046),
.B(n_97),
.C(n_100),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_1049),
.B(n_1048),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_1042),
.B(n_102),
.C(n_103),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1042),
.A2(n_734),
.B1(n_858),
.B2(n_111),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_1042),
.A2(n_105),
.B(n_106),
.C(n_112),
.Y(n_1061)
);

NAND4xp75_ASAP7_75t_L g1062 ( 
.A(n_1040),
.B(n_113),
.C(n_115),
.D(n_116),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1058),
.B(n_118),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1056),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1061),
.A2(n_119),
.B(n_122),
.C(n_123),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_1050),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1057),
.Y(n_1068)
);

CKINVDCx6p67_ASAP7_75t_R g1069 ( 
.A(n_1051),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1059),
.B(n_1056),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_1062),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1064),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1069),
.A2(n_1060),
.B1(n_1054),
.B2(n_1052),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1065),
.A2(n_1070),
.B1(n_1067),
.B2(n_1068),
.Y(n_1074)
);

XOR2x1_ASAP7_75t_L g1075 ( 
.A(n_1063),
.B(n_1055),
.Y(n_1075)
);

OA22x2_ASAP7_75t_L g1076 ( 
.A1(n_1071),
.A2(n_124),
.B1(n_130),
.B2(n_131),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_SL g1077 ( 
.A1(n_1071),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_1066),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1064),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1079),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1072),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1074),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1080),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1073),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_1075),
.B(n_1078),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1085),
.Y(n_1086)
);

NAND5xp2_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_1082),
.C(n_1076),
.D(n_1077),
.E(n_1081),
.Y(n_1087)
);

OAI222xp33_ASAP7_75t_L g1088 ( 
.A1(n_1086),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.C1(n_151),
.C2(n_152),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1087),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1088),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_1091),
.A2(n_164),
.B(n_165),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1090),
.B(n_166),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1093),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_1094)
);

AOI211xp5_ASAP7_75t_L g1095 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_172),
.C(n_173),
.Y(n_1095)
);


endmodule