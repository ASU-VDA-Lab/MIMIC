module fake_jpeg_10880_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_66),
.Y(n_68)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_42),
.B1(n_57),
.B2(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_57),
.B1(n_42),
.B2(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_76),
.B1(n_8),
.B2(n_9),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_45),
.B1(n_51),
.B2(n_54),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_65),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_49),
.B1(n_41),
.B2(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_3),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_61),
.B(n_66),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_25),
.B(n_14),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_62),
.B1(n_49),
.B2(n_64),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_97),
.B1(n_11),
.B2(n_12),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_8),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_20),
.C(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_11),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_97),
.B1(n_84),
.B2(n_96),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_72),
.B1(n_77),
.B2(n_13),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_108),
.B1(n_15),
.B2(n_16),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_24),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_111),
.B(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_117),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_95),
.C(n_88),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_37),
.C(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_108),
.C(n_105),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_102),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_123),
.A3(n_124),
.B1(n_121),
.B2(n_114),
.C1(n_104),
.C2(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_121),
.Y(n_130)
);

AOI311xp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_28),
.A3(n_30),
.B(n_31),
.C(n_35),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_99),
.B(n_36),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_105),
.Y(n_133)
);


endmodule