module fake_jpeg_14123_n_634 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_634);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_634;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx2_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_68),
.B(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_59),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_73),
.B(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_80),
.Y(n_132)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_85),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_88),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_29),
.B(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_90),
.B(n_96),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g215 ( 
.A(n_91),
.Y(n_215)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_93),
.B(n_53),
.Y(n_187)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_37),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_55),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_58),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_121),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_52),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_20),
.Y(n_186)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_23),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_49),
.B1(n_36),
.B2(n_46),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_131),
.A2(n_136),
.B1(n_144),
.B2(n_180),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_67),
.B1(n_87),
.B2(n_84),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_138),
.B(n_141),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_142),
.B(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_74),
.A2(n_36),
.B1(n_53),
.B2(n_57),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_78),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_68),
.B(n_49),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_210),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_39),
.B1(n_49),
.B2(n_46),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_164),
.A2(n_28),
.B1(n_30),
.B2(n_125),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_78),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_72),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_79),
.A2(n_30),
.B1(n_32),
.B2(n_57),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_187),
.B(n_188),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_65),
.B(n_48),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_66),
.B(n_48),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_189),
.B(n_190),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_45),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_45),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_194),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_35),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_95),
.B(n_35),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_196),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_34),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_61),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_94),
.B(n_34),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_39),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_75),
.B(n_22),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_128),
.B(n_32),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_217),
.B(n_249),
.Y(n_332)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_168),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_260),
.Y(n_295)
);

OR2x2_ASAP7_75t_SL g223 ( 
.A(n_160),
.B(n_128),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_223),
.B(n_224),
.Y(n_315)
);

INVx2_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_135),
.A2(n_91),
.B1(n_123),
.B2(n_97),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g341 ( 
.A1(n_225),
.A2(n_236),
.B1(n_258),
.B2(n_259),
.Y(n_341)
);

CKINVDCx12_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_226),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_227),
.A2(n_239),
.B1(n_150),
.B2(n_176),
.Y(n_314)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

CKINVDCx10_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_229),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_28),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_288),
.Y(n_298)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_105),
.B1(n_111),
.B2(n_107),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_237),
.B(n_270),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_83),
.B1(n_62),
.B2(n_99),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_137),
.A2(n_88),
.B1(n_98),
.B2(n_117),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_180),
.A2(n_104),
.B1(n_103),
.B2(n_122),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_131),
.A2(n_118),
.B1(n_113),
.B2(n_5),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_244),
.A2(n_257),
.B1(n_242),
.B2(n_230),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_245),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_210),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_262),
.Y(n_293)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_139),
.Y(n_252)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_132),
.B(n_4),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_254),
.B(n_255),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_155),
.B(n_157),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_140),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_154),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_212),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_278),
.Y(n_304)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_209),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_183),
.B(n_11),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_151),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_265),
.Y(n_349)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_173),
.B(n_11),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g268 ( 
.A1(n_152),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g324 ( 
.A1(n_268),
.A2(n_277),
.B1(n_286),
.B2(n_171),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_209),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_172),
.Y(n_272)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_133),
.Y(n_273)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g275 ( 
.A(n_214),
.Y(n_275)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_146),
.Y(n_276)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_210),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_133),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_281),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_202),
.A2(n_13),
.B1(n_14),
.B2(n_171),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_150),
.C(n_214),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_200),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_159),
.B(n_182),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_162),
.Y(n_310)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_269),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_153),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_285),
.B1(n_291),
.B2(n_201),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_153),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g286 ( 
.A1(n_152),
.A2(n_14),
.B1(n_198),
.B2(n_165),
.Y(n_286)
);

CKINVDCx12_ASAP7_75t_R g287 ( 
.A(n_167),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_287),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_185),
.B(n_198),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_185),
.B(n_165),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_163),
.Y(n_325)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_200),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_243),
.A2(n_143),
.B(n_204),
.C(n_151),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_301),
.B(n_327),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_309),
.B(n_323),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_314),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_248),
.A2(n_147),
.B1(n_143),
.B2(n_199),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_313),
.A2(n_339),
.B1(n_340),
.B2(n_344),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_217),
.B(n_211),
.CI(n_162),
.CON(n_316),
.SN(n_316)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_316),
.B(n_330),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_204),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_325),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_224),
.B(n_211),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_208),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_243),
.B(n_208),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_331),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_227),
.A2(n_163),
.B1(n_199),
.B2(n_179),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_333),
.A2(n_336),
.B1(n_264),
.B2(n_252),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_237),
.A2(n_179),
.B1(n_213),
.B2(n_147),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_277),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_243),
.B(n_169),
.C(n_158),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_342),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_282),
.A2(n_158),
.B1(n_176),
.B2(n_169),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_240),
.B(n_145),
.C(n_213),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_257),
.A2(n_161),
.B1(n_145),
.B2(n_149),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_246),
.B(n_161),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_350),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_244),
.A2(n_149),
.B1(n_282),
.B2(n_288),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_286),
.B1(n_229),
.B2(n_268),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_231),
.B(n_241),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_339),
.A2(n_235),
.B1(n_280),
.B2(n_290),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_353),
.A2(n_356),
.B1(n_372),
.B2(n_337),
.Y(n_403)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_354),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_298),
.A2(n_286),
.B1(n_256),
.B2(n_220),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_358),
.A2(n_300),
.B(n_342),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_329),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_349),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_362),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_232),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_361),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_306),
.Y(n_362)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_364),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_270),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_378),
.Y(n_401)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_366),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_233),
.B1(n_275),
.B2(n_245),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_368),
.A2(n_319),
.B1(n_322),
.B2(n_262),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_223),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_268),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_296),
.Y(n_375)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_268),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_379),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_305),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_293),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_395),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_350),
.B(n_332),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_277),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_385),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_317),
.B(n_277),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_386),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_286),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_390),
.Y(n_429)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx13_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_392),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_331),
.B(n_253),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_315),
.C(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_394),
.A2(n_348),
.B1(n_340),
.B2(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_294),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_293),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_396),
.B(n_328),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_400),
.B(n_417),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

BUFx12f_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_403),
.A2(n_420),
.B1(n_428),
.B2(n_391),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_352),
.A2(n_301),
.A3(n_324),
.B1(n_327),
.B2(n_297),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_424),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_407),
.A2(n_411),
.B1(n_421),
.B2(n_423),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_352),
.A2(n_297),
.B1(n_324),
.B2(n_315),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_386),
.Y(n_412)
);

INVx13_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_371),
.A2(n_293),
.B(n_338),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_415),
.A2(n_432),
.B(n_393),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_331),
.C(n_327),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_419),
.B(n_374),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_310),
.B1(n_341),
.B2(n_300),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_389),
.A2(n_218),
.B1(n_228),
.B2(n_326),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_354),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_431),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_376),
.A2(n_310),
.B1(n_311),
.B2(n_302),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_383),
.A2(n_311),
.B1(n_308),
.B2(n_303),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_379),
.Y(n_431)
);

OAI22x1_ASAP7_75t_L g435 ( 
.A1(n_377),
.A2(n_321),
.B1(n_319),
.B2(n_312),
.Y(n_435)
);

OA22x2_ASAP7_75t_L g453 ( 
.A1(n_435),
.A2(n_380),
.B1(n_396),
.B2(n_351),
.Y(n_453)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_437),
.A2(n_439),
.B1(n_442),
.B2(n_468),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_403),
.A2(n_381),
.B1(n_394),
.B2(n_385),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_460),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_429),
.A2(n_381),
.B1(n_384),
.B2(n_363),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_362),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_446),
.B(n_457),
.Y(n_476)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_426),
.Y(n_447)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_447),
.Y(n_482)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_356),
.Y(n_451)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_388),
.B(n_377),
.C(n_387),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_R g474 ( 
.A(n_453),
.B(n_435),
.Y(n_474)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_411),
.A2(n_353),
.B1(n_388),
.B2(n_391),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_459),
.B1(n_463),
.B2(n_464),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_382),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_363),
.B1(n_391),
.B2(n_351),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_462),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_375),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_418),
.B1(n_415),
.B2(n_405),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_388),
.B1(n_373),
.B2(n_370),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_360),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_465),
.B(n_469),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_466),
.A2(n_432),
.B(n_417),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_418),
.A2(n_378),
.B1(n_390),
.B2(n_326),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_413),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_470),
.B(n_430),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

NOR4xp25_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_433),
.C(n_405),
.D(n_419),
.Y(n_475)
);

NOR3xp33_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_453),
.C(n_455),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_478),
.Y(n_507)
);

OA22x2_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_435),
.B1(n_406),
.B2(n_407),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_438),
.B(n_400),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_480),
.B(n_366),
.Y(n_521)
);

OAI21x1_ASAP7_75t_SL g505 ( 
.A1(n_481),
.A2(n_450),
.B(n_448),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_404),
.C(n_423),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_491),
.C(n_492),
.Y(n_510)
);

BUFx12_ASAP7_75t_L g488 ( 
.A(n_445),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_488),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_401),
.C(n_434),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_442),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_434),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_495),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_467),
.B(n_461),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_399),
.Y(n_497)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_497),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_451),
.B(n_399),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_491),
.C(n_486),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_431),
.Y(n_501)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_501),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_445),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_398),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_468),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_453),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_SL g546 ( 
.A(n_505),
.B(n_507),
.C(n_516),
.Y(n_546)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_496),
.Y(n_506)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_506),
.Y(n_539)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_483),
.A2(n_439),
.B1(n_450),
.B2(n_452),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_509),
.A2(n_514),
.B1(n_482),
.B2(n_473),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_512),
.B(n_532),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_513),
.B(n_529),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_503),
.A2(n_421),
.B1(n_456),
.B2(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_516),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_489),
.A2(n_453),
.B(n_443),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_525),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_476),
.A2(n_449),
.B1(n_447),
.B2(n_460),
.Y(n_519)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_416),
.C(n_467),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_523),
.C(n_500),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_498),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_481),
.B(n_409),
.C(n_425),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_524),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_489),
.A2(n_398),
.B(n_454),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_526),
.Y(n_533)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_528),
.Y(n_551)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_479),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_530),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_498),
.A2(n_458),
.B1(n_441),
.B2(n_425),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_531),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_395),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_538),
.Y(n_563)
);

FAx1_ASAP7_75t_SL g537 ( 
.A(n_507),
.B(n_487),
.CI(n_474),
.CON(n_537),
.SN(n_537)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_547),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_487),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_555),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_499),
.C(n_477),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_545),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_499),
.C(n_478),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_546),
.A2(n_517),
.B(n_525),
.Y(n_557)
);

FAx1_ASAP7_75t_SL g547 ( 
.A(n_520),
.B(n_478),
.CI(n_485),
.CON(n_547),
.SN(n_547)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_478),
.C(n_485),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_549),
.B(n_554),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_471),
.C(n_482),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_521),
.B(n_471),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_529),
.B1(n_528),
.B2(n_514),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_557),
.B(n_555),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_542),
.Y(n_558)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

A2O1A1O1Ixp25_ASAP7_75t_L g559 ( 
.A1(n_535),
.A2(n_517),
.B(n_506),
.C(n_508),
.D(n_522),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_559),
.B(n_560),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_533),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_553),
.Y(n_561)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_561),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_554),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_566),
.Y(n_583)
);

BUFx12_ASAP7_75t_L g565 ( 
.A(n_537),
.Y(n_565)
);

INVx11_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_551),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_569),
.A2(n_543),
.B1(n_539),
.B2(n_540),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_515),
.C(n_504),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_570),
.B(n_572),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_509),
.C(n_518),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_536),
.A2(n_527),
.B1(n_484),
.B2(n_473),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_537),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_511),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_574),
.B(n_575),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_527),
.C(n_409),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_472),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_576),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_541),
.C(n_545),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_578),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_575),
.B(n_549),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_580),
.A2(n_588),
.B1(n_589),
.B2(n_565),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_563),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_534),
.C(n_546),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_591),
.C(n_568),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_559),
.B(n_556),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_572),
.B(n_538),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_563),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_547),
.C(n_472),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_596),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_595),
.B(n_598),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_568),
.C(n_569),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_592),
.A2(n_567),
.B(n_557),
.Y(n_597)
);

AOI31xp67_ASAP7_75t_L g611 ( 
.A1(n_597),
.A2(n_588),
.A3(n_589),
.B(n_583),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_600),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_586),
.A2(n_565),
.B1(n_547),
.B2(n_441),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_590),
.B(n_488),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_601),
.B(n_603),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_488),
.C(n_364),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_602),
.B(n_606),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_355),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_584),
.A2(n_367),
.B1(n_303),
.B2(n_307),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_605),
.A2(n_307),
.B1(n_308),
.B2(n_284),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_579),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_583),
.C(n_591),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_609),
.B(n_613),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_604),
.A2(n_582),
.B(n_592),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_610),
.A2(n_278),
.B(n_221),
.Y(n_621)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_611),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_594),
.B(n_581),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_614),
.Y(n_619)
);

AOI322xp5_ASAP7_75t_L g617 ( 
.A1(n_607),
.A2(n_597),
.A3(n_580),
.B1(n_603),
.B2(n_601),
.C1(n_392),
.C2(n_291),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_617),
.B(n_622),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_621),
.A2(n_623),
.B(n_250),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_285),
.C(n_251),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_609),
.A2(n_615),
.B(n_616),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_611),
.C(n_612),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_624),
.A2(n_626),
.B(n_627),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_618),
.Y(n_627)
);

AOI322xp5_ASAP7_75t_L g628 ( 
.A1(n_625),
.A2(n_619),
.A3(n_322),
.B1(n_345),
.B2(n_318),
.C1(n_271),
.C2(n_219),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_619),
.Y(n_630)
);

AOI322xp5_ASAP7_75t_L g631 ( 
.A1(n_630),
.A2(n_629),
.A3(n_345),
.B1(n_318),
.B2(n_276),
.C1(n_272),
.C2(n_247),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_631),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_632),
.B(n_238),
.C(n_234),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_633),
.Y(n_634)
);


endmodule