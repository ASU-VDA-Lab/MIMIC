module fake_jpeg_2239_n_497 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_133;
wire n_132;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_63),
.Y(n_143)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_74),
.Y(n_108)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_13),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_31),
.Y(n_112)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_89),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_13),
.C(n_12),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_44),
.B(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_94),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_92),
.Y(n_151)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_98),
.Y(n_124)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_116),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_31),
.B1(n_24),
.B2(n_36),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_63),
.B1(n_24),
.B2(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_34),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_18),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_59),
.B(n_18),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_46),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_38),
.B1(n_27),
.B2(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_71),
.B(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_25),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_84),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_78),
.B(n_30),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_157),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_87),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_158),
.A2(n_163),
.B1(n_169),
.B2(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_177),
.C(n_178),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_111),
.A2(n_54),
.B1(n_91),
.B2(n_96),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_33),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_199),
.Y(n_212)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_114),
.A2(n_43),
.B(n_42),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_122),
.B(n_142),
.Y(n_209)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx12_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_109),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_24),
.B1(n_65),
.B2(n_37),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_122),
.A2(n_42),
.B1(n_37),
.B2(n_43),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_15),
.B1(n_34),
.B2(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_124),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_192),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_194),
.Y(n_204)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_197),
.Y(n_207)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_110),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_108),
.B(n_98),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_201),
.Y(n_224)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_0),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_209),
.A2(n_194),
.B(n_156),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_210),
.A2(n_35),
.B1(n_178),
.B2(n_161),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_128),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_215),
.B(n_218),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_165),
.A2(n_150),
.B1(n_125),
.B2(n_110),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_169),
.B1(n_158),
.B2(n_159),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_165),
.B(n_151),
.CI(n_134),
.CON(n_218),
.SN(n_218)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_219),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_171),
.A2(n_188),
.B(n_168),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_226),
.A2(n_192),
.B(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_164),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_35),
.Y(n_258)
);

INVx4_ASAP7_75t_SL g238 ( 
.A(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_240),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_248),
.B1(n_254),
.B2(n_100),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_213),
.B(n_180),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_245),
.B(n_258),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_182),
.B1(n_184),
.B2(n_187),
.Y(n_247)
);

OAI22x1_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_263),
.B1(n_221),
.B2(n_95),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_218),
.B1(n_212),
.B2(n_213),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_202),
.C(n_189),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_266),
.C(n_205),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_160),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_257),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_252),
.B1(n_222),
.B2(n_230),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_179),
.B1(n_174),
.B2(n_199),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_218),
.A2(n_146),
.B1(n_104),
.B2(n_136),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_207),
.B(n_229),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_224),
.B(n_204),
.Y(n_271)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_215),
.B(n_170),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_262),
.Y(n_290)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_181),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_203),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_131),
.C(n_201),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_271),
.B(n_274),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_239),
.A2(n_224),
.B1(n_211),
.B2(n_216),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_279),
.B1(n_281),
.B2(n_265),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_293),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_208),
.B(n_211),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_289),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_220),
.B1(n_237),
.B2(n_233),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_220),
.B1(n_233),
.B2(n_232),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_242),
.A2(n_175),
.B1(n_196),
.B2(n_146),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_232),
.B1(n_200),
.B2(n_206),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_229),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_223),
.C(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_172),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_250),
.B1(n_259),
.B2(n_264),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_256),
.A2(n_205),
.B1(n_227),
.B2(n_225),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_225),
.B1(n_223),
.B2(n_203),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_241),
.B1(n_261),
.B2(n_246),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_296),
.A2(n_238),
.B1(n_118),
.B2(n_148),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_309),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_308),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_266),
.B(n_238),
.C(n_255),
.Y(n_302)
);

AO21x2_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_296),
.B(n_273),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_257),
.B(n_263),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_303),
.A2(n_306),
.B(n_280),
.Y(n_340)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_258),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_312),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_274),
.A2(n_243),
.B(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_240),
.B(n_103),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

AO22x1_ASAP7_75t_L g312 ( 
.A1(n_269),
.A2(n_221),
.B1(n_234),
.B2(n_227),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_246),
.Y(n_314)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_191),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_318),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_191),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_295),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_320),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_286),
.B(n_131),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_136),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_323),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_286),
.B(n_79),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_275),
.B(n_293),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_336),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_298),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_330),
.A2(n_315),
.B1(n_302),
.B2(n_312),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_284),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_344),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_332),
.B1(n_315),
.B2(n_308),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_314),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_313),
.B(n_284),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_337),
.B(n_312),
.Y(n_371)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_340),
.B(n_346),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_268),
.Y(n_342)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_287),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_318),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_288),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_166),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_319),
.A2(n_277),
.B1(n_292),
.B2(n_268),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_280),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_299),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_320),
.C(n_299),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_365),
.C(n_375),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_358),
.A2(n_366),
.B1(n_333),
.B2(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_305),
.C(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_378),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_353),
.A2(n_300),
.B1(n_315),
.B2(n_326),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_369),
.B1(n_372),
.B2(n_380),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_298),
.C(n_324),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_339),
.B1(n_333),
.B2(n_334),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_368),
.A2(n_370),
.B1(n_376),
.B2(n_377),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_328),
.A2(n_339),
.B1(n_353),
.B2(n_334),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_371),
.B(n_381),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_342),
.A2(n_302),
.B1(n_292),
.B2(n_285),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_302),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_333),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_282),
.C(n_302),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_332),
.A2(n_307),
.B1(n_282),
.B2(n_240),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_348),
.A2(n_118),
.B1(n_148),
.B2(n_142),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_354),
.B(n_10),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_342),
.A2(n_105),
.B1(n_132),
.B2(n_129),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_166),
.C(n_105),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_327),
.C(n_350),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_382),
.A2(n_340),
.B(n_333),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_384),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_406),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_389),
.A2(n_373),
.B1(n_372),
.B2(n_386),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_349),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_397),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_349),
.C(n_348),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_370),
.A2(n_336),
.B1(n_351),
.B2(n_343),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_394),
.A2(n_403),
.B1(n_404),
.B2(n_106),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_356),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_395),
.Y(n_413)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_341),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_341),
.C(n_343),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_377),
.C(n_368),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_345),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_402),
.Y(n_412)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_379),
.A2(n_345),
.B1(n_355),
.B2(n_352),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_327),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_390),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_373),
.A2(n_352),
.B(n_338),
.Y(n_406)
);

XOR2x2_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_234),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_400),
.Y(n_427)
);

BUFx12f_ASAP7_75t_SL g408 ( 
.A(n_391),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_408),
.A2(n_407),
.B(n_406),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_415),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_371),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_414),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_383),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_404),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_420),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_424),
.Y(n_440)
);

AOI322xp5_ASAP7_75t_SL g422 ( 
.A1(n_399),
.A2(n_376),
.A3(n_364),
.B1(n_380),
.B2(n_360),
.C1(n_166),
.C2(n_132),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_422),
.B(n_428),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_360),
.C(n_129),
.Y(n_424)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_426),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_411),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_106),
.C(n_115),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_388),
.C(n_401),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_430),
.B(n_441),
.Y(n_448)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_387),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_436),
.Y(n_447)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_423),
.Y(n_434)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_394),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_384),
.B(n_389),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_438),
.A2(n_442),
.B(n_61),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_428),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_419),
.A2(n_386),
.B1(n_398),
.B2(n_400),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_427),
.A2(n_398),
.B(n_127),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_444),
.A2(n_415),
.B(n_408),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_413),
.A2(n_61),
.B1(n_56),
.B2(n_115),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_446),
.A2(n_56),
.B1(n_76),
.B2(n_95),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_430),
.B(n_416),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_450),
.B(n_451),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_429),
.B(n_425),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_421),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_454),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_409),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_444),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_449),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_457),
.A2(n_459),
.B(n_455),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_459),
.A2(n_460),
.B1(n_437),
.B2(n_62),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_431),
.A2(n_76),
.B1(n_97),
.B2(n_77),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_461),
.A2(n_446),
.B1(n_441),
.B2(n_97),
.Y(n_463)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_470),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_448),
.A2(n_457),
.B(n_453),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_466),
.A2(n_471),
.B(n_462),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_443),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_472),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_443),
.C(n_437),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_SL g474 ( 
.A(n_469),
.B(n_473),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_458),
.A2(n_439),
.B(n_73),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_70),
.C(n_66),
.Y(n_473)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_476),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_57),
.B(n_51),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_477),
.A2(n_478),
.B(n_480),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_10),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_472),
.A2(n_49),
.B1(n_48),
.B2(n_28),
.Y(n_480)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g485 ( 
.A1(n_479),
.A2(n_469),
.B(n_467),
.C(n_473),
.D(n_11),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_486),
.A3(n_487),
.B1(n_483),
.B2(n_484),
.C1(n_2),
.C2(n_3),
.Y(n_489)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g486 ( 
.A1(n_482),
.A2(n_12),
.B(n_11),
.C(n_8),
.D(n_28),
.Y(n_486)
);

AOI31xp67_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_11),
.A3(n_1),
.B(n_2),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_23),
.C(n_1),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_481),
.Y(n_490)
);

AOI21xp33_ASAP7_75t_L g493 ( 
.A1(n_489),
.A2(n_491),
.B(n_3),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_490),
.A2(n_0),
.B(n_1),
.Y(n_492)
);

AOI322xp5_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_478),
.A3(n_23),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_5),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_SL g494 ( 
.A(n_492),
.B(n_493),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_4),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_4),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_496),
.B(n_4),
.Y(n_497)
);


endmodule