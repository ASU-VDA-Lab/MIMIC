module fake_jpeg_18816_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_14),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_39),
.B1(n_36),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_71)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_66),
.Y(n_78)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_1),
.B(n_2),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_71),
.B(n_10),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_56),
.B(n_60),
.C(n_3),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_5),
.C(n_6),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_76),
.B(n_65),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_11),
.B(n_12),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_80),
.A2(n_81),
.B1(n_77),
.B2(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_78),
.B(n_65),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_82),
.A3(n_18),
.B1(n_20),
.B2(n_22),
.C1(n_23),
.C2(n_24),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_15),
.B1(n_25),
.B2(n_27),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_72),
.C(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);


endmodule