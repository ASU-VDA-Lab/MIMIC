module real_jpeg_28836_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_0),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_25),
.B1(n_28),
.B2(n_55),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_25),
.B1(n_28),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_25),
.B1(n_28),
.B2(n_85),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_64),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_6),
.A2(n_64),
.B(n_134),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_11),
.B(n_25),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_6),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_42),
.B1(n_174),
.B2(n_187),
.Y(n_189)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_73),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_71),
.Y(n_179)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_12),
.A2(n_25),
.B1(n_28),
.B2(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_107),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_24),
.A2(n_37),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_24),
.A2(n_37),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_37),
.B1(n_141),
.B2(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_24),
.B(n_78),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_32),
.B(n_78),
.C(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_28),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_32),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_31),
.A2(n_65),
.A3(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_32),
.B(n_62),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_53),
.B(n_56),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_37),
.A2(n_142),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_46),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_44),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_42),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_42),
.A2(n_48),
.B1(n_179),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_43),
.B(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_43),
.A2(n_47),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_43),
.A2(n_173),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_48),
.B(n_78),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.C(n_74),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_54),
.B(n_57),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_59)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_68),
.B1(n_70),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_60),
.A2(n_68),
.B1(n_115),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_75),
.B1(n_82),
.B2(n_102),
.Y(n_101)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.CON(n_75),
.SN(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.Y(n_82)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_100),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_103),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.C(n_113),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_108),
.A2(n_109),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.C(n_118),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_202),
.B(n_208),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_153),
.B(n_201),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_143),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_127),
.B(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.C(n_139),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_128),
.A2(n_129),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_150),
.C(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_195),
.B(n_200),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_175),
.B(n_194),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_156),
.B(n_163),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_183),
.B(n_193),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_181),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_188),
.B(n_192),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);


endmodule