module fake_jpeg_15691_n_78 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

INVx11_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_1),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_38),
.B1(n_21),
.B2(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_50),
.B1(n_3),
.B2(n_5),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_58),
.Y(n_69)
);

AOI322xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.A3(n_62),
.B1(n_68),
.B2(n_63),
.C1(n_57),
.C2(n_59),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_52),
.C(n_64),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_17),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_26),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_29),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_30),
.C(n_31),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_59),
.B1(n_53),
.B2(n_57),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_53),
.Y(n_78)
);


endmodule