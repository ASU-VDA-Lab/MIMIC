module fake_jpeg_17298_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_43),
.B1(n_57),
.B2(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_84),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_0),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_48),
.B(n_49),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_58),
.C(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_54),
.B1(n_52),
.B2(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_63),
.B1(n_59),
.B2(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_42),
.Y(n_111)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_96),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_106),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_104),
.Y(n_118)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_3),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_58),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g113 ( 
.A(n_85),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_127),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_119),
.B(n_124),
.C(n_96),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_115),
.B(n_117),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_124),
.B(n_116),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_142),
.C(n_137),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_25),
.B1(n_39),
.B2(n_8),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_24),
.B(n_38),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_23),
.B(n_37),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_22),
.B(n_36),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_21),
.B(n_32),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_158),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_20),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_53),
.C(n_107),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_19),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_18),
.B(n_33),
.Y(n_163)
);


endmodule