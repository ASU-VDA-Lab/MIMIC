module fake_jpeg_16275_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_40),
.B(n_47),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_21),
.A2(n_19),
.B(n_22),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_43),
.B(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_24),
.C(n_16),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_59),
.Y(n_75)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_26),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_69),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_27),
.B1(n_19),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_74),
.B1(n_8),
.B2(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_41),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_73),
.B(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_27),
.B1(n_19),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_27),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_24),
.B1(n_16),
.B2(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_32),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_91),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_24),
.B1(n_28),
.B2(n_36),
.Y(n_112)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_32),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_15),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_18),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_36),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_8),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_18),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_12),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_109),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_127),
.B1(n_87),
.B2(n_81),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_36),
.C(n_7),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_133),
.C(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_134),
.Y(n_146)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_36),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_3),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_67),
.B(n_71),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_11),
.C(n_13),
.Y(n_133)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_135),
.B(n_80),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_104),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_82),
.A2(n_14),
.B1(n_73),
.B2(n_86),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_67),
.B1(n_71),
.B2(n_102),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_153),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_94),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_154),
.B(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_133),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_159),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_65),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_155),
.C(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_157),
.B1(n_165),
.B2(n_106),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_87),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_64),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_64),
.C(n_81),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_75),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_105),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_166),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_87),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_88),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_76),
.C(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_169),
.Y(n_183)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_139),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_76),
.C(n_78),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_90),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_117),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_114),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_114),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_110),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_111),
.C(n_110),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_110),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_165),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_117),
.B1(n_108),
.B2(n_127),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_121),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_154),
.B(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_153),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_136),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_111),
.C(n_115),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_112),
.B1(n_121),
.B2(n_119),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_171),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_119),
.B1(n_130),
.B2(n_129),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_106),
.B1(n_115),
.B2(n_95),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_161),
.B(n_154),
.C(n_144),
.D(n_151),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_203),
.B(n_205),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_193),
.B(n_195),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_151),
.C(n_140),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_204),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_174),
.C(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_175),
.B(n_156),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_160),
.B(n_146),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_219),
.B(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_147),
.B1(n_160),
.B2(n_168),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_194),
.B1(n_173),
.B2(n_134),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_176),
.B(n_145),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_145),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_107),
.B(n_136),
.Y(n_219)
);

NOR4xp25_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_181),
.C(n_178),
.D(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_230),
.C(n_212),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_215),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_203),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_233),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_187),
.C(n_179),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_107),
.B(n_125),
.C(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_223),
.B(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_205),
.B1(n_207),
.B2(n_210),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_229),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_202),
.C(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_201),
.B1(n_219),
.B2(n_206),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_245),
.B(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_200),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_212),
.C(n_213),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_253),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_242),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_223),
.B(n_224),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_254),
.B(n_255),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_227),
.B(n_235),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_231),
.Y(n_256)
);

AOI31xp67_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_240),
.A3(n_229),
.B(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_245),
.C(n_230),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_233),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_261),
.B(n_221),
.Y(n_263)
);

OAI211xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_225),
.B(n_228),
.C(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_222),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_252),
.A3(n_201),
.B1(n_221),
.B2(n_247),
.C1(n_229),
.C2(n_241),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_260),
.C(n_258),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_266),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_261),
.C(n_257),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_107),
.B(n_200),
.C(n_233),
.D(n_268),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);


endmodule