module fake_jpeg_20158_n_268 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_268);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_12),
.B(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_10),
.Y(n_35)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_12),
.B1(n_22),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_55),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_63),
.B1(n_26),
.B2(n_28),
.Y(n_75)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_65),
.Y(n_68)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_34),
.B1(n_42),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_76),
.B1(n_29),
.B2(n_13),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_34),
.B1(n_42),
.B2(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_26),
.B1(n_49),
.B2(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_84),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_55),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_48),
.B1(n_55),
.B2(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_96),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_32),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_21),
.C(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_102),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_84),
.B1(n_75),
.B2(n_76),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_66),
.B(n_79),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_26),
.B(n_29),
.C(n_28),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_54),
.B(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_29),
.B1(n_37),
.B2(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_79),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_99),
.B1(n_91),
.B2(n_16),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_115),
.B1(n_69),
.B2(n_80),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_78),
.B(n_20),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_89),
.B(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_116),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_69),
.B1(n_66),
.B2(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_99),
.B(n_70),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_139),
.B(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_129),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22x1_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_104),
.B1(n_99),
.B2(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_134),
.B1(n_146),
.B2(n_147),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_148),
.B1(n_121),
.B2(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_86),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_144),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_97),
.B1(n_100),
.B2(n_86),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_114),
.B(n_119),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_99),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_20),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_13),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_70),
.B1(n_21),
.B2(n_24),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_17),
.B1(n_16),
.B2(n_22),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_12),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_153),
.C(n_154),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_117),
.B(n_123),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_168),
.B1(n_169),
.B2(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_122),
.B1(n_17),
.B2(n_51),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_140),
.B1(n_148),
.B2(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_18),
.B(n_19),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_14),
.C(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_18),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_138),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_168),
.B(n_163),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_187),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_146),
.B1(n_147),
.B2(n_23),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_156),
.B1(n_173),
.B2(n_159),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_180),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_171),
.C(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_205),
.C(n_188),
.Y(n_212)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_163),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_179),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_210),
.B1(n_189),
.B2(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_156),
.C(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_182),
.B1(n_178),
.B2(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_224),
.B1(n_177),
.B2(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_192),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_211),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_205),
.C(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_206),
.B1(n_183),
.B2(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_185),
.B1(n_177),
.B2(n_203),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_233),
.C(n_227),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_196),
.B1(n_201),
.B2(n_191),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_241),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_191),
.B(n_6),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_245),
.B(n_7),
.Y(n_251)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_6),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_6),
.B(n_7),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_250),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_237),
.C(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_258),
.C(n_15),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_238),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_252),
.B(n_23),
.C(n_15),
.D(n_14),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g261 ( 
.A(n_259),
.B(n_256),
.C(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_15),
.C(n_23),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_262),
.B(n_23),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_23),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_14),
.B(n_3),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_265),
.A2(n_0),
.B(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_4),
.C(n_5),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_5),
.B1(n_248),
.B2(n_240),
.Y(n_268)
);


endmodule