module real_jpeg_25472_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_112, n_7, n_3, n_5, n_4, n_105, n_109, n_1, n_16, n_15, n_13, n_113, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_16;
input n_15;
input n_13;
input n_113;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_1),
.B(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_2),
.B(n_38),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_7),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_7),
.B(n_24),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_9),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_12),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_13),
.B(n_87),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_90),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_18),
.CI(n_22),
.CON(n_17),
.SN(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_97),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_21),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_21),
.B(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B(n_100),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_94),
.B(n_99),
.Y(n_31)
);

OAI321xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_86),
.A3(n_89),
.B1(n_92),
.B2(n_93),
.C(n_103),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_80),
.B(n_85),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_75),
.B(n_79),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_70),
.B(n_74),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B(n_69),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_63),
.B(n_68),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_59),
.B(n_62),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_52),
.B(n_58),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_98),
.Y(n_99)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_104),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_105),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_106),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_107),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_108),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_109),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_110),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_111),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_112),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_113),
.Y(n_91)
);


endmodule