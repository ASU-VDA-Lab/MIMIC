module fake_jpeg_4956_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_21),
.B1(n_19),
.B2(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_40),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_21),
.B(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_3),
.CI(n_5),
.CON(n_60),
.SN(n_60)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_14),
.B1(n_18),
.B2(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_27),
.C(n_31),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_24),
.C(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_1),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_57),
.B1(n_60),
.B2(n_41),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_9),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_2),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_41),
.CON(n_64),
.SN(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_56),
.B(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_46),
.B1(n_50),
.B2(n_60),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_50),
.B1(n_60),
.B2(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_44),
.B1(n_24),
.B2(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_75),
.B(n_64),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_75),
.B(n_62),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_63),
.C(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_63),
.C(n_76),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_93),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_68),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_68),
.B(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_100),
.Y(n_102)
);

NAND4xp25_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_97),
.C(n_47),
.D(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_47),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.Y(n_105)
);


endmodule