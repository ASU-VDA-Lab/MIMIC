module fake_aes_1998_n_43 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVxp67_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_0), .B(n_6), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_9), .A2(n_2), .B(n_10), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_8), .B(n_5), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_14), .B(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_11), .B(n_1), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx4_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_15), .B1(n_12), .B2(n_13), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_22), .B(n_13), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_19), .A2(n_15), .B1(n_12), .B2(n_16), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_20), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
OR2x6_ASAP7_75t_L g28 ( .A(n_25), .B(n_22), .Y(n_28) );
NAND4xp25_ASAP7_75t_L g29 ( .A(n_26), .B(n_18), .C(n_19), .D(n_21), .Y(n_29) );
NOR2x1_ASAP7_75t_R g30 ( .A(n_28), .B(n_22), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
INVxp67_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_31), .B(n_29), .Y(n_34) );
AOI311xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_28), .A3(n_21), .B(n_23), .C(n_6), .Y(n_35) );
INVxp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
NOR2xp33_ASAP7_75t_L g37 ( .A(n_33), .B(n_24), .Y(n_37) );
AOI21xp33_ASAP7_75t_SL g38 ( .A1(n_36), .A2(n_3), .B(n_7), .Y(n_38) );
OR3x2_ASAP7_75t_L g39 ( .A(n_35), .B(n_7), .C(n_37), .Y(n_39) );
INVxp67_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
AOI22xp5_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_38), .B1(n_39), .B2(n_41), .Y(n_43) );
endmodule