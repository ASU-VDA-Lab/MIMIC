module fake_jpeg_15471_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_35),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_33),
.A2(n_34),
.B1(n_21),
.B2(n_23),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_2),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_4),
.B(n_5),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_4),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_24),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_15),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_35),
.C(n_42),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_6),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_27),
.B2(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_66),
.B1(n_69),
.B2(n_76),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_46),
.B1(n_40),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_11),
.B1(n_69),
.B2(n_57),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_24),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

AO21x2_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_23),
.B(n_20),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_75),
.B1(n_54),
.B2(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_21),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_80),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_90),
.C(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_95),
.B(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_52),
.B1(n_69),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_69),
.B1(n_54),
.B2(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_73),
.B1(n_72),
.B2(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_54),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_93),
.C(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_108),
.C(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_51),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_107),
.B1(n_109),
.B2(n_99),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_95),
.B(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_102),
.B(n_108),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_78),
.C(n_86),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_85),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_112),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22x1_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_91),
.B1(n_106),
.B2(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_119),
.B1(n_108),
.B2(n_111),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_91),
.B1(n_101),
.B2(n_98),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_100),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_114),
.B(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_123),
.B(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_122),
.C(n_117),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_115),
.C(n_118),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_117),
.B1(n_121),
.B2(n_115),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B(n_129),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_130),
.A3(n_127),
.B1(n_128),
.B2(n_133),
.C(n_129),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_141)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_141),
.B(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_142),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_135),
.Y(n_145)
);


endmodule