module fake_jpeg_23925_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_0),
.Y(n_37)
);

NAND2x1_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_0),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_2),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_59),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_33),
.B1(n_29),
.B2(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_72),
.B1(n_79),
.B2(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_33),
.B1(n_29),
.B2(n_36),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_27),
.B(n_24),
.C(n_23),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_19),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_64),
.B(n_12),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_81),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_27),
.B1(n_34),
.B2(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_47),
.B1(n_43),
.B2(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_108),
.B1(n_63),
.B2(n_70),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_114),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_52),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_78),
.B(n_67),
.C(n_56),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_150),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_102),
.B1(n_119),
.B2(n_115),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_65),
.B(n_77),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_143),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_74),
.B1(n_53),
.B2(n_73),
.Y(n_138)
);

AO22x2_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_107),
.B1(n_109),
.B2(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_74),
.B1(n_53),
.B2(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_94),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_70),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_97),
.C(n_115),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_68),
.B1(n_73),
.B2(n_71),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_102),
.B1(n_119),
.B2(n_106),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_85),
.C(n_66),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_135),
.C(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_107),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_177),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_112),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_6),
.B(n_7),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_149),
.Y(n_178)
);

AOI22x1_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_76),
.B1(n_111),
.B2(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_159),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_116),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_168),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_150),
.B1(n_137),
.B2(n_127),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_95),
.B1(n_93),
.B2(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_95),
.B1(n_93),
.B2(n_13),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_187),
.C(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_189),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_141),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_195),
.B1(n_176),
.B2(n_155),
.C(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_129),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_126),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_122),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_171),
.B1(n_163),
.B2(n_181),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_210),
.B1(n_212),
.B2(n_199),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_166),
.B(n_171),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_206),
.B(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_208),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_172),
.B1(n_155),
.B2(n_177),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_213),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_195),
.A2(n_188),
.B(n_172),
.C(n_169),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_217),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_179),
.C(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_227),
.C(n_153),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

OA21x2_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_210),
.B(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_218),
.B1(n_228),
.B2(n_224),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_162),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_153),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_136),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_136),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_234),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_223),
.C(n_225),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_215),
.B(n_219),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_216),
.C(n_124),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_245),
.Y(n_253)
);

XOR2x1_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_227),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_231),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_221),
.B(n_230),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_131),
.Y(n_256)
);

OAI321xp33_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_246),
.A3(n_244),
.B1(n_241),
.B2(n_240),
.C(n_15),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_14),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_252),
.C(n_12),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_254),
.CI(n_257),
.CON(n_261),
.SN(n_261)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_14),
.B(n_15),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_262),
.B(n_260),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_258),
.Y(n_264)
);


endmodule