module fake_jpeg_14358_n_433 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_433);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_45),
.B(n_52),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_57),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_70),
.Y(n_112)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_35),
.Y(n_121)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_25),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_36),
.Y(n_115)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_81),
.Y(n_110)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_25),
.B1(n_40),
.B2(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_87),
.A2(n_95),
.B1(n_107),
.B2(n_137),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_42),
.B1(n_24),
.B2(n_33),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_94),
.B1(n_109),
.B2(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_36),
.B(n_42),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_92),
.B(n_37),
.CI(n_3),
.CON(n_164),
.SN(n_164)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_42),
.B1(n_24),
.B2(n_33),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_39),
.B1(n_31),
.B2(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_40),
.B1(n_38),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_130),
.B1(n_78),
.B2(n_63),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_42),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_121),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_61),
.B1(n_69),
.B2(n_56),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_33),
.B1(n_31),
.B2(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_30),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_27),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_116),
.B(n_117),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_26),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_43),
.B(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_134),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_54),
.A2(n_31),
.B1(n_39),
.B2(n_22),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_37),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_62),
.A2(n_39),
.B1(n_31),
.B2(n_37),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_37),
.B1(n_16),
.B2(n_5),
.Y(n_137)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_51),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_140),
.B(n_141),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_83),
.B(n_81),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_142),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_75),
.B(n_64),
.C(n_49),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_143),
.A2(n_149),
.B(n_146),
.C(n_181),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_144),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_212)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_132),
.B1(n_114),
.B2(n_123),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_148),
.A2(n_164),
.B(n_146),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_92),
.A2(n_77),
.B1(n_59),
.B2(n_46),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_150),
.B(n_156),
.Y(n_218)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_151),
.Y(n_220)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_152),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_101),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_160),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_37),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_162),
.B(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_2),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_169),
.B(n_184),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_174),
.Y(n_234)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_130),
.B1(n_131),
.B2(n_128),
.Y(n_192)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_179),
.Y(n_203)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_180),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_183),
.Y(n_229)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_84),
.B(n_3),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_110),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_188),
.Y(n_193)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_96),
.B(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_6),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_98),
.B(n_6),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_191),
.B1(n_160),
.B2(n_159),
.Y(n_221)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_91),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_188),
.B1(n_154),
.B2(n_153),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_194),
.A2(n_211),
.B(n_234),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_196),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_122),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_201),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_105),
.B1(n_131),
.B2(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_198),
.A2(n_212),
.B1(n_226),
.B2(n_230),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_129),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_214),
.C(n_233),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_136),
.B(n_129),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_205),
.A2(n_213),
.B(n_215),
.Y(n_244)
);

AOI22x1_ASAP7_75t_L g211 ( 
.A1(n_149),
.A2(n_105),
.B1(n_136),
.B2(n_9),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_148),
.A2(n_10),
.B(n_11),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_139),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_172),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_12),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_164),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_149),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_177),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_178),
.B1(n_138),
.B2(n_191),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_143),
.B(n_142),
.C(n_145),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_152),
.C(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_258),
.B1(n_274),
.B2(n_278),
.Y(n_285)
);

OAI22x1_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_143),
.B1(n_183),
.B2(n_179),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_254),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_143),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_249),
.B(n_266),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_248),
.B1(n_260),
.B2(n_262),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_185),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_259),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_192),
.A2(n_182),
.B1(n_173),
.B2(n_180),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_159),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_174),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_272),
.B(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_197),
.B(n_170),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_249),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_230),
.B1(n_215),
.B2(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_206),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_193),
.B1(n_211),
.B2(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_214),
.C(n_193),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_250),
.C(n_259),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_211),
.A2(n_216),
.B1(n_213),
.B2(n_203),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_203),
.A2(n_237),
.B1(n_196),
.B2(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_275),
.B1(n_248),
.B2(n_246),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_273),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_221),
.A2(n_227),
.B1(n_235),
.B2(n_199),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_202),
.A2(n_234),
.B1(n_225),
.B2(n_195),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_232),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_204),
.B1(n_220),
.B2(n_231),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_195),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_276),
.B(n_279),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_204),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_199),
.A2(n_228),
.B1(n_230),
.B2(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_224),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_283),
.A2(n_303),
.B1(n_310),
.B2(n_280),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_257),
.B(n_255),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_298),
.C(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_274),
.B1(n_270),
.B2(n_245),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_305),
.B1(n_285),
.B2(n_301),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_255),
.A2(n_245),
.B(n_266),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_301),
.B(n_294),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_261),
.C(n_250),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_256),
.C(n_244),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_260),
.B(n_242),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_304),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_251),
.A2(n_274),
.B1(n_264),
.B2(n_267),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_277),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_270),
.B1(n_278),
.B2(n_241),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_267),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_275),
.B(n_240),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_312),
.C(n_291),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_247),
.B1(n_268),
.B2(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_249),
.B(n_252),
.C(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_316),
.B(n_342),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_324),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_318),
.A2(n_326),
.B1(n_332),
.B2(n_287),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_282),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_307),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_330),
.Y(n_357)
);

OAI22x1_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_285),
.B1(n_305),
.B2(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_331),
.C(n_325),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_293),
.C(n_306),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_294),
.C(n_288),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_303),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_308),
.A2(n_296),
.B1(n_280),
.B2(n_297),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_333),
.A2(n_338),
.B1(n_309),
.B2(n_313),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_284),
.B(n_290),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_335),
.Y(n_365)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_314),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_336),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_337),
.A2(n_287),
.B(n_316),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_288),
.B1(n_297),
.B2(n_302),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_286),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g349 ( 
.A(n_339),
.B(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_343),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_314),
.B(n_312),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_345),
.C(n_346),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_299),
.C(n_309),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_318),
.B1(n_332),
.B2(n_320),
.Y(n_373)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_338),
.B(n_333),
.Y(n_367)
);

INVx13_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_327),
.C(n_322),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_357),
.C(n_363),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_339),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_361),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_343),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_331),
.C(n_337),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_340),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_319),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_354),
.B(n_361),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_326),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_374),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_366),
.B(n_329),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_370),
.B(n_378),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_372),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_352),
.B1(n_353),
.B2(n_358),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_319),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_320),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_379),
.C(n_380),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_341),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_357),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_323),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_347),
.A2(n_335),
.B1(n_348),
.B2(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_384),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_362),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_344),
.B(n_362),
.Y(n_385)
);

XOR2x1_ASAP7_75t_SL g397 ( 
.A(n_385),
.B(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_387),
.A2(n_375),
.B(n_390),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_353),
.B1(n_359),
.B2(n_344),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_389),
.Y(n_406)
);

OAI321xp33_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_359),
.A3(n_365),
.B1(n_355),
.B2(n_349),
.C(n_360),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_355),
.B(n_365),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_390),
.A2(n_401),
.B(n_391),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g392 ( 
.A1(n_381),
.A2(n_369),
.A3(n_383),
.B1(n_370),
.B2(n_351),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_398),
.Y(n_408)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_394),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_351),
.C(n_360),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_399),
.C(n_393),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_397),
.B(n_398),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_369),
.A2(n_376),
.B1(n_368),
.B2(n_374),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_375),
.C(n_377),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_401),
.A2(n_385),
.B1(n_380),
.B2(n_371),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_402),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_409),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_410),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_405),
.A2(n_386),
.B(n_389),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_393),
.C(n_395),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_388),
.C(n_400),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_413),
.A2(n_415),
.B(n_417),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_406),
.A2(n_391),
.B(n_397),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_400),
.C(n_387),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_408),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_420),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_414),
.A2(n_406),
.B1(n_411),
.B2(n_407),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_405),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_422),
.A2(n_423),
.B(n_413),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_410),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_424),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g426 ( 
.A1(n_419),
.A2(n_404),
.B(n_416),
.C(n_392),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_SL g428 ( 
.A(n_426),
.B(n_407),
.C(n_408),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_425),
.B(n_421),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_427),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_423),
.C(n_416),
.Y(n_431)
);

BUFx24_ASAP7_75t_SL g432 ( 
.A(n_431),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_432),
.B(n_396),
.Y(n_433)
);


endmodule