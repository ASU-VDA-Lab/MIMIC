module fake_ariane_385_n_4866 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_4866);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_4866;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4688;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4834;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_4770;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_4586;
wire n_1469;
wire n_4342;
wire n_4692;
wire n_4557;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2334;
wire n_2135;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_4475;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_610;
wire n_4403;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_1430;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_4626;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_4178;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4547;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_4058;
wire n_952;
wire n_864;
wire n_4090;
wire n_2446;
wire n_4819;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_4813;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2461;
wire n_2207;
wire n_2702;
wire n_3719;
wire n_4363;
wire n_2731;
wire n_3703;
wire n_634;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_2238;
wire n_1503;
wire n_2529;
wire n_2374;
wire n_4103;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_1181;
wire n_3435;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_4841;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_4683;
wire n_737;
wire n_2873;
wire n_2653;
wire n_1298;
wire n_1745;
wire n_4610;
wire n_1366;
wire n_4674;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_4028;
wire n_4796;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_4736;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_4842;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_4416;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4439;
wire n_870;
wire n_2547;
wire n_4600;
wire n_3382;
wire n_1453;
wire n_945;
wire n_958;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_4575;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_813;
wire n_4660;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4106;
wire n_4853;
wire n_4589;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_4581;
wire n_2960;
wire n_4260;
wire n_665;
wire n_754;
wire n_4625;
wire n_3270;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_829;
wire n_1761;
wire n_4148;
wire n_4814;
wire n_1062;
wire n_4845;
wire n_738;
wire n_3679;
wire n_4702;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_4512;
wire n_2342;
wire n_4590;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_4038;
wire n_3856;
wire n_4132;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_4500;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_4734;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_4722;
wire n_2914;
wire n_4824;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_4515;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3890;
wire n_4741;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_4136;
wire n_4604;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4567;
wire n_4176;
wire n_1207;
wire n_4760;
wire n_4124;
wire n_3606;
wire n_786;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_4797;
wire n_4823;
wire n_3474;
wire n_2232;
wire n_4488;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_4831;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_1512;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_4782;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_4608;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_4597;
wire n_4560;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_3948;
wire n_4621;
wire n_4839;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_4546;
wire n_1889;
wire n_587;
wire n_1977;
wire n_4768;
wire n_2650;
wire n_693;
wire n_863;
wire n_1254;
wire n_3960;
wire n_4454;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_611;
wire n_2060;
wire n_1295;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_3883;
wire n_1013;
wire n_4576;
wire n_4032;
wire n_4018;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_661;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_3003;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_4572;
wire n_4505;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_3739;
wire n_3962;
wire n_1597;
wire n_4082;
wire n_4476;
wire n_2942;
wire n_4680;
wire n_1771;
wire n_2902;
wire n_4541;
wire n_4360;
wire n_1544;
wire n_579;
wire n_3271;
wire n_4540;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_2382;
wire n_1213;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_4443;
wire n_1021;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_4854;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_4815;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_4665;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_4593;
wire n_942;
wire n_4562;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_2909;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_3554;
wire n_4276;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_4747;
wire n_1830;
wire n_3850;
wire n_4529;
wire n_575;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_4498;
wire n_772;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_4432;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_4495;
wire n_2800;
wire n_2568;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_4737;
wire n_4801;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_4109;
wire n_3777;
wire n_4108;
wire n_4502;
wire n_4530;
wire n_4774;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_4740;
wire n_3588;
wire n_1108;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_4115;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_652;
wire n_1819;
wire n_4850;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_4513;
wire n_1179;
wire n_4311;
wire n_3284;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_696;
wire n_4775;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_4827;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_4786;
wire n_2791;
wire n_762;
wire n_1468;
wire n_1253;
wire n_1661;
wire n_4378;
wire n_555;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_4459;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_4594;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_4709;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4642;
wire n_4233;
wire n_3538;
wire n_4791;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_4718;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_4029;
wire n_3875;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_4794;
wire n_2745;
wire n_4843;
wire n_2087;
wire n_669;
wire n_1491;
wire n_2628;
wire n_931;
wire n_3219;
wire n_3362;
wire n_619;
wire n_967;
wire n_1083;
wire n_3937;
wire n_4130;
wire n_4763;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_746;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_615;
wire n_4587;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_4456;
wire n_4795;
wire n_4838;
wire n_1312;
wire n_4508;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2601;
wire n_2172;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_815;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_2668;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_3257;
wire n_650;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2557;
wire n_2898;
wire n_2695;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_712;
wire n_3567;
wire n_909;
wire n_4003;
wire n_1392;
wire n_767;
wire n_2795;
wire n_1832;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_4438;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_3884;
wire n_4433;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_4492;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_965;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_4806;
wire n_4861;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_4445;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_4254;
wire n_4462;
wire n_2507;
wire n_4219;
wire n_4484;
wire n_3438;
wire n_4723;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_4451;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_3661;
wire n_2223;
wire n_3082;
wire n_836;
wire n_1279;
wire n_3415;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_4784;
wire n_1247;
wire n_4234;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_2632;
wire n_1255;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_4613;
wire n_4836;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_3971;
wire n_4315;
wire n_706;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_4442;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_4857;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_4494;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_4207;
wire n_3711;
wire n_4201;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_4725;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_4719;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_4751;
wire n_3994;
wire n_4636;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_4563;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_4049;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_4522;
wire n_2718;
wire n_4263;
wire n_720;
wire n_4707;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_4426;
wire n_3876;
wire n_4588;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_4634;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_4658;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4186;
wire n_1501;
wire n_4089;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_4699;
wire n_1198;
wire n_4096;
wire n_4506;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_4728;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_4643;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_4713;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_4543;
wire n_4788;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_4818;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_4555;
wire n_1901;
wire n_647;
wire n_2055;
wire n_4486;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_600;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_4441;
wire n_1906;
wire n_4323;
wire n_3039;
wire n_1899;
wire n_2195;
wire n_3922;
wire n_4447;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_4640;
wire n_1467;
wire n_4780;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_4458;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_4523;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_604;
wire n_677;
wire n_3705;
wire n_3022;
wire n_703;
wire n_3983;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_681;
wire n_3477;
wire n_3286;
wire n_4480;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_707;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_4583;
wire n_3788;
wire n_3939;
wire n_590;
wire n_2075;
wire n_699;
wire n_727;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3837;
wire n_3835;
wire n_1015;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2418;
wire n_3260;
wire n_3349;
wire n_3819;
wire n_3761;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_4348;
wire n_1602;
wire n_4616;
wire n_688;
wire n_4771;
wire n_4457;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_4773;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3205;
wire n_3051;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_729;
wire n_3403;
wire n_887;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_4661;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_4856;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_1402;
wire n_957;
wire n_1242;
wire n_3957;
wire n_2754;
wire n_2774;
wire n_2707;
wire n_4580;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_4826;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_861;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_877;
wire n_3995;
wire n_1119;
wire n_4460;
wire n_3713;
wire n_4670;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_4798;
wire n_4648;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_4848;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4461;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_4615;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_4844;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_2949;
wire n_888;
wire n_2894;
wire n_2300;
wire n_845;
wire n_3896;
wire n_4067;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_4551;
wire n_3214;
wire n_551;
wire n_3551;
wire n_4521;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_4677;
wire n_1844;
wire n_4525;
wire n_2283;
wire n_582;
wire n_2526;
wire n_3364;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_710;
wire n_2994;
wire n_1919;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_4324;
wire n_842;
wire n_3626;
wire n_1898;
wire n_4428;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_4598;
wire n_4729;
wire n_4464;
wire n_4463;
wire n_1793;
wire n_4446;
wire n_4789;
wire n_3180;
wire n_3648;
wire n_4662;
wire n_3423;
wire n_4800;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_742;
wire n_1388;
wire n_2119;
wire n_1266;
wire n_1719;
wire n_2742;
wire n_1540;
wire n_769;
wire n_3671;
wire n_4396;
wire n_4440;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_4425;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_4565;
wire n_744;
wire n_2821;
wire n_3491;
wire n_1895;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_4781;
wire n_3064;
wire n_2904;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_4828;
wire n_1860;
wire n_1734;
wire n_3065;
wire n_4652;
wire n_3016;
wire n_4114;
wire n_4552;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_837;
wire n_812;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_4482;
wire n_2480;
wire n_606;
wire n_3024;
wire n_951;
wire n_4528;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_4863;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4859;
wire n_4568;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_4811;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4424;
wire n_4429;
wire n_3340;
wire n_4351;
wire n_4192;
wire n_4779;
wire n_2140;
wire n_1748;
wire n_873;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_4524;
wire n_1538;
wire n_4865;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_4646;
wire n_4657;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_4436;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_4545;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_4758;
wire n_3685;
wire n_4840;
wire n_811;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_624;
wire n_3507;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_4535;
wire n_2492;
wire n_3864;
wire n_4694;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_4664;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_2265;
wire n_687;
wire n_4633;
wire n_4708;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_2627;
wire n_1786;
wire n_4050;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_642;
wire n_2106;
wire n_1804;
wire n_1406;
wire n_4717;
wire n_595;
wire n_4306;
wire n_4739;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_4671;
wire n_2272;
wire n_3266;
wire n_4766;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_4558;
wire n_1318;
wire n_854;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_805;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4511;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_4675;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1856;
wire n_1476;
wire n_1733;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_1524;
wire n_3925;
wire n_2928;
wire n_4651;
wire n_4689;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_4748;
wire n_961;
wire n_4537;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_4618;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_4847;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_4846;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_2295;
wire n_4076;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_4704;
wire n_3129;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_4427;
wire n_4805;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1324;
wire n_2528;
wire n_1778;
wire n_3640;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4822;
wire n_686;
wire n_4279;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1759;
wire n_1557;
wire n_2325;
wire n_1829;
wire n_4330;
wire n_1130;
wire n_4635;
wire n_4724;
wire n_1450;
wire n_4152;
wire n_4744;
wire n_3718;
wire n_4706;
wire n_2022;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_4666;
wire n_4764;
wire n_4783;
wire n_3017;
wire n_2986;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_2546;
wire n_2890;
wire n_3381;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_897;
wire n_3455;
wire n_807;
wire n_949;
wire n_3736;
wire n_4466;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_2760;
wire n_1864;
wire n_3907;
wire n_4603;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4419;
wire n_4835;
wire n_1151;
wire n_4595;
wire n_554;
wire n_960;
wire n_4420;
wire n_4703;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3605;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_4721;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4404;
wire n_4742;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_4630;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_4829;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_4617;
wire n_818;
wire n_4377;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_4790;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4732;
wire n_4301;
wire n_3573;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_4727;
wire n_1303;
wire n_4561;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_4641;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_2610;
wire n_1593;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_4825;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_4712;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_2804;
wire n_1288;
wire n_2475;
wire n_1185;
wire n_858;
wire n_2173;
wire n_3982;
wire n_4715;
wire n_4817;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_4755;
wire n_2771;
wire n_4799;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_4202;
wire n_4536;
wire n_2044;
wire n_4534;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_4437;
wire n_1192;
wire n_3738;
wire n_3098;
wire n_894;
wire n_1380;
wire n_4503;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_562;
wire n_4070;
wire n_2020;
wire n_748;
wire n_3987;
wire n_2310;
wire n_4249;
wire n_4418;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_4769;
wire n_914;
wire n_4582;
wire n_689;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_4450;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_4412;
wire n_576;
wire n_843;
wire n_2647;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4370;
wire n_3444;
wire n_4368;
wire n_4682;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_4816;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_4184;
wire n_846;
wire n_4430;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_4810;
wire n_2450;
wire n_2411;
wire n_4631;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1955;
wire n_1504;
wire n_2431;
wire n_2110;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3322;
wire n_2666;
wire n_3289;
wire n_4538;
wire n_4544;
wire n_1370;
wire n_1603;
wire n_728;
wire n_4191;
wire n_4409;
wire n_4478;
wire n_2935;
wire n_2401;
wire n_4246;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_4355;
wire n_2863;
wire n_2588;
wire n_2331;
wire n_4632;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_4061;
wire n_2658;
wire n_623;
wire n_3587;
wire n_3509;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_4601;
wire n_3344;
wire n_4754;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_4531;
wire n_4155;
wire n_3376;
wire n_810;
wire n_4278;
wire n_4518;
wire n_4710;
wire n_1959;
wire n_1290;
wire n_3770;
wire n_3497;
wire n_617;
wire n_4375;
wire n_4542;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_4532;
wire n_4685;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_4684;
wire n_743;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_3790;
wire n_4711;
wire n_907;
wire n_2749;
wire n_2592;
wire n_1454;
wire n_660;
wire n_3490;
wire n_2459;
wire n_962;
wire n_4413;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2751;
wire n_2566;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_3251;
wire n_673;
wire n_3288;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_571;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_4821;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_4650;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_4164;
wire n_4126;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_3363;
wire n_1994;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_3836;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_4860;
wire n_4469;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_4455;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4366;
wire n_1584;
wire n_1157;
wire n_4384;
wire n_848;
wire n_4639;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_4733;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_1814;
wire n_4210;
wire n_4577;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_692;
wire n_4208;
wire n_3442;
wire n_3972;
wire n_2054;
wire n_4623;
wire n_2315;
wire n_1857;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_4509;
wire n_2073;
wire n_2150;
wire n_4481;
wire n_4004;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_621;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_4804;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_4669;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_585;
wire n_3092;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_875;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_622;
wire n_1626;
wire n_3436;
wire n_4620;
wire n_4584;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_4759;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_3751;
wire n_2299;
wire n_4388;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_4477;
wire n_1621;
wire n_4110;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_4411;
wire n_1221;
wire n_4217;
wire n_4585;
wire n_1785;
wire n_792;
wire n_1262;
wire n_4271;
wire n_1942;
wire n_3406;
wire n_2180;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_580;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_4687;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_4785;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_4605;
wire n_4720;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_4649;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_2465;
wire n_3610;
wire n_1407;
wire n_2865;
wire n_1204;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_4762;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_4592;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_3677;
wire n_2010;
wire n_1564;
wire n_4832;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_4820;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4644;
wire n_4086;
wire n_4752;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_4746;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_4656;
wire n_4862;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_4672;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_653;
wire n_1445;
wire n_3034;
wire n_1317;
wire n_4858;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_4435;
wire n_783;
wire n_4778;
wire n_4053;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_4750;
wire n_3177;
wire n_4667;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_4496;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_4596;
wire n_4673;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_4628;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_4837;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_788;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_4738;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_4554;
wire n_2630;
wire n_591;
wire n_4105;
wire n_4526;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_1663;
wire n_3114;
wire n_919;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_4578;
wire n_1458;
wire n_679;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_3360;
wire n_4470;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_2787;
wire n_765;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_4659;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2556;
wire n_2440;
wire n_2186;
wire n_2215;
wire n_1530;
wire n_4057;
wire n_2770;
wire n_4550;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4647;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_4144;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_2012;
wire n_1937;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_4849;
wire n_4726;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_733;
wire n_2212;
wire n_761;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_4434;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_4499;
wire n_2569;
wire n_758;
wire n_4504;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_2897;
wire n_816;
wire n_4339;
wire n_1322;
wire n_3273;
wire n_4812;
wire n_4497;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_4510;
wire n_835;
wire n_3155;
wire n_4855;
wire n_4300;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4169;
wire n_4024;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4472;
wire n_4253;
wire n_1865;
wire n_1710;
wire n_2641;
wire n_2522;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_1792;
wire n_4064;
wire n_3351;
wire n_2062;
wire n_4489;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_4519;
wire n_1099;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_4564;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_4787;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_4681;
wire n_3778;
wire n_4654;
wire n_831;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_4566;
wire n_3970;
wire n_4371;
wire n_778;
wire n_2351;
wire n_1619;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_2784;
wire n_1902;
wire n_3898;
wire n_4414;
wire n_2541;
wire n_694;
wire n_1643;
wire n_4185;
wire n_3188;
wire n_3232;
wire n_3001;
wire n_1320;
wire n_4448;
wire n_1113;
wire n_4749;
wire n_3218;
wire n_2347;
wire n_4676;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_2538;
wire n_1845;
wire n_4295;
wire n_3932;
wire n_2101;
wire n_2577;
wire n_1934;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_4579;
wire n_4507;
wire n_2104;
wire n_4756;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_2552;
wire n_671;
wire n_1533;
wire n_2372;
wire n_1470;
wire n_1806;
wire n_3445;
wire n_4087;
wire n_4776;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_4473;
wire n_4619;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_4471;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_904;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_4691;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_4449;
wire n_3285;
wire n_3824;
wire n_4607;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_4753;
wire n_1150;
wire n_4266;
wire n_977;
wire n_2339;
wire n_3846;
wire n_4803;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_4407;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4373;
wire n_2472;
wire n_4695;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_4479;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_4668;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_4777;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_4743;
wire n_3371;
wire n_1781;
wire n_4571;
wire n_709;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_809;
wire n_3194;
wire n_3143;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_4415;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_3461;
wire n_3366;
wire n_2430;
wire n_2504;
wire n_910;
wire n_4211;
wire n_3094;
wire n_939;
wire n_1410;
wire n_2297;
wire n_741;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4700;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_4679;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_4408;
wire n_1983;
wire n_2982;
wire n_1273;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_4767;
wire n_2913;
wire n_993;
wire n_4569;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_4483;
wire n_3672;
wire n_922;
wire n_1004;
wire n_3061;
wire n_1810;
wire n_2587;
wire n_3504;
wire n_2839;
wire n_1347;
wire n_4693;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_4548;
wire n_4487;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_4807;
wire n_3556;
wire n_4539;
wire n_896;
wire n_4574;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_4698;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_3918;
wire n_716;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_4501;
wire n_4808;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_3244;
wire n_4383;
wire n_4830;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_596;
wire n_3112;
wire n_2051;
wire n_954;
wire n_1821;
wire n_1168;
wire n_4095;
wire n_4444;
wire n_4663;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_4624;
wire n_4485;
wire n_656;
wire n_574;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_4678;
wire n_2585;
wire n_1591;
wire n_664;
wire n_3293;
wire n_2995;
wire n_3361;
wire n_4533;
wire n_4287;
wire n_1683;
wire n_2582;
wire n_1229;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_4686;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3895;
wire n_3779;
wire n_4627;
wire n_3149;
wire n_1063;
wire n_4761;
wire n_3934;
wire n_4556;
wire n_991;
wire n_2205;
wire n_2275;
wire n_2183;
wire n_4338;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_4606;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_4573;
wire n_938;
wire n_1891;
wire n_4520;
wire n_1328;
wire n_895;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_3058;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_2792;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_4553;
wire n_4465;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3592;
wire n_3557;
wire n_3725;
wire n_3986;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_937;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_4772;
wire n_4612;
wire n_4852;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_3128;
wire n_1827;
wire n_4149;
wire n_4120;
wire n_866;
wire n_925;
wire n_4335;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2880;
wire n_2819;
wire n_3075;
wire n_3030;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_4614;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_4629;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_4516;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_4716;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_4730;
wire n_773;
wire n_3221;
wire n_2798;
wire n_2316;
wire n_3217;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_4599;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4622;
wire n_4222;
wire n_803;
wire n_2514;
wire n_1871;
wire n_718;
wire n_4757;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_3249;
wire n_1870;
wire n_3430;
wire n_3483;
wire n_4591;
wire n_4046;
wire n_4467;
wire n_4701;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_782;
wire n_3489;
wire n_3083;
wire n_4570;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_4696;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_4655;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_3041;
wire n_1989;
wire n_1421;
wire n_2423;
wire n_2689;
wire n_2208;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_4493;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_4645;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_4851;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_2345;
wire n_4417;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx3_ASAP7_75t_L g550 ( 
.A(n_158),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_193),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_71),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_239),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_192),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_278),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_511),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_17),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_11),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_411),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_294),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_158),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_407),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_498),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_543),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_200),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_405),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_430),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_248),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_202),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_390),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_278),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_478),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_456),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_517),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_534),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_338),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_269),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_352),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_196),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_371),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_25),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_287),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_402),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_0),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_124),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_331),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_184),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_147),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_387),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_208),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_222),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_488),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_110),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_376),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_183),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_360),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_40),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g600 ( 
.A(n_24),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_213),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_62),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_84),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_96),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_380),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_419),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_83),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_504),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_383),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_546),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_139),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_525),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_166),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_174),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_208),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_404),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_410),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_118),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_439),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_394),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_329),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_60),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_1),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_418),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_78),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_59),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_129),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_81),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_224),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_130),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_16),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_440),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_23),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_70),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_300),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_378),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_363),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_444),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_391),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_120),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_140),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_400),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_522),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_81),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_62),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_523),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_309),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_362),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_114),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_279),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_449),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_457),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_540),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_239),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_248),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_389),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_77),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_489),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_331),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_136),
.Y(n_665)
);

INVxp33_ASAP7_75t_SL g666 ( 
.A(n_146),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_15),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_9),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_539),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_434),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_431),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_5),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_520),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_191),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_279),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_184),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_225),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_24),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_367),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_108),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_283),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_265),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_526),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_75),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_379),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_61),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_35),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_85),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_312),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_103),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_460),
.Y(n_691)
);

CKINVDCx16_ASAP7_75t_R g692 ( 
.A(n_502),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_284),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_438),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_353),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_267),
.Y(n_696)
);

BUFx5_ASAP7_75t_L g697 ( 
.A(n_55),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_521),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_61),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_269),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_417),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_509),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_51),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_117),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_166),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_13),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_209),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_386),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_134),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_157),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_253),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_204),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_39),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_13),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_263),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_76),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_226),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_464),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_194),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_251),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_188),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_392),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_441),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_506),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_510),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_313),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_255),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_427),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_480),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_277),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_335),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_263),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_393),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_530),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_547),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_151),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_109),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_133),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_433),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_200),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_108),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_178),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_341),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_235),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_219),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_254),
.Y(n_746)
);

CKINVDCx14_ASAP7_75t_R g747 ( 
.A(n_225),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_533),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_381),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_538),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_496),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_145),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_80),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_544),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_280),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_162),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_157),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_518),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_537),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_320),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_58),
.Y(n_761)
);

CKINVDCx11_ASAP7_75t_R g762 ( 
.A(n_507),
.Y(n_762)
);

BUFx2_ASAP7_75t_SL g763 ( 
.A(n_43),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_372),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_428),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_177),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_243),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_211),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_466),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_532),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_467),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_227),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_542),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_297),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_396),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_205),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_458),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_30),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_188),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_406),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_290),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_448),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_535),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_107),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_19),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_334),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_485),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_531),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_293),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_315),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_515),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_349),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_416),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_38),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_357),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_27),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_343),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_337),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_499),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_462),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_275),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_334),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_260),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_179),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_32),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_20),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_297),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_167),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_28),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_476),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_314),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_527),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_354),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_60),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_126),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_365),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_129),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_329),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_463),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_92),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_186),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_281),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_217),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_491),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_377),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_103),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_253),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_133),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_55),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_1),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_296),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_210),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_70),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_58),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_174),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_173),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_270),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_3),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_123),
.Y(n_839)
);

BUFx2_ASAP7_75t_SL g840 ( 
.A(n_49),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_106),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_326),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_505),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_176),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_548),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_280),
.Y(n_846)
);

CKINVDCx14_ASAP7_75t_R g847 ( 
.A(n_172),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_89),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_83),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_113),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_319),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_162),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_374),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_333),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_134),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_146),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_274),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_306),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_241),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_194),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_259),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_170),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_337),
.Y(n_863)
);

BUFx10_ASAP7_75t_L g864 ( 
.A(n_483),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_345),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_26),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_370),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_204),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_541),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_351),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_210),
.Y(n_871)
);

CKINVDCx14_ASAP7_75t_R g872 ( 
.A(n_136),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_295),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_176),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_294),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_119),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_202),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_395),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_501),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_26),
.Y(n_880)
);

BUFx10_ASAP7_75t_L g881 ( 
.A(n_549),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_164),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_182),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_469),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_88),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_209),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_185),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_302),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_255),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_254),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_29),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_459),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_151),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_109),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_484),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_481),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_282),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_99),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_412),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_312),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_322),
.Y(n_901)
);

BUFx5_ASAP7_75t_L g902 ( 
.A(n_453),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_59),
.Y(n_903)
);

CKINVDCx16_ASAP7_75t_R g904 ( 
.A(n_375),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_142),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_63),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_86),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_10),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_69),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_23),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_179),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_126),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_235),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_167),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_322),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_9),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_110),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_508),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_116),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_273),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_524),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_317),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_149),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_432),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_189),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_293),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_445),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_119),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_274),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_173),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_138),
.Y(n_931)
);

CKINVDCx14_ASAP7_75t_R g932 ( 
.A(n_226),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_35),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_320),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_88),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_358),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_536),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_165),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_319),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_369),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_54),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_528),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_177),
.Y(n_943)
);

CKINVDCx16_ASAP7_75t_R g944 ( 
.A(n_332),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_295),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_398),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_308),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_63),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_333),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_106),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_170),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_339),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_5),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_53),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_513),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_172),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_291),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_425),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_205),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_261),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_91),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_232),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_245),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_221),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_247),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_414),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_222),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_409),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_335),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_104),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_435),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_242),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_30),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_361),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_622),
.Y(n_975)
);

INVxp33_ASAP7_75t_L g976 ( 
.A(n_861),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_697),
.Y(n_977)
);

CKINVDCx16_ASAP7_75t_R g978 ( 
.A(n_747),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_600),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_550),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_550),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_666),
.B(n_0),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_550),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_697),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_848),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_848),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_697),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_697),
.Y(n_988)
);

CKINVDCx16_ASAP7_75t_R g989 ( 
.A(n_847),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_848),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_697),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_561),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_872),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_561),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_620),
.Y(n_995)
);

CKINVDCx16_ASAP7_75t_R g996 ( 
.A(n_932),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_609),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_817),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_620),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_705),
.Y(n_1000)
);

INVxp67_ASAP7_75t_SL g1001 ( 
.A(n_705),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_820),
.Y(n_1002)
);

INVxp33_ASAP7_75t_SL g1003 ( 
.A(n_862),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_697),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_820),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_956),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_956),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_959),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_609),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_817),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_697),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_692),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_959),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_857),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_600),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_692),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_857),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_551),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_758),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_562),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_551),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_556),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_586),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_556),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_558),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_655),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_558),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_655),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_758),
.Y(n_1029)
);

INVxp33_ASAP7_75t_L g1030 ( 
.A(n_581),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_581),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_686),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_601),
.Y(n_1033)
);

INVxp33_ASAP7_75t_L g1034 ( 
.A(n_601),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_602),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_593),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_602),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_553),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_553),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_560),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_560),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_598),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_686),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_598),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_904),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_555),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_605),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_586),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_586),
.Y(n_1049)
);

CKINVDCx16_ASAP7_75t_R g1050 ( 
.A(n_740),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_605),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_586),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_614),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_904),
.Y(n_1054)
);

INVxp67_ASAP7_75t_SL g1055 ( 
.A(n_586),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_762),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_614),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_790),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_628),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_628),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_647),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_790),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_790),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_647),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_577),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_661),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_661),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_694),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_790),
.Y(n_1069)
);

INVxp33_ASAP7_75t_SL g1070 ( 
.A(n_795),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_740),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_694),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_753),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_577),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_702),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_562),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_753),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_702),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_593),
.Y(n_1079)
);

INVxp67_ASAP7_75t_SL g1080 ( 
.A(n_790),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_763),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_724),
.Y(n_1082)
);

BUFx2_ASAP7_75t_SL g1083 ( 
.A(n_577),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_724),
.B(n_2),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_965),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_944),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_743),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_743),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_750),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_733),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_944),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_750),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_764),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_606),
.Y(n_1094)
);

BUFx8_ASAP7_75t_SL g1095 ( 
.A(n_589),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_603),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_965),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_603),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_969),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_965),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_969),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_615),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_615),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_590),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_617),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_617),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_624),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_606),
.Y(n_1108)
);

INVxp33_ASAP7_75t_SL g1109 ( 
.A(n_552),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_606),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_624),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_625),
.Y(n_1112)
);

INVxp33_ASAP7_75t_SL g1113 ( 
.A(n_554),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_965),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_763),
.Y(n_1115)
);

CKINVDCx14_ASAP7_75t_R g1116 ( 
.A(n_576),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_616),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_965),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_864),
.Y(n_1119)
);

INVxp33_ASAP7_75t_SL g1120 ( 
.A(n_563),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_764),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_625),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_627),
.Y(n_1123)
);

INVxp67_ASAP7_75t_SL g1124 ( 
.A(n_627),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_864),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_630),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_630),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_840),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_864),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_770),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_881),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_607),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_634),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_770),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_634),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_733),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_813),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_645),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_813),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_645),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_650),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_650),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_665),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_881),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_771),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_665),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_865),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_672),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_672),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_662),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_771),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_674),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_674),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_678),
.Y(n_1154)
);

INVxp33_ASAP7_75t_SL g1155 ( 
.A(n_567),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_675),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_678),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_681),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_681),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_682),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_682),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_616),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_635),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_688),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_688),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_689),
.Y(n_1166)
);

INVxp33_ASAP7_75t_L g1167 ( 
.A(n_689),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_706),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_800),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_706),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_840),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_709),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_709),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_717),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_R g1175 ( 
.A(n_569),
.B(n_340),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_717),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_570),
.Y(n_1177)
);

INVxp33_ASAP7_75t_L g1178 ( 
.A(n_719),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_881),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_968),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_800),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_719),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_736),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_812),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_736),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_772),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_772),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_778),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_778),
.Y(n_1189)
);

CKINVDCx16_ASAP7_75t_R g1190 ( 
.A(n_715),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_779),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_779),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_781),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_573),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_781),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_786),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_786),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_578),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_815),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_720),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_815),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_822),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_822),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_826),
.Y(n_1204)
);

INVxp33_ASAP7_75t_L g1205 ( 
.A(n_826),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_834),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_635),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_834),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_760),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_865),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_837),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_837),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_846),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_846),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_571),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_850),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_580),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_850),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_812),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_860),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_860),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_824),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_871),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_579),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_871),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_591),
.Y(n_1226)
);

CKINVDCx16_ASAP7_75t_R g1227 ( 
.A(n_715),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_873),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_873),
.Y(n_1229)
);

INVxp33_ASAP7_75t_L g1230 ( 
.A(n_880),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_880),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_571),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_619),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_883),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_824),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_843),
.Y(n_1236)
);

INVxp33_ASAP7_75t_SL g1237 ( 
.A(n_583),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_843),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_715),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_640),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_767),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_867),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_867),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_878),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_878),
.Y(n_1245)
);

INVxp33_ASAP7_75t_L g1246 ( 
.A(n_883),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_892),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_768),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_885),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_885),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_891),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_892),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_691),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_759),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_891),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_797),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_898),
.Y(n_1257)
);

INVxp33_ASAP7_75t_L g1258 ( 
.A(n_898),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_906),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_906),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_895),
.Y(n_1261)
);

INVxp33_ASAP7_75t_SL g1262 ( 
.A(n_584),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_895),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_L g1264 ( 
.A(n_798),
.B(n_2),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_913),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_913),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_918),
.Y(n_1267)
);

CKINVDCx16_ASAP7_75t_R g1268 ( 
.A(n_715),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_920),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_920),
.Y(n_1270)
);

INVxp33_ASAP7_75t_SL g1271 ( 
.A(n_587),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_929),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_929),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_930),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_853),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_930),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_943),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_943),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_918),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_940),
.Y(n_1280)
);

INVxp33_ASAP7_75t_SL g1281 ( 
.A(n_597),
.Y(n_1281)
);

INVxp33_ASAP7_75t_SL g1282 ( 
.A(n_599),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_940),
.B(n_3),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_948),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_794),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_948),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_798),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_952),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_952),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_960),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_960),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_585),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_588),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_588),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_592),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_585),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_592),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_684),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_806),
.Y(n_1299)
);

CKINVDCx14_ASAP7_75t_R g1300 ( 
.A(n_921),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_684),
.Y(n_1301)
);

INVxp33_ASAP7_75t_L g1302 ( 
.A(n_828),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_971),
.Y(n_1303)
);

INVxp33_ASAP7_75t_SL g1304 ( 
.A(n_604),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_801),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_807),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_828),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_841),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_629),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_801),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_611),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_841),
.Y(n_1312)
);

INVxp33_ASAP7_75t_SL g1313 ( 
.A(n_623),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_631),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_844),
.B(n_4),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_844),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_886),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_827),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_886),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_889),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_922),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_629),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_643),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_889),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_939),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_939),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_632),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_643),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_633),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_685),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_637),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_829),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_922),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_803),
.B(n_4),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_934),
.B(n_6),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_866),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_738),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_622),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_595),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_638),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_970),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_639),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_738),
.Y(n_1343)
);

INVxp33_ASAP7_75t_SL g1344 ( 
.A(n_646),
.Y(n_1344)
);

INVxp33_ASAP7_75t_L g1345 ( 
.A(n_685),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1070),
.B(n_819),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_975),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1302),
.B(n_738),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_975),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_975),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1065),
.B(n_773),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_975),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1020),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1020),
.B(n_618),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1023),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1076),
.B(n_618),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_975),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1345),
.B(n_995),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1338),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1338),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1180),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1049),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_978),
.B(n_738),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1065),
.B(n_773),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1076),
.Y(n_1365)
);

BUFx8_ASAP7_75t_L g1366 ( 
.A(n_1099),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1338),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1070),
.B(n_557),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1049),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1090),
.Y(n_1370)
);

AND2x6_ASAP7_75t_L g1371 ( 
.A(n_1038),
.B(n_899),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1056),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_L g1373 ( 
.A(n_1330),
.B(n_564),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1338),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1052),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1052),
.Y(n_1376)
);

BUFx8_ASAP7_75t_SL g1377 ( 
.A(n_1095),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1090),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1028),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_989),
.B(n_776),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1136),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1337),
.B(n_613),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1338),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1001),
.B(n_663),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1330),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1343),
.B(n_663),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1007),
.B(n_793),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_996),
.B(n_776),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1058),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1056),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1050),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1121),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1058),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1261),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1048),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1121),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1062),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1136),
.B(n_1137),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1261),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1062),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1073),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1118),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1134),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1137),
.B(n_793),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1036),
.B(n_899),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1086),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_984),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1118),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1267),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1180),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1139),
.B(n_1147),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_984),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1267),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1134),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1139),
.B(n_572),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1145),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1147),
.B(n_612),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1300),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_988),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_993),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1055),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_988),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_991),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_993),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_991),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1043),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1079),
.B(n_695),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1004),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1004),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1145),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1011),
.Y(n_1431)
);

INVx5_ASAP7_75t_L g1432 ( 
.A(n_1011),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1210),
.B(n_701),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1081),
.B(n_780),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_977),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1210),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1074),
.B(n_1094),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1083),
.B(n_776),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1091),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1151),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_977),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_987),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1292),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_987),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1292),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1038),
.B(n_559),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1116),
.B(n_565),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1074),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1063),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_979),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1083),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_980),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1179),
.B(n_566),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1069),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1179),
.B(n_568),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1039),
.B(n_659),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1296),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1101),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1094),
.B(n_574),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1108),
.B(n_575),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1296),
.Y(n_1461)
);

INVx5_ASAP7_75t_L g1462 ( 
.A(n_1309),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1039),
.B(n_677),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1309),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1080),
.B(n_582),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1099),
.B(n_776),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1085),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_SL g1468 ( 
.A(n_997),
.B(n_1009),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1151),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1169),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_997),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1097),
.B(n_594),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1009),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1100),
.B(n_596),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1114),
.B(n_608),
.Y(n_1475)
);

AND2x6_ASAP7_75t_L g1476 ( 
.A(n_1040),
.B(n_622),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1322),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1108),
.B(n_610),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1040),
.B(n_711),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1110),
.B(n_621),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1169),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_979),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1322),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1323),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1110),
.B(n_626),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1041),
.B(n_789),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1041),
.B(n_876),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1311),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1012),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1115),
.B(n_636),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1119),
.B(n_641),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_981),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1323),
.Y(n_1493)
);

BUFx8_ASAP7_75t_SL g1494 ( 
.A(n_1104),
.Y(n_1494)
);

CKINVDCx6p67_ASAP7_75t_R g1495 ( 
.A(n_1190),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1181),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_983),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1181),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_976),
.B(n_849),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1184),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1184),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1119),
.B(n_642),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_985),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1015),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1042),
.B(n_907),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1128),
.B(n_644),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1042),
.B(n_622),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_986),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1044),
.B(n_961),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1219),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1022),
.B(n_849),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1219),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1222),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1125),
.B(n_648),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1015),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_990),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1044),
.B(n_622),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_992),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1222),
.Y(n_1519)
);

BUFx8_ASAP7_75t_SL g1520 ( 
.A(n_1104),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1026),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1171),
.B(n_651),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_994),
.Y(n_1523)
);

INVx5_ASAP7_75t_L g1524 ( 
.A(n_1252),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1012),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1047),
.B(n_792),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1016),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1125),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1252),
.Y(n_1529)
);

INVx5_ASAP7_75t_L g1530 ( 
.A(n_1263),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1263),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1016),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1129),
.B(n_653),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1340),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1030),
.B(n_849),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1341),
.B(n_656),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_999),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1328),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1129),
.B(n_657),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1328),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1019),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1311),
.Y(n_1542)
);

BUFx8_ASAP7_75t_SL g1543 ( 
.A(n_1132),
.Y(n_1543)
);

INVx5_ASAP7_75t_L g1544 ( 
.A(n_1215),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1047),
.B(n_1051),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1215),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1215),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1051),
.B(n_792),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1284),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1053),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1131),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1284),
.Y(n_1552)
);

AND2x6_ASAP7_75t_L g1553 ( 
.A(n_1053),
.B(n_792),
.Y(n_1553)
);

INVx5_ASAP7_75t_L g1554 ( 
.A(n_1232),
.Y(n_1554)
);

INVx6_ASAP7_75t_L g1555 ( 
.A(n_1227),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1117),
.B(n_658),
.Y(n_1556)
);

INVx5_ASAP7_75t_L g1557 ( 
.A(n_1232),
.Y(n_1557)
);

INVx5_ASAP7_75t_L g1558 ( 
.A(n_1232),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1301),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1117),
.B(n_669),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1026),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1131),
.B(n_670),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1057),
.Y(n_1563)
);

INVx5_ASAP7_75t_L g1564 ( 
.A(n_1301),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1057),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1059),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1059),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1060),
.B(n_792),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1034),
.B(n_849),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1301),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1144),
.B(n_671),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1303),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1060),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1162),
.B(n_673),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1061),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1061),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1167),
.B(n_912),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1064),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1178),
.B(n_912),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1064),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1066),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1019),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1032),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1066),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1144),
.B(n_679),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1032),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1067),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1067),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1000),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1068),
.B(n_1072),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1068),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1072),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1075),
.B(n_792),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1075),
.Y(n_1594)
);

INVx5_ASAP7_75t_L g1595 ( 
.A(n_1162),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1124),
.B(n_683),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1078),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1126),
.B(n_698),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1078),
.B(n_927),
.Y(n_1599)
);

INVx5_ASAP7_75t_L g1600 ( 
.A(n_1163),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1082),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1127),
.B(n_708),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1071),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1177),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1082),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1087),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1217),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1029),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1002),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1087),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1088),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1314),
.Y(n_1612)
);

BUFx12f_ASAP7_75t_L g1613 ( 
.A(n_1029),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1045),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1088),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1149),
.B(n_1159),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1205),
.B(n_912),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1166),
.B(n_718),
.Y(n_1618)
);

AND2x6_ASAP7_75t_L g1619 ( 
.A(n_1089),
.B(n_927),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1089),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1183),
.B(n_1188),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1092),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1092),
.Y(n_1623)
);

BUFx12f_ASAP7_75t_L g1624 ( 
.A(n_1045),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1093),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1230),
.B(n_912),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1195),
.B(n_722),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1093),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1202),
.B(n_723),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1246),
.B(n_595),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1258),
.B(n_595),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1130),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1130),
.Y(n_1633)
);

INVx6_ASAP7_75t_L g1634 ( 
.A(n_1239),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1203),
.B(n_725),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1340),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1270),
.B(n_728),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1235),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1005),
.B(n_729),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1071),
.Y(n_1640)
);

INVxp33_ASAP7_75t_SL g1641 ( 
.A(n_1054),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1235),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1236),
.B(n_927),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1006),
.B(n_734),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1236),
.B(n_1238),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1319),
.B(n_649),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1008),
.B(n_735),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1013),
.B(n_739),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1238),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1242),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1243),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1163),
.B(n_652),
.Y(n_1653)
);

BUFx8_ASAP7_75t_L g1654 ( 
.A(n_1207),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1244),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1207),
.B(n_748),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1244),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1441),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1427),
.B(n_1054),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1427),
.B(n_1245),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1452),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1452),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1412),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1412),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1422),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1422),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1379),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1549),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1545),
.B(n_1268),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1348),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1423),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1423),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1549),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1549),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1549),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1391),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1434),
.B(n_1245),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1435),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1419),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1434),
.B(n_1247),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1552),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1385),
.B(n_1247),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1435),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1441),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1401),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1406),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1552),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1370),
.B(n_1192),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1385),
.B(n_1279),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1426),
.Y(n_1690)
);

AND2x6_ASAP7_75t_L g1691 ( 
.A(n_1438),
.B(n_1279),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1419),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1442),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1442),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1385),
.B(n_1358),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1419),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1552),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1441),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1441),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1370),
.B(n_1280),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1353),
.B(n_1264),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1353),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1444),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1419),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1365),
.B(n_1287),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1444),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1439),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1394),
.B(n_1280),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1552),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1565),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1565),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1425),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1565),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1458),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1545),
.B(n_1287),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1425),
.Y(n_1716)
);

AND2x6_ASAP7_75t_L g1717 ( 
.A(n_1446),
.B(n_927),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1545),
.B(n_1305),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1444),
.Y(n_1719)
);

CKINVDCx16_ASAP7_75t_R g1720 ( 
.A(n_1420),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1565),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1365),
.B(n_1305),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1566),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1566),
.Y(n_1724)
);

AND2x6_ASAP7_75t_L g1725 ( 
.A(n_1446),
.B(n_927),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1566),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1378),
.B(n_1315),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1566),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1446),
.B(n_1046),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1444),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1425),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1555),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1630),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1425),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1576),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1378),
.B(n_1315),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1428),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1352),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1381),
.B(n_1018),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1428),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1428),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1428),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1352),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1429),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1429),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1534),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1576),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1381),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1590),
.B(n_1021),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1436),
.B(n_1024),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1429),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1436),
.B(n_1025),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1590),
.B(n_1027),
.Y(n_1753)
);

AND3x2_ASAP7_75t_L g1754 ( 
.A(n_1372),
.B(n_1339),
.C(n_1014),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1576),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1411),
.B(n_1031),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1576),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1590),
.B(n_1033),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1580),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1429),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1431),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1394),
.B(n_1314),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1636),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1394),
.B(n_1327),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1399),
.B(n_1327),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1580),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1368),
.A2(n_982),
.B1(n_1003),
.B2(n_1109),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1431),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1431),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1580),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1580),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1431),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1377),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1362),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1631),
.Y(n_1775)
);

AND2x6_ASAP7_75t_L g1776 ( 
.A(n_1456),
.B(n_936),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1420),
.B(n_1217),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1399),
.B(n_1329),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1511),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1352),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1645),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1362),
.Y(n_1782)
);

BUFx8_ASAP7_75t_L g1783 ( 
.A(n_1361),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1369),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1587),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1587),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1587),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1595),
.B(n_1109),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1369),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1399),
.B(n_1329),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1587),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1375),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1594),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1594),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1375),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1409),
.B(n_1331),
.Y(n_1796)
);

CKINVDCx11_ASAP7_75t_R g1797 ( 
.A(n_1361),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1409),
.B(n_1331),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1376),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1500),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1376),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1393),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1594),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1594),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1409),
.B(n_1413),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1597),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1500),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1500),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1411),
.B(n_1035),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1500),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1413),
.B(n_1344),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1597),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1393),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1346),
.A2(n_1132),
.B1(n_1156),
.B2(n_1150),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1645),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1645),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1456),
.B(n_1463),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1535),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1397),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1597),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1411),
.B(n_1037),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1597),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1510),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1413),
.B(n_1344),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1606),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1456),
.B(n_1096),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1510),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1463),
.B(n_1098),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1510),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1377),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1606),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1606),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1606),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1595),
.B(n_1600),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1451),
.B(n_1113),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1611),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1397),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1463),
.B(n_1102),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1651),
.A2(n_1084),
.B(n_1283),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1479),
.B(n_1103),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1595),
.B(n_1113),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1479),
.B(n_1105),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1479),
.B(n_1106),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1611),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1510),
.Y(n_1845)
);

INVx6_ASAP7_75t_L g1846 ( 
.A(n_1546),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1611),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1513),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1486),
.B(n_1107),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1611),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1645),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1620),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1620),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1408),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1417),
.B(n_1120),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1408),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1620),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1464),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1494),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1487),
.B(n_1111),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1620),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1638),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1464),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1483),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1368),
.A2(n_1003),
.B1(n_1155),
.B2(n_1120),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1505),
.B(n_1112),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1595),
.B(n_1155),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1638),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1513),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1595),
.B(n_1237),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1483),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1550),
.A2(n_1123),
.B(n_1122),
.Y(n_1874)
);

BUFx10_ASAP7_75t_L g1875 ( 
.A(n_1346),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1493),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1513),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1550),
.A2(n_1135),
.B(n_1133),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1638),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1351),
.A2(n_1237),
.B1(n_1271),
.B2(n_1262),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1493),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1638),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1417),
.B(n_1262),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1645),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1505),
.B(n_1138),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1645),
.Y(n_1886)
);

AND2x2_ASAP7_75t_SL g1887 ( 
.A(n_1505),
.B(n_1334),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1513),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1496),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1496),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1642),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1642),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1642),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1519),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1529),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1642),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1519),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1417),
.B(n_1271),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1649),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1494),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1649),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1445),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1600),
.B(n_1281),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1509),
.B(n_1140),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1649),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1649),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1655),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1509),
.B(n_1141),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1445),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1655),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1445),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1445),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1655),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1457),
.Y(n_1914)
);

CKINVDCx8_ASAP7_75t_R g1915 ( 
.A(n_1418),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1655),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1657),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1657),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1457),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1433),
.B(n_1313),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1509),
.B(n_1142),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1657),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1569),
.B(n_1143),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1457),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1476),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1577),
.Y(n_1926)
);

BUFx12f_ASAP7_75t_L g1927 ( 
.A(n_1366),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1657),
.Y(n_1928)
);

OR2x6_ASAP7_75t_L g1929 ( 
.A(n_1410),
.B(n_1471),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1563),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1579),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1575),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1584),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1457),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1453),
.B(n_1281),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1461),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1461),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1588),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1529),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1591),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1601),
.Y(n_1941)
);

AND2x6_ASAP7_75t_L g1942 ( 
.A(n_1363),
.B(n_936),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1625),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1433),
.B(n_1282),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1567),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1455),
.B(n_1282),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1567),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1573),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1461),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1573),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1617),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1433),
.B(n_1304),
.Y(n_1952)
);

CKINVDCx20_ASAP7_75t_R g1953 ( 
.A(n_1520),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1600),
.B(n_1304),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1578),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1578),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1461),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1477),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1581),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1581),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1626),
.B(n_1146),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1592),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1592),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1578),
.Y(n_1964)
);

OA21x2_ASAP7_75t_L g1965 ( 
.A1(n_1605),
.A2(n_1152),
.B(n_1148),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1373),
.B(n_1153),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1450),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1605),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1477),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1546),
.B(n_1313),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1622),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1610),
.Y(n_1972)
);

INVx4_ASAP7_75t_L g1973 ( 
.A(n_1622),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1610),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1482),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1654),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1615),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1615),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1354),
.B(n_1356),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1628),
.A2(n_1157),
.B(n_1154),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1628),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1633),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1654),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1622),
.B(n_1158),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1477),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1623),
.B(n_1160),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1477),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1633),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1529),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1546),
.B(n_1194),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_L g1991 ( 
.A(n_1448),
.B(n_1175),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1650),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1650),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1484),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1484),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1559),
.B(n_1570),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1652),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1484),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1484),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1663),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1817),
.B(n_1646),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1663),
.Y(n_2002)
);

OR2x6_ASAP7_75t_L g2003 ( 
.A(n_1929),
.B(n_1410),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1678),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1664),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1660),
.B(n_1536),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1664),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1973),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1665),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1665),
.Y(n_2010)
);

INVxp67_ASAP7_75t_SL g2011 ( 
.A(n_1781),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1874),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1874),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1773),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1666),
.Y(n_2015)
);

INVx4_ASAP7_75t_L g2016 ( 
.A(n_1886),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1659),
.B(n_1641),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1677),
.B(n_1536),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1781),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1874),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1817),
.B(n_1646),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1973),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1678),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1666),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1973),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1887),
.B(n_1448),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1887),
.B(n_1528),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1671),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1683),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1671),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1680),
.B(n_1528),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1773),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1830),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1683),
.Y(n_2034)
);

BUFx10_ASAP7_75t_L g2035 ( 
.A(n_1835),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1855),
.B(n_1551),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1693),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1672),
.Y(n_2038)
);

CKINVDCx20_ASAP7_75t_R g2039 ( 
.A(n_1814),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1672),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1693),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1694),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1781),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1691),
.B(n_1551),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1883),
.B(n_1468),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1898),
.B(n_1600),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1694),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1858),
.A2(n_1351),
.B1(n_1364),
.B2(n_1499),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1846),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1889),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1830),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1920),
.B(n_1600),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1815),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1944),
.B(n_1952),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1859),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1859),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1865),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1865),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_1815),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1866),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1889),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1691),
.B(n_1556),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1858),
.B(n_1518),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1890),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1866),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1873),
.Y(n_2066)
);

INVxp33_ASAP7_75t_L g2067 ( 
.A(n_1690),
.Y(n_2067)
);

OAI22xp33_ASAP7_75t_SL g2068 ( 
.A1(n_1767),
.A2(n_1364),
.B1(n_1233),
.B2(n_1240),
.Y(n_2068)
);

INVx4_ASAP7_75t_L g2069 ( 
.A(n_1886),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_1815),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1688),
.B(n_1604),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1873),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1876),
.Y(n_2073)
);

INVx3_ASAP7_75t_L g2074 ( 
.A(n_1816),
.Y(n_2074)
);

INVx4_ASAP7_75t_L g2075 ( 
.A(n_1886),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_1816),
.Y(n_2076)
);

OAI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_1867),
.A2(n_1334),
.B1(n_1335),
.B2(n_1604),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1746),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1691),
.B(n_1556),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1876),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1890),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1894),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1816),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_L g2084 ( 
.A(n_1691),
.B(n_1851),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1894),
.Y(n_2085)
);

NAND2xp33_ASAP7_75t_L g2086 ( 
.A(n_1691),
.B(n_1851),
.Y(n_2086)
);

INVxp67_ASAP7_75t_SL g2087 ( 
.A(n_1851),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_L g2088 ( 
.A(n_1691),
.B(n_1488),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1667),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1688),
.B(n_1641),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1881),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1881),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1695),
.B(n_1560),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1878),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1884),
.Y(n_2095)
);

BUFx10_ASAP7_75t_L g2096 ( 
.A(n_1935),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1688),
.B(n_1542),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1860),
.B(n_1623),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1946),
.A2(n_1632),
.B1(n_1382),
.B2(n_1623),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1878),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_L g2101 ( 
.A(n_1884),
.B(n_1612),
.Y(n_2101)
);

NAND3xp33_ASAP7_75t_L g2102 ( 
.A(n_1991),
.B(n_1574),
.C(n_1560),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1679),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1878),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1774),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1774),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1965),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1782),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1875),
.B(n_1437),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1965),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1984),
.B(n_1574),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1782),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1897),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1784),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1880),
.B(n_1437),
.Y(n_2115)
);

NAND2xp33_ASAP7_75t_SL g2116 ( 
.A(n_1970),
.B(n_1478),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1860),
.B(n_1466),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1875),
.B(n_1555),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1984),
.B(n_1656),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1875),
.B(n_1555),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1702),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1986),
.B(n_1656),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1784),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1986),
.B(n_1490),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1923),
.B(n_1490),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_1667),
.Y(n_2126)
);

OAI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1779),
.A2(n_1818),
.B1(n_1931),
.B2(n_1926),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_1884),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1789),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1797),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1923),
.B(n_1506),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1897),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1789),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1961),
.B(n_1506),
.Y(n_2134)
);

INVxp67_ASAP7_75t_SL g2135 ( 
.A(n_1679),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_1953),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1961),
.B(n_1522),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1792),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1792),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1965),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1795),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1795),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_1846),
.Y(n_2143)
);

INVxp67_ASAP7_75t_SL g2144 ( 
.A(n_1679),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1702),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1980),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1799),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1980),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1669),
.B(n_1979),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1980),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1846),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1955),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_SL g2153 ( 
.A(n_1929),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1955),
.B(n_1522),
.Y(n_2154)
);

AND3x1_ASAP7_75t_L g2155 ( 
.A(n_1715),
.B(n_1382),
.C(n_1653),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1799),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1669),
.B(n_1480),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1955),
.B(n_1616),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1801),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1979),
.B(n_1485),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1956),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1801),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1802),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1802),
.Y(n_2164)
);

AND3x1_ASAP7_75t_L g2165 ( 
.A(n_1715),
.B(n_1502),
.C(n_1491),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1956),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1813),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1813),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1956),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1819),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1964),
.B(n_1621),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1819),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1837),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1837),
.Y(n_2174)
);

INVxp67_ASAP7_75t_SL g2175 ( 
.A(n_1679),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1854),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_1846),
.Y(n_2177)
);

AOI21x1_ASAP7_75t_L g2178 ( 
.A1(n_1854),
.A2(n_1526),
.B(n_1517),
.Y(n_2178)
);

NAND2xp33_ASAP7_75t_SL g2179 ( 
.A(n_1788),
.B(n_1514),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1856),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1670),
.B(n_1634),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1746),
.B(n_1634),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1856),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1964),
.B(n_1632),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1979),
.B(n_1533),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1964),
.Y(n_2186)
);

INVx2_ASAP7_75t_SL g2187 ( 
.A(n_1729),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1971),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1971),
.B(n_1632),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1971),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1945),
.Y(n_2191)
);

NAND3xp33_ASAP7_75t_L g2192 ( 
.A(n_1991),
.B(n_1460),
.C(n_1459),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1947),
.Y(n_2193)
);

NOR2x1p5_ASAP7_75t_L g2194 ( 
.A(n_1861),
.B(n_1495),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1700),
.B(n_1717),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1948),
.Y(n_2196)
);

OR2x6_ASAP7_75t_L g2197 ( 
.A(n_1929),
.B(n_1471),
.Y(n_2197)
);

INVxp67_ASAP7_75t_L g2198 ( 
.A(n_1763),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1811),
.B(n_1539),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_1763),
.B(n_1634),
.Y(n_2200)
);

AND2x6_ASAP7_75t_L g2201 ( 
.A(n_1826),
.B(n_1380),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1950),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1824),
.B(n_1562),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_1676),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1959),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_1658),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1717),
.B(n_1405),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1679),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_1692),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1960),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_1676),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1962),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_1996),
.B(n_1571),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1963),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1930),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1932),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1717),
.B(n_1405),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_1729),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1968),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1972),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1974),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1717),
.B(n_1596),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1826),
.B(n_1585),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_1800),
.Y(n_2224)
);

NAND3xp33_ASAP7_75t_L g2225 ( 
.A(n_1733),
.B(n_1460),
.C(n_1459),
.Y(n_2225)
);

BUFx3_ASAP7_75t_L g2226 ( 
.A(n_1748),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1717),
.B(n_1725),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1977),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1717),
.B(n_1598),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1658),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1978),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1981),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1826),
.B(n_1602),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1982),
.Y(n_2234)
);

NAND2xp33_ASAP7_75t_L g2235 ( 
.A(n_1762),
.B(n_902),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1842),
.B(n_1388),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1988),
.Y(n_2237)
);

INVxp33_ASAP7_75t_L g2238 ( 
.A(n_1707),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_1658),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1992),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1842),
.B(n_1843),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1993),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1842),
.B(n_1618),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_1686),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_1843),
.B(n_1627),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1705),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1933),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1997),
.Y(n_2248)
);

INVx5_ASAP7_75t_L g2249 ( 
.A(n_1692),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1748),
.Y(n_2250)
);

OAI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_1951),
.A2(n_1775),
.B1(n_1335),
.B2(n_1990),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1699),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1699),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_1843),
.B(n_1629),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_1868),
.B(n_1908),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1938),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_1686),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1940),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1725),
.B(n_1635),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1721),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1721),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1868),
.B(n_1200),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1725),
.B(n_1637),
.Y(n_2263)
);

CKINVDCx8_ASAP7_75t_R g2264 ( 
.A(n_1720),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1868),
.B(n_1424),
.Y(n_2265)
);

BUFx3_ASAP7_75t_L g2266 ( 
.A(n_1732),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1725),
.B(n_1386),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1728),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1703),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1703),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1908),
.B(n_1424),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_1684),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1706),
.Y(n_2273)
);

OAI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_1777),
.A2(n_1607),
.B1(n_1489),
.B2(n_1525),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1706),
.Y(n_2275)
);

INVxp67_ASAP7_75t_SL g2276 ( 
.A(n_1692),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1728),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1719),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1908),
.B(n_1473),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1755),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1705),
.B(n_1473),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1719),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1828),
.B(n_1332),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1730),
.Y(n_2284)
);

AND2x6_ASAP7_75t_L g2285 ( 
.A(n_1828),
.B(n_1517),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1725),
.B(n_1386),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1725),
.B(n_1776),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1730),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1755),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_1684),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1757),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_1967),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1757),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1759),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1731),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1838),
.B(n_1241),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1731),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1759),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1941),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1705),
.B(n_1489),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1737),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1943),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_1722),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_1722),
.B(n_1525),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_1975),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1737),
.Y(n_2306)
);

NOR2x1p5_ASAP7_75t_L g2307 ( 
.A(n_1861),
.B(n_1495),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_1684),
.Y(n_2308)
);

NAND3xp33_ASAP7_75t_L g2309 ( 
.A(n_1718),
.B(n_1224),
.C(n_1198),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1740),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_1698),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1776),
.B(n_1559),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1776),
.B(n_1559),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1668),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1673),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1764),
.B(n_1765),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_1714),
.B(n_1299),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_1722),
.B(n_1527),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_1776),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1740),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_1778),
.B(n_1226),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1674),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1675),
.Y(n_2323)
);

INVx4_ASAP7_75t_L g2324 ( 
.A(n_1800),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1741),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1741),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1681),
.Y(n_2327)
);

AO21x2_ASAP7_75t_L g2328 ( 
.A1(n_1687),
.A2(n_1404),
.B(n_1639),
.Y(n_2328)
);

NAND3xp33_ASAP7_75t_L g2329 ( 
.A(n_1718),
.B(n_1342),
.C(n_1607),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_1692),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_1698),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1756),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1756),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_1838),
.B(n_1336),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_1692),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_1696),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1790),
.B(n_1796),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1697),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1709),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1710),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_1798),
.B(n_1226),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1696),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1701),
.B(n_1527),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_SL g2344 ( 
.A1(n_1953),
.A2(n_1150),
.B1(n_1209),
.B2(n_1156),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_1788),
.A2(n_1354),
.B1(n_1356),
.B2(n_1465),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_L g2346 ( 
.A(n_1841),
.B(n_1233),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_1841),
.B(n_1240),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2006),
.B(n_1839),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2299),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_2103),
.Y(n_2350)
);

XOR2xp5_ASAP7_75t_L g2351 ( 
.A(n_2014),
.B(n_1900),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2299),
.Y(n_2352)
);

INVxp67_ASAP7_75t_SL g2353 ( 
.A(n_2084),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2266),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2283),
.B(n_1840),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2017),
.B(n_1869),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2018),
.B(n_1839),
.Y(n_2357)
);

NOR2xp67_ASAP7_75t_L g2358 ( 
.A(n_2182),
.B(n_1927),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2302),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2302),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2246),
.B(n_2303),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2246),
.B(n_1749),
.Y(n_2362)
);

XOR2xp5_ASAP7_75t_L g2363 ( 
.A(n_2014),
.B(n_1900),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2215),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2216),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2283),
.B(n_1840),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2126),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2000),
.Y(n_2368)
);

XOR2xp5_ASAP7_75t_L g2369 ( 
.A(n_2032),
.B(n_1209),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2247),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2256),
.Y(n_2371)
);

CKINVDCx20_ASAP7_75t_R g2372 ( 
.A(n_2136),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2258),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2296),
.B(n_2334),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2098),
.Y(n_2375)
);

CKINVDCx20_ASAP7_75t_R g2376 ( 
.A(n_2136),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2098),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2296),
.B(n_1849),
.Y(n_2378)
);

INVxp67_ASAP7_75t_SL g2379 ( 
.A(n_2084),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2303),
.B(n_1749),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2260),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2260),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2334),
.B(n_1849),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2031),
.B(n_1869),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2261),
.Y(n_2385)
);

INVxp33_ASAP7_75t_L g2386 ( 
.A(n_2317),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2261),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2262),
.B(n_1862),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2268),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2262),
.B(n_1862),
.Y(n_2390)
);

BUFx3_ASAP7_75t_L g2391 ( 
.A(n_2266),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2268),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2000),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2204),
.B(n_1504),
.Y(n_2394)
);

HB1xp67_ASAP7_75t_L g2395 ( 
.A(n_2089),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2089),
.B(n_2257),
.Y(n_2396)
);

XNOR2x1_ASAP7_75t_L g2397 ( 
.A(n_2077),
.B(n_1253),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2277),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2002),
.Y(n_2399)
);

AND2x6_ASAP7_75t_L g2400 ( 
.A(n_2043),
.B(n_1753),
.Y(n_2400)
);

CKINVDCx20_ASAP7_75t_R g2401 ( 
.A(n_2032),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2277),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2280),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2280),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2289),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2109),
.B(n_1915),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2289),
.Y(n_2407)
);

NAND2x1p5_ASAP7_75t_L g2408 ( 
.A(n_2143),
.B(n_1896),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2291),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2291),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2293),
.Y(n_2411)
);

XOR2x2_ASAP7_75t_L g2412 ( 
.A(n_2344),
.B(n_1754),
.Y(n_2412)
);

INVxp67_ASAP7_75t_SL g2413 ( 
.A(n_2086),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2293),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2294),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2294),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2298),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2298),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2193),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2193),
.Y(n_2420)
);

XOR2xp5_ASAP7_75t_L g2421 ( 
.A(n_2033),
.B(n_1248),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2124),
.B(n_2111),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2205),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2205),
.Y(n_2424)
);

NAND2xp33_ASAP7_75t_R g2425 ( 
.A(n_2033),
.B(n_1572),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2210),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2002),
.Y(n_2427)
);

XNOR2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2130),
.B(n_1976),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2210),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2257),
.B(n_1885),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2214),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2214),
.Y(n_2432)
);

INVxp67_ASAP7_75t_L g2433 ( 
.A(n_2211),
.Y(n_2433)
);

AND2x6_ASAP7_75t_L g2434 ( 
.A(n_2043),
.B(n_1753),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2292),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2219),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2219),
.Y(n_2437)
);

INVxp67_ASAP7_75t_SL g2438 ( 
.A(n_2086),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_2115),
.B(n_1872),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2149),
.B(n_1872),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2232),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2232),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2119),
.B(n_1839),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2122),
.B(n_1758),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2234),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2005),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2234),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_SL g2448 ( 
.A(n_2003),
.Y(n_2448)
);

CKINVDCx20_ASAP7_75t_R g2449 ( 
.A(n_2051),
.Y(n_2449)
);

INVx2_ASAP7_75t_SL g2450 ( 
.A(n_2317),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2237),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2005),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2007),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2237),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2242),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2187),
.B(n_1885),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2151),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2242),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2161),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2161),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2007),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2054),
.B(n_1903),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2166),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2166),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2169),
.Y(n_2465)
);

XOR2xp5_ASAP7_75t_L g2466 ( 
.A(n_2051),
.B(n_1248),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2169),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2009),
.Y(n_2468)
);

BUFx6f_ASAP7_75t_SL g2469 ( 
.A(n_2003),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2191),
.Y(n_2470)
);

AND2x2_ASAP7_75t_SL g2471 ( 
.A(n_2088),
.B(n_1976),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2009),
.Y(n_2472)
);

XNOR2x2_ASAP7_75t_L g2473 ( 
.A(n_2346),
.B(n_1904),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2191),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2196),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2196),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_SL g2477 ( 
.A(n_2264),
.B(n_1927),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2187),
.B(n_1904),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2130),
.Y(n_2479)
);

XNOR2xp5_ASAP7_75t_L g2480 ( 
.A(n_2274),
.B(n_1285),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_2264),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2093),
.B(n_1903),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2218),
.B(n_1921),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_2292),
.Y(n_2484)
);

NAND2xp33_ASAP7_75t_R g2485 ( 
.A(n_2197),
.B(n_1418),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2202),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2202),
.Y(n_2487)
);

CKINVDCx20_ASAP7_75t_R g2488 ( 
.A(n_2305),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2212),
.Y(n_2489)
);

XNOR2xp5_ASAP7_75t_L g2490 ( 
.A(n_2039),
.B(n_1285),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2212),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2125),
.B(n_1758),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2220),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2103),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2220),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2221),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2221),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2062),
.A2(n_1689),
.B(n_1682),
.Y(n_2498)
);

INVx1_ASAP7_75t_SL g2499 ( 
.A(n_2305),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2103),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2228),
.Y(n_2501)
);

XOR2xp5_ASAP7_75t_L g2502 ( 
.A(n_2039),
.B(n_1306),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2010),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2228),
.Y(n_2504)
);

AND2x6_ASAP7_75t_L g2505 ( 
.A(n_2043),
.B(n_1921),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2231),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2026),
.B(n_1954),
.Y(n_2507)
);

XOR2x2_ASAP7_75t_L g2508 ( 
.A(n_2068),
.B(n_1521),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2231),
.Y(n_2509)
);

CKINVDCx20_ASAP7_75t_R g2510 ( 
.A(n_2244),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2218),
.B(n_1253),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2240),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2240),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2248),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2027),
.B(n_1954),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2010),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2248),
.Y(n_2517)
);

CKINVDCx20_ASAP7_75t_R g2518 ( 
.A(n_2078),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2188),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2131),
.B(n_1661),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2188),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2004),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2001),
.B(n_1254),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2004),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2023),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2134),
.B(n_1662),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2015),
.Y(n_2527)
);

AND2x6_ASAP7_75t_L g2528 ( 
.A(n_2053),
.B(n_1966),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2023),
.Y(n_2529)
);

BUFx6f_ASAP7_75t_L g2530 ( 
.A(n_2103),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2015),
.Y(n_2531)
);

XOR2xp5_ASAP7_75t_L g2532 ( 
.A(n_2165),
.B(n_1306),
.Y(n_2532)
);

XOR2xp5_ASAP7_75t_L g2533 ( 
.A(n_2067),
.B(n_1318),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2137),
.B(n_1776),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2029),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2157),
.B(n_1727),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2029),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2034),
.Y(n_2538)
);

XOR2x2_ASAP7_75t_L g2539 ( 
.A(n_2155),
.B(n_1561),
.Y(n_2539)
);

INVxp67_ASAP7_75t_SL g2540 ( 
.A(n_2016),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2016),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2034),
.Y(n_2542)
);

CKINVDCx20_ASAP7_75t_R g2543 ( 
.A(n_2198),
.Y(n_2543)
);

XNOR2x2_ASAP7_75t_L g2544 ( 
.A(n_2347),
.B(n_1318),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2024),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2001),
.B(n_1254),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2037),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2021),
.B(n_1256),
.Y(n_2548)
);

AND2x6_ASAP7_75t_L g2549 ( 
.A(n_2053),
.B(n_1966),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2037),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2236),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2096),
.B(n_2090),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2332),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2333),
.Y(n_2554)
);

CKINVDCx16_ASAP7_75t_R g2555 ( 
.A(n_2003),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2200),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2153),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2024),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2050),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2021),
.B(n_1256),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2238),
.B(n_1583),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2028),
.Y(n_2562)
);

INVx3_ASAP7_75t_L g2563 ( 
.A(n_2151),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2158),
.B(n_1776),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2050),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2103),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2061),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2117),
.B(n_1275),
.Y(n_2568)
);

OAI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2079),
.A2(n_1708),
.B(n_1711),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2061),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2064),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2064),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2081),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2081),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2082),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2082),
.Y(n_2576)
);

NAND2x1p5_ASAP7_75t_L g2577 ( 
.A(n_2143),
.B(n_1896),
.Y(n_2577)
);

INVx2_ASAP7_75t_SL g2578 ( 
.A(n_2236),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2028),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2085),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2030),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2096),
.B(n_1727),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2085),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2113),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_L g2585 ( 
.A(n_2096),
.B(n_1727),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2113),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2132),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2132),
.Y(n_2588)
);

CKINVDCx20_ASAP7_75t_R g2589 ( 
.A(n_2003),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2097),
.B(n_1736),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2241),
.B(n_1756),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2199),
.B(n_1736),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2030),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2038),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2038),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2314),
.Y(n_2596)
);

CKINVDCx20_ASAP7_75t_R g2597 ( 
.A(n_2197),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2203),
.B(n_1736),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2117),
.B(n_1275),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2314),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2063),
.B(n_1983),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2315),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2315),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2322),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2063),
.B(n_1983),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2322),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_SL g2607 ( 
.A(n_2197),
.B(n_1915),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2323),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2323),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2143),
.B(n_1701),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2327),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2255),
.B(n_1809),
.Y(n_2612)
);

INVxp67_ASAP7_75t_SL g2613 ( 
.A(n_2016),
.Y(n_2613)
);

NAND2x1p5_ASAP7_75t_L g2614 ( 
.A(n_2143),
.B(n_1896),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2327),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2338),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2338),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2339),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2339),
.Y(n_2619)
);

CKINVDCx20_ASAP7_75t_R g2620 ( 
.A(n_2197),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2035),
.B(n_2223),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2340),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2340),
.Y(n_2623)
);

CKINVDCx20_ASAP7_75t_R g2624 ( 
.A(n_2118),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2063),
.B(n_1685),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2186),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2035),
.B(n_1809),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2041),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2171),
.B(n_1966),
.Y(n_2629)
);

INVxp33_ASAP7_75t_L g2630 ( 
.A(n_2181),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2151),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2035),
.B(n_1809),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2041),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2071),
.B(n_1821),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2042),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2042),
.Y(n_2636)
);

XOR2xp5_ASAP7_75t_L g2637 ( 
.A(n_2329),
.B(n_1572),
.Y(n_2637)
);

INVx2_ASAP7_75t_SL g2638 ( 
.A(n_2265),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2047),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2120),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2045),
.B(n_1821),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2047),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2040),
.Y(n_2643)
);

NAND2xp33_ASAP7_75t_R g2644 ( 
.A(n_2044),
.B(n_1586),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2040),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2160),
.B(n_1821),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2055),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2316),
.B(n_1942),
.Y(n_2648)
);

BUFx2_ASAP7_75t_L g2649 ( 
.A(n_2201),
.Y(n_2649)
);

INVxp67_ASAP7_75t_SL g2650 ( 
.A(n_2069),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2055),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2056),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2152),
.B(n_1942),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2153),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2056),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2069),
.B(n_1698),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2143),
.B(n_1701),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2185),
.B(n_1739),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2321),
.B(n_1603),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2057),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2057),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2058),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2058),
.Y(n_2663)
);

CKINVDCx20_ASAP7_75t_R g2664 ( 
.A(n_2281),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2271),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2095),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2127),
.B(n_1640),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2060),
.Y(n_2668)
);

INVxp67_ASAP7_75t_SL g2669 ( 
.A(n_2069),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2060),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2341),
.B(n_1739),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2065),
.Y(n_2672)
);

CKINVDCx16_ASAP7_75t_R g2673 ( 
.A(n_2153),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2065),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2066),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2066),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2102),
.B(n_1739),
.Y(n_2677)
);

NAND2x1p5_ASAP7_75t_L g2678 ( 
.A(n_2075),
.B(n_1925),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2048),
.B(n_1390),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2072),
.Y(n_2680)
);

XOR2xp5_ASAP7_75t_L g2681 ( 
.A(n_2192),
.B(n_1077),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2072),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2075),
.B(n_1738),
.Y(n_2683)
);

INVxp67_ASAP7_75t_SL g2684 ( 
.A(n_2075),
.Y(n_2684)
);

NOR2x1_ASAP7_75t_L g2685 ( 
.A(n_2194),
.B(n_1929),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2152),
.B(n_1942),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2121),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2152),
.B(n_1942),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2285),
.Y(n_2689)
);

INVxp33_ASAP7_75t_SL g2690 ( 
.A(n_2099),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2073),
.Y(n_2691)
);

INVxp33_ASAP7_75t_L g2692 ( 
.A(n_2309),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2073),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2080),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2080),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2091),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2091),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2233),
.B(n_1750),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2422),
.B(n_2201),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2397),
.A2(n_2201),
.B1(n_1532),
.B2(n_1582),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2630),
.B(n_1077),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_L g2702 ( 
.A(n_2356),
.B(n_1515),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_2473),
.A2(n_2201),
.B1(n_2088),
.B2(n_2285),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2368),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2422),
.B(n_2201),
.Y(n_2705)
);

INVxp67_ASAP7_75t_SL g2706 ( 
.A(n_2353),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2350),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2671),
.B(n_2201),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2356),
.B(n_1515),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2393),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2671),
.B(n_2285),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2556),
.B(n_1520),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2690),
.B(n_2251),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2399),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2427),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2391),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2492),
.B(n_2285),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2446),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2492),
.B(n_2285),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2444),
.B(n_2285),
.Y(n_2720)
);

NAND2xp33_ASAP7_75t_L g2721 ( 
.A(n_2400),
.B(n_2008),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2349),
.Y(n_2722)
);

NOR3xp33_ASAP7_75t_L g2723 ( 
.A(n_2659),
.B(n_2225),
.C(n_2036),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2444),
.B(n_2243),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2367),
.B(n_1543),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2352),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2374),
.B(n_2245),
.Y(n_2727)
);

AOI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_2532),
.A2(n_1942),
.B1(n_2254),
.B2(n_1356),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2355),
.B(n_1750),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2430),
.B(n_1750),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2366),
.B(n_1752),
.Y(n_2731)
);

NOR2xp67_ASAP7_75t_L g2732 ( 
.A(n_2481),
.B(n_1532),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2452),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2378),
.B(n_1752),
.Y(n_2734)
);

A2O1A1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2482),
.A2(n_2439),
.B(n_2384),
.C(n_2462),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2383),
.B(n_1752),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2388),
.B(n_2121),
.Y(n_2737)
);

NAND2xp33_ASAP7_75t_SL g2738 ( 
.A(n_2624),
.B(n_2307),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2591),
.B(n_2145),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2390),
.B(n_2145),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2435),
.B(n_1543),
.Y(n_2741)
);

AOI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2348),
.A2(n_2337),
.B(n_2213),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2499),
.B(n_2692),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2359),
.Y(n_2744)
);

INVxp67_ASAP7_75t_L g2745 ( 
.A(n_2395),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2360),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2395),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2520),
.B(n_2226),
.Y(n_2748)
);

A2O1A1Ixp33_ASAP7_75t_L g2749 ( 
.A1(n_2482),
.A2(n_2179),
.B(n_2116),
.C(n_2101),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2396),
.B(n_2300),
.Y(n_2750)
);

OAI22xp5_ASAP7_75t_L g2751 ( 
.A1(n_2540),
.A2(n_2154),
.B1(n_2008),
.B2(n_2025),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2348),
.A2(n_2189),
.B(n_2184),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2453),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2364),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2520),
.B(n_2226),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2484),
.B(n_2250),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2526),
.B(n_2456),
.Y(n_2757)
);

AND2x2_ASAP7_75t_SL g2758 ( 
.A(n_2471),
.B(n_2101),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2526),
.B(n_2478),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2483),
.B(n_2250),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2592),
.B(n_1384),
.Y(n_2761)
);

AOI221xp5_ASAP7_75t_L g2762 ( 
.A1(n_2679),
.A2(n_1321),
.B1(n_1310),
.B2(n_1010),
.C(n_1164),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2518),
.A2(n_1582),
.B1(n_1608),
.B2(n_1541),
.Y(n_2763)
);

AOI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2544),
.A2(n_2539),
.B1(n_2681),
.B2(n_2508),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2461),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2625),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_SL g2767 ( 
.A(n_2477),
.B(n_1783),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2592),
.B(n_1387),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2598),
.B(n_1942),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2598),
.B(n_1415),
.Y(n_2770)
);

INVx8_ASAP7_75t_L g2771 ( 
.A(n_2400),
.Y(n_2771)
);

INVx3_ASAP7_75t_L g2772 ( 
.A(n_2350),
.Y(n_2772)
);

INVx2_ASAP7_75t_SL g2773 ( 
.A(n_2394),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_L g2774 ( 
.A1(n_2471),
.A2(n_1354),
.B1(n_2105),
.B2(n_2092),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2629),
.B(n_2190),
.Y(n_2775)
);

BUFx3_ASAP7_75t_L g2776 ( 
.A(n_2488),
.Y(n_2776)
);

AND3x1_ASAP7_75t_L g2777 ( 
.A(n_2607),
.B(n_1797),
.C(n_1783),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2629),
.B(n_2190),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2384),
.B(n_2190),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2523),
.B(n_2304),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2546),
.B(n_2318),
.Y(n_2781)
);

OAI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2540),
.A2(n_2008),
.B1(n_2025),
.B2(n_2022),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2362),
.B(n_2345),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2357),
.A2(n_2092),
.B1(n_2106),
.B2(n_2105),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2362),
.B(n_1398),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2548),
.B(n_1518),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2582),
.B(n_2585),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2380),
.B(n_1570),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2350),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2380),
.B(n_1570),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2536),
.B(n_1355),
.Y(n_2791)
);

INVxp67_ASAP7_75t_L g2792 ( 
.A(n_2450),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2536),
.B(n_1395),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_SL g2794 ( 
.A(n_2582),
.B(n_2095),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2585),
.B(n_2095),
.Y(n_2795)
);

INVx5_ASAP7_75t_L g2796 ( 
.A(n_2400),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2627),
.B(n_2128),
.Y(n_2797)
);

INVx3_ASAP7_75t_L g2798 ( 
.A(n_2494),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2543),
.A2(n_1608),
.B1(n_1613),
.B2(n_1541),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2551),
.B(n_1421),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2551),
.B(n_1449),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2560),
.B(n_1523),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2591),
.B(n_2279),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2375),
.B(n_1454),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2377),
.B(n_1467),
.Y(n_2805)
);

AND2x6_ASAP7_75t_SL g2806 ( 
.A(n_2369),
.B(n_1783),
.Y(n_2806)
);

AOI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2510),
.A2(n_1614),
.B1(n_1624),
.B2(n_1613),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2698),
.B(n_1654),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2627),
.B(n_2128),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2667),
.B(n_1614),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2541),
.A2(n_2025),
.B1(n_2022),
.B2(n_2049),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2698),
.B(n_2632),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2632),
.B(n_2128),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2541),
.A2(n_2022),
.B1(n_2177),
.B2(n_2049),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2646),
.B(n_2207),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2640),
.B(n_1624),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2433),
.B(n_2116),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2357),
.A2(n_2106),
.B1(n_2112),
.B2(n_2108),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2468),
.Y(n_2819)
);

NAND2x1_ASAP7_75t_L g2820 ( 
.A(n_2666),
.B(n_2224),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2646),
.B(n_2217),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2590),
.B(n_1366),
.Y(n_2822)
);

NAND2xp33_ASAP7_75t_L g2823 ( 
.A(n_2400),
.B(n_2177),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2433),
.B(n_2568),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2439),
.A2(n_2108),
.B1(n_2114),
.B2(n_2112),
.Y(n_2825)
);

OR2x6_ASAP7_75t_L g2826 ( 
.A(n_2649),
.B(n_2343),
.Y(n_2826)
);

INVxp33_ASAP7_75t_L g2827 ( 
.A(n_2533),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2590),
.B(n_1366),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2425),
.A2(n_2179),
.B1(n_935),
.B2(n_941),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2472),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2658),
.B(n_1523),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2503),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2406),
.B(n_2046),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2658),
.B(n_1537),
.Y(n_2834)
);

NAND3xp33_ASAP7_75t_L g2835 ( 
.A(n_2677),
.B(n_2213),
.C(n_2052),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2561),
.B(n_2621),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2621),
.B(n_1447),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2612),
.B(n_1537),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_SL g2839 ( 
.A(n_2401),
.B(n_874),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2470),
.A2(n_2123),
.B1(n_2129),
.B2(n_2114),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2365),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2599),
.B(n_1589),
.Y(n_2842)
);

AOI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2425),
.A2(n_972),
.B1(n_2019),
.B2(n_2011),
.Y(n_2843)
);

BUFx3_ASAP7_75t_L g2844 ( 
.A(n_2449),
.Y(n_2844)
);

NOR2xp67_ASAP7_75t_L g2845 ( 
.A(n_2354),
.B(n_2311),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2612),
.B(n_1589),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2505),
.B(n_1609),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2505),
.A2(n_2511),
.B1(n_2440),
.B2(n_2400),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_2601),
.B(n_2053),
.Y(n_2849)
);

INVxp67_ASAP7_75t_L g2850 ( 
.A(n_2634),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2505),
.B(n_1609),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2505),
.B(n_1501),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2516),
.Y(n_2853)
);

BUFx5_ASAP7_75t_L g2854 ( 
.A(n_2434),
.Y(n_2854)
);

INVx2_ASAP7_75t_SL g2855 ( 
.A(n_2479),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2505),
.B(n_1501),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2370),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2605),
.B(n_2059),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_SL g2859 ( 
.A(n_2552),
.B(n_2059),
.Y(n_2859)
);

HB1xp67_ASAP7_75t_L g2860 ( 
.A(n_2689),
.Y(n_2860)
);

OR2x2_ASAP7_75t_L g2861 ( 
.A(n_2386),
.B(n_998),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2527),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2552),
.B(n_2578),
.Y(n_2863)
);

AND2x6_ASAP7_75t_SL g2864 ( 
.A(n_2421),
.B(n_1161),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2462),
.B(n_2206),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2371),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2474),
.A2(n_2123),
.B1(n_2133),
.B2(n_2129),
.Y(n_2867)
);

NOR2xp67_ASAP7_75t_L g2868 ( 
.A(n_2358),
.B(n_2331),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2361),
.B(n_2059),
.Y(n_2869)
);

AND2x2_ASAP7_75t_SL g2870 ( 
.A(n_2555),
.B(n_2267),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2373),
.Y(n_2871)
);

NOR3xp33_ASAP7_75t_L g2872 ( 
.A(n_2677),
.B(n_1333),
.C(n_2235),
.Y(n_2872)
);

BUFx2_ASAP7_75t_L g2873 ( 
.A(n_2372),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2419),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2494),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2361),
.B(n_2070),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2634),
.B(n_1501),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2641),
.B(n_2206),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2641),
.B(n_2206),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2440),
.B(n_2230),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2420),
.B(n_2230),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2423),
.B(n_2230),
.Y(n_2882)
);

NOR2x1p5_ASAP7_75t_L g2883 ( 
.A(n_2557),
.B(n_2286),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2424),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2494),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2426),
.B(n_2239),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2689),
.B(n_2070),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2429),
.B(n_2239),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2475),
.A2(n_2138),
.B1(n_2139),
.B2(n_2133),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2431),
.Y(n_2890)
);

INVxp67_ASAP7_75t_L g2891 ( 
.A(n_2528),
.Y(n_2891)
);

NOR2xp67_ASAP7_75t_L g2892 ( 
.A(n_2687),
.B(n_2239),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2466),
.B(n_2272),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2531),
.Y(n_2894)
);

INVx2_ASAP7_75t_SL g2895 ( 
.A(n_2673),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2637),
.B(n_2507),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2432),
.B(n_2272),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2507),
.B(n_2272),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2545),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2515),
.B(n_2290),
.Y(n_2900)
);

AOI221xp5_ASAP7_75t_L g2901 ( 
.A1(n_2515),
.A2(n_1168),
.B1(n_1172),
.B2(n_1170),
.C(n_1165),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2436),
.B(n_2290),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2437),
.B(n_2290),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2476),
.A2(n_2139),
.B1(n_2141),
.B2(n_2138),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2441),
.B(n_2308),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2442),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2480),
.B(n_1017),
.Y(n_2907)
);

INVx2_ASAP7_75t_SL g2908 ( 
.A(n_2654),
.Y(n_2908)
);

OAI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2353),
.A2(n_1652),
.B1(n_660),
.B2(n_664),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2638),
.B(n_2308),
.Y(n_2910)
);

OR2x6_ASAP7_75t_L g2911 ( 
.A(n_2665),
.B(n_2319),
.Y(n_2911)
);

AND2x4_ASAP7_75t_SL g2912 ( 
.A(n_2376),
.B(n_2308),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2558),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2562),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2445),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2664),
.B(n_2311),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2447),
.B(n_2311),
.Y(n_2917)
);

INVxp67_ASAP7_75t_L g2918 ( 
.A(n_2528),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2412),
.B(n_1392),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2451),
.B(n_2331),
.Y(n_2920)
);

AND2x6_ASAP7_75t_L g2921 ( 
.A(n_2666),
.B(n_2070),
.Y(n_2921)
);

AOI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2434),
.A2(n_2087),
.B1(n_2074),
.B2(n_2083),
.Y(n_2922)
);

NAND2xp33_ASAP7_75t_L g2923 ( 
.A(n_2434),
.B(n_2500),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2454),
.B(n_2331),
.Y(n_2924)
);

INVx2_ASAP7_75t_SL g2925 ( 
.A(n_2685),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2455),
.B(n_2140),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2458),
.B(n_2140),
.Y(n_2927)
);

BUFx5_ASAP7_75t_L g2928 ( 
.A(n_2434),
.Y(n_2928)
);

OAI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2379),
.A2(n_667),
.B1(n_668),
.B2(n_654),
.Y(n_2929)
);

AOI221xp5_ASAP7_75t_L g2930 ( 
.A1(n_2443),
.A2(n_1176),
.B1(n_1182),
.B2(n_1174),
.C(n_1173),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2579),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2581),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2528),
.B(n_2549),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2434),
.A2(n_2074),
.B1(n_2083),
.B2(n_2076),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2596),
.Y(n_2935)
);

A2O1A1Ixp33_ASAP7_75t_L g2936 ( 
.A1(n_2648),
.A2(n_2229),
.B(n_2259),
.C(n_2222),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2528),
.B(n_1644),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2553),
.B(n_1805),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2600),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_2500),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2351),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2528),
.B(n_1647),
.Y(n_2942)
);

OAI22xp33_ASAP7_75t_L g2943 ( 
.A1(n_2379),
.A2(n_680),
.B1(n_687),
.B2(n_676),
.Y(n_2943)
);

AOI22xp33_ASAP7_75t_L g2944 ( 
.A1(n_2486),
.A2(n_2142),
.B1(n_2147),
.B2(n_2141),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2602),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2549),
.B(n_1648),
.Y(n_2946)
);

BUFx8_ASAP7_75t_L g2947 ( 
.A(n_2448),
.Y(n_2947)
);

NOR2x1p5_ASAP7_75t_L g2948 ( 
.A(n_2428),
.B(n_1492),
.Y(n_2948)
);

INVx2_ASAP7_75t_SL g2949 ( 
.A(n_2363),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2554),
.B(n_1834),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2593),
.Y(n_2951)
);

OR2x6_ASAP7_75t_L g2952 ( 
.A(n_2610),
.B(n_2319),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2613),
.B(n_2074),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2613),
.B(n_2076),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2650),
.B(n_2076),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2594),
.Y(n_2956)
);

BUFx3_ASAP7_75t_L g2957 ( 
.A(n_2589),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2650),
.B(n_2083),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2443),
.B(n_2252),
.Y(n_2959)
);

OAI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2413),
.A2(n_693),
.B1(n_696),
.B2(n_690),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2595),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2413),
.B(n_2252),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2490),
.B(n_1392),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2549),
.B(n_2142),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2549),
.B(n_2147),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2487),
.A2(n_2159),
.B1(n_2162),
.B2(n_2156),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2626),
.B(n_1834),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2603),
.B(n_2275),
.Y(n_2968)
);

OAI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2438),
.A2(n_700),
.B1(n_703),
.B2(n_699),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2549),
.B(n_2156),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2489),
.A2(n_2162),
.B1(n_2163),
.B2(n_2159),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2604),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2606),
.B(n_2163),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2669),
.B(n_2208),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2662),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2597),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2608),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2672),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2609),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2611),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2615),
.Y(n_2981)
);

CKINVDCx5p33_ASAP7_75t_R g2982 ( 
.A(n_2485),
.Y(n_2982)
);

A2O1A1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_2648),
.A2(n_2263),
.B(n_2195),
.C(n_2235),
.Y(n_2983)
);

BUFx6f_ASAP7_75t_L g2984 ( 
.A(n_2500),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2669),
.B(n_2208),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2620),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2616),
.B(n_2164),
.Y(n_2987)
);

AOI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2438),
.A2(n_2312),
.B1(n_2313),
.B2(n_2224),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2617),
.B(n_2164),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2502),
.B(n_1392),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2491),
.A2(n_2495),
.B1(n_2496),
.B2(n_2493),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2618),
.B(n_2167),
.Y(n_2992)
);

NOR2xp33_ASAP7_75t_L g2993 ( 
.A(n_2619),
.B(n_2253),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2622),
.B(n_2167),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2623),
.B(n_2269),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_SL g2996 ( 
.A1(n_2485),
.A2(n_707),
.B1(n_710),
.B2(n_704),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2497),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2684),
.B(n_2208),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2501),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2693),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2504),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2684),
.B(n_2208),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2381),
.B(n_2382),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2385),
.B(n_2168),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2387),
.B(n_2168),
.Y(n_3005)
);

AND2x6_ASAP7_75t_SL g3006 ( 
.A(n_2534),
.B(n_1185),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2389),
.B(n_2170),
.Y(n_3007)
);

CKINVDCx20_ASAP7_75t_R g3008 ( 
.A(n_2530),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2392),
.B(n_2170),
.Y(n_3009)
);

O2A1O1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2534),
.A2(n_1503),
.B(n_1508),
.C(n_1497),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2530),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2398),
.B(n_2270),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2402),
.B(n_2172),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2403),
.B(n_2270),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_SL g3015 ( 
.A(n_2530),
.B(n_2208),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2697),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2522),
.Y(n_3017)
);

OAI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2713),
.A2(n_2404),
.B1(n_2407),
.B2(n_2405),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2702),
.B(n_2448),
.Y(n_3019)
);

AOI21xp5_ASAP7_75t_L g3020 ( 
.A1(n_2706),
.A2(n_2498),
.B(n_2683),
.Y(n_3020)
);

AOI33xp33_ASAP7_75t_L g3021 ( 
.A1(n_2762),
.A2(n_1191),
.A3(n_1187),
.B1(n_1193),
.B2(n_1189),
.B3(n_1186),
.Y(n_3021)
);

AOI21xp33_ASAP7_75t_L g3022 ( 
.A1(n_2810),
.A2(n_2644),
.B(n_2509),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2757),
.B(n_2759),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2766),
.B(n_1396),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2836),
.B(n_2409),
.Y(n_3025)
);

OAI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2735),
.A2(n_2498),
.B(n_2569),
.Y(n_3026)
);

A2O1A1Ixp33_ASAP7_75t_L g3027 ( 
.A1(n_2837),
.A2(n_2411),
.B(n_2414),
.C(n_2410),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2706),
.A2(n_2683),
.B(n_2656),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2721),
.A2(n_2656),
.B(n_2569),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2764),
.A2(n_2506),
.B1(n_2513),
.B2(n_2512),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2749),
.A2(n_2686),
.B(n_2653),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2823),
.A2(n_2686),
.B(n_2653),
.Y(n_3032)
);

A2O1A1Ixp33_ASAP7_75t_L g3033 ( 
.A1(n_2848),
.A2(n_2416),
.B(n_2417),
.C(n_2415),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2742),
.A2(n_2688),
.B(n_2563),
.Y(n_3034)
);

NAND2x1p5_ASAP7_75t_L g3035 ( 
.A(n_2796),
.B(n_2657),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2773),
.B(n_2418),
.Y(n_3036)
);

AOI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2742),
.A2(n_2688),
.B(n_2563),
.Y(n_3037)
);

O2A1O1Ixp33_ASAP7_75t_L g3038 ( 
.A1(n_2709),
.A2(n_1516),
.B(n_1197),
.C(n_1199),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2703),
.A2(n_2525),
.B1(n_2529),
.B2(n_2524),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2751),
.A2(n_2631),
.B(n_2457),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2730),
.B(n_2514),
.Y(n_3041)
);

CKINVDCx11_ASAP7_75t_R g3042 ( 
.A(n_2806),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2812),
.B(n_2566),
.Y(n_3043)
);

OAI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2779),
.A2(n_2564),
.B(n_2521),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2758),
.B(n_2566),
.Y(n_3045)
);

AOI21xp33_ASAP7_75t_L g3046 ( 
.A1(n_2929),
.A2(n_2644),
.B(n_2517),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_SL g3047 ( 
.A(n_2758),
.B(n_2566),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2782),
.A2(n_2631),
.B(n_2457),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2754),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2919),
.B(n_1396),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2764),
.A2(n_2469),
.B1(n_2537),
.B2(n_2535),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2841),
.Y(n_3052)
);

OAI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2835),
.A2(n_2564),
.B(n_2519),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2923),
.A2(n_2144),
.B(n_2135),
.Y(n_3054)
);

A2O1A1Ixp33_ASAP7_75t_L g3055 ( 
.A1(n_2711),
.A2(n_2542),
.B(n_2547),
.C(n_2538),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2752),
.A2(n_2209),
.B(n_2175),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2701),
.B(n_2469),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2865),
.A2(n_2460),
.B(n_2459),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2863),
.B(n_2330),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2811),
.A2(n_2276),
.B(n_2330),
.Y(n_3060)
);

AO21x1_ASAP7_75t_L g3061 ( 
.A1(n_2962),
.A2(n_2559),
.B(n_2550),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_3017),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2775),
.A2(n_2335),
.B(n_2330),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2704),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2710),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2857),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_2796),
.B(n_2330),
.Y(n_3067)
);

OAI21xp33_ASAP7_75t_L g3068 ( 
.A1(n_2839),
.A2(n_744),
.B(n_726),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2714),
.Y(n_3069)
);

AOI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2778),
.A2(n_2335),
.B(n_2330),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2850),
.B(n_2743),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2850),
.B(n_2565),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2796),
.B(n_2335),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2745),
.B(n_2567),
.Y(n_3074)
);

INVx4_ASAP7_75t_L g3075 ( 
.A(n_2796),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2789),
.Y(n_3076)
);

O2A1O1Ixp33_ASAP7_75t_L g3077 ( 
.A1(n_2817),
.A2(n_1201),
.B(n_1204),
.C(n_1196),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2745),
.B(n_2570),
.Y(n_3078)
);

BUFx3_ASAP7_75t_L g3079 ( 
.A(n_2716),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2814),
.A2(n_2342),
.B(n_2335),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2715),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2898),
.A2(n_2342),
.B(n_2335),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2747),
.B(n_2571),
.Y(n_3083)
);

INVxp67_ASAP7_75t_L g3084 ( 
.A(n_2963),
.Y(n_3084)
);

A2O1A1Ixp33_ASAP7_75t_L g3085 ( 
.A1(n_2703),
.A2(n_2573),
.B(n_2574),
.C(n_2572),
.Y(n_3085)
);

NOR2x1_ASAP7_75t_L g3086 ( 
.A(n_2844),
.B(n_2575),
.Y(n_3086)
);

AOI21xp33_ASAP7_75t_L g3087 ( 
.A1(n_2909),
.A2(n_2328),
.B(n_2576),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2747),
.B(n_2580),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2866),
.Y(n_3089)
);

A2O1A1Ixp33_ASAP7_75t_L g3090 ( 
.A1(n_3003),
.A2(n_2584),
.B(n_2586),
.C(n_2583),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2724),
.A2(n_2588),
.B1(n_2587),
.B2(n_2464),
.Y(n_3091)
);

INVxp67_ASAP7_75t_L g3092 ( 
.A(n_2824),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2761),
.B(n_2463),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2768),
.B(n_2465),
.Y(n_3094)
);

O2A1O1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2929),
.A2(n_1208),
.B(n_1211),
.C(n_1206),
.Y(n_3095)
);

OAI321xp33_ASAP7_75t_L g3096 ( 
.A1(n_2829),
.A2(n_1325),
.A3(n_1326),
.B1(n_1324),
.B2(n_1297),
.C(n_1294),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2900),
.A2(n_2342),
.B(n_2336),
.Y(n_3097)
);

AND2x2_ASAP7_75t_SL g3098 ( 
.A(n_2777),
.B(n_2012),
.Y(n_3098)
);

INVx4_ASAP7_75t_L g3099 ( 
.A(n_2771),
.Y(n_3099)
);

BUFx2_ASAP7_75t_L g3100 ( 
.A(n_2776),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2896),
.B(n_2467),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2708),
.B(n_2336),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2959),
.A2(n_2342),
.B(n_2336),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2871),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2959),
.A2(n_2342),
.B(n_2336),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2722),
.Y(n_3106)
);

INVx1_ASAP7_75t_SL g3107 ( 
.A(n_3008),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2865),
.A2(n_2336),
.B(n_2324),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2718),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2748),
.A2(n_2324),
.B(n_2224),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2990),
.B(n_1396),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2755),
.A2(n_2324),
.B(n_2249),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_2808),
.B(n_1472),
.Y(n_3113)
);

OAI21xp33_ASAP7_75t_L g3114 ( 
.A1(n_2943),
.A2(n_2969),
.B(n_2960),
.Y(n_3114)
);

A2O1A1Ixp33_ASAP7_75t_L g3115 ( 
.A1(n_2833),
.A2(n_1723),
.B(n_1724),
.C(n_1713),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2733),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_2739),
.B(n_2249),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2770),
.B(n_1403),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2726),
.Y(n_3119)
);

OAI21x1_ASAP7_75t_SL g3120 ( 
.A1(n_2880),
.A2(n_2178),
.B(n_2253),
.Y(n_3120)
);

INVx3_ASAP7_75t_L g3121 ( 
.A(n_2771),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2907),
.B(n_1403),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2727),
.B(n_1403),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2962),
.A2(n_2249),
.B(n_2408),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2762),
.B(n_1414),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2753),
.Y(n_3126)
);

NAND2xp33_ASAP7_75t_L g3127 ( 
.A(n_2921),
.B(n_2408),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2842),
.B(n_1414),
.Y(n_3128)
);

AOI211xp5_ASAP7_75t_L g3129 ( 
.A1(n_2996),
.A2(n_1213),
.B(n_1214),
.C(n_1212),
.Y(n_3129)
);

AOI21x1_ASAP7_75t_L g3130 ( 
.A1(n_2974),
.A2(n_2020),
.B(n_2013),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2699),
.A2(n_2249),
.B(n_2577),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2744),
.Y(n_3132)
);

BUFx3_ASAP7_75t_L g3133 ( 
.A(n_2947),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_2864),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2746),
.Y(n_3135)
);

HB1xp67_ASAP7_75t_L g3136 ( 
.A(n_2792),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2705),
.A2(n_2249),
.B(n_2577),
.Y(n_3137)
);

NOR3xp33_ASAP7_75t_L g3138 ( 
.A(n_2943),
.B(n_1218),
.C(n_1216),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_2861),
.B(n_2873),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2822),
.B(n_1474),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2794),
.A2(n_2614),
.B(n_2328),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_2893),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2786),
.B(n_1414),
.Y(n_3143)
);

A2O1A1Ixp33_ASAP7_75t_L g3144 ( 
.A1(n_2950),
.A2(n_1735),
.B(n_1747),
.C(n_1726),
.Y(n_3144)
);

OAI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2983),
.A2(n_1770),
.B(n_1766),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2874),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2816),
.A2(n_713),
.B1(n_714),
.B2(n_712),
.Y(n_3147)
);

AO21x1_ASAP7_75t_L g3148 ( 
.A1(n_2872),
.A2(n_2633),
.B(n_2628),
.Y(n_3148)
);

AOI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2795),
.A2(n_2614),
.B(n_2328),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2802),
.B(n_1416),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_2784),
.A2(n_2100),
.B(n_2094),
.Y(n_3151)
);

AOI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2741),
.A2(n_2712),
.B1(n_2725),
.B2(n_2843),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2792),
.B(n_1416),
.Y(n_3153)
);

AND3x1_ASAP7_75t_SL g3154 ( 
.A(n_2948),
.B(n_1221),
.C(n_1220),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2765),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2789),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2729),
.B(n_1416),
.Y(n_3157)
);

A2O1A1Ixp33_ASAP7_75t_L g3158 ( 
.A1(n_3010),
.A2(n_1785),
.B(n_1786),
.C(n_1771),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2731),
.B(n_1430),
.Y(n_3159)
);

O2A1O1Ixp5_ASAP7_75t_L g3160 ( 
.A1(n_2787),
.A2(n_1791),
.B(n_1793),
.C(n_1787),
.Y(n_3160)
);

NOR2x1_ASAP7_75t_R g3161 ( 
.A(n_2982),
.B(n_716),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2815),
.B(n_2635),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2734),
.B(n_1430),
.Y(n_3163)
);

AO21x1_ASAP7_75t_L g3164 ( 
.A1(n_2872),
.A2(n_2639),
.B(n_2636),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_2737),
.Y(n_3165)
);

INVxp67_ASAP7_75t_L g3166 ( 
.A(n_2780),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2797),
.A2(n_2107),
.B(n_2104),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2809),
.A2(n_2146),
.B(n_2110),
.Y(n_3168)
);

NOR2x1p5_ASAP7_75t_SL g3169 ( 
.A(n_2854),
.B(n_2148),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2750),
.B(n_1430),
.Y(n_3170)
);

INVx3_ASAP7_75t_L g3171 ( 
.A(n_2771),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2819),
.Y(n_3172)
);

BUFx4f_ASAP7_75t_L g3173 ( 
.A(n_2870),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2813),
.A2(n_2150),
.B(n_2678),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2739),
.B(n_2642),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2926),
.A2(n_2678),
.B(n_2645),
.Y(n_3176)
);

AOI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2781),
.A2(n_2803),
.B1(n_2828),
.B2(n_2916),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2736),
.B(n_1440),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_2927),
.A2(n_2647),
.B(n_2643),
.Y(n_3179)
);

NOR2xp67_ASAP7_75t_L g3180 ( 
.A(n_2908),
.B(n_2651),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2740),
.B(n_1440),
.Y(n_3181)
);

INVx2_ASAP7_75t_SL g3182 ( 
.A(n_2947),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2827),
.B(n_1475),
.Y(n_3183)
);

O2A1O1Ixp5_ASAP7_75t_L g3184 ( 
.A1(n_2985),
.A2(n_1803),
.B(n_1804),
.C(n_1794),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2998),
.A2(n_2655),
.B(n_2652),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2830),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2800),
.B(n_1440),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_2821),
.B(n_2660),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_L g3189 ( 
.A(n_2803),
.B(n_721),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_2789),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_SL g3191 ( 
.A(n_2717),
.B(n_2661),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2801),
.B(n_1469),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_3002),
.A2(n_2668),
.B(n_2663),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2884),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2953),
.A2(n_2674),
.B(n_2670),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2912),
.B(n_1469),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2890),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_2954),
.A2(n_2676),
.B(n_2675),
.Y(n_3198)
);

AOI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_2955),
.A2(n_2682),
.B(n_2680),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2760),
.B(n_1469),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2855),
.B(n_727),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2958),
.A2(n_2694),
.B(n_2691),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2906),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2915),
.B(n_1470),
.Y(n_3204)
);

HB1xp67_ASAP7_75t_L g3205 ( 
.A(n_2860),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_2938),
.A2(n_2696),
.B(n_2695),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_2719),
.B(n_2720),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2935),
.B(n_1470),
.Y(n_3208)
);

OAI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3010),
.A2(n_1812),
.B(n_1806),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2936),
.A2(n_2297),
.B(n_2295),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2939),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2945),
.B(n_1470),
.Y(n_3212)
);

INVx11_ASAP7_75t_L g3213 ( 
.A(n_2921),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2700),
.B(n_730),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2832),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_2986),
.B(n_1481),
.Y(n_3216)
);

OAI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_2972),
.A2(n_1225),
.B1(n_1228),
.B2(n_1223),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2853),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2941),
.B(n_731),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_2870),
.B(n_2269),
.Y(n_3220)
);

INVxp67_ASAP7_75t_L g3221 ( 
.A(n_2949),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2977),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2979),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_2878),
.A2(n_2297),
.B(n_2295),
.Y(n_3224)
);

OR2x6_ASAP7_75t_L g3225 ( 
.A(n_2826),
.B(n_2227),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2879),
.A2(n_2306),
.B(n_2301),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_2937),
.A2(n_2306),
.B(n_2301),
.Y(n_3227)
);

AO21x1_ASAP7_75t_L g3228 ( 
.A1(n_2909),
.A2(n_1822),
.B(n_1820),
.Y(n_3228)
);

OR2x6_ASAP7_75t_L g3229 ( 
.A(n_2826),
.B(n_2287),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2980),
.B(n_1481),
.Y(n_3230)
);

AO21x1_ASAP7_75t_L g3231 ( 
.A1(n_2967),
.A2(n_1831),
.B(n_1825),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2862),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_2957),
.B(n_1481),
.Y(n_3233)
);

AND2x4_ASAP7_75t_L g3234 ( 
.A(n_2826),
.B(n_2883),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_2976),
.B(n_2895),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2981),
.B(n_1498),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_2891),
.B(n_2273),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2942),
.A2(n_2320),
.B(n_2310),
.Y(n_3238)
);

NOR3xp33_ASAP7_75t_L g3239 ( 
.A(n_2960),
.B(n_1231),
.C(n_1229),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2901),
.B(n_1498),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2997),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2901),
.B(n_1498),
.Y(n_3242)
);

OAI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_2969),
.A2(n_1249),
.B1(n_1250),
.B2(n_1234),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2946),
.A2(n_1833),
.B(n_1832),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3015),
.A2(n_2320),
.B(n_2310),
.Y(n_3245)
);

OAI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2922),
.A2(n_1844),
.B(n_1836),
.Y(n_3246)
);

BUFx3_ASAP7_75t_L g3247 ( 
.A(n_3011),
.Y(n_3247)
);

OR2x2_ASAP7_75t_L g3248 ( 
.A(n_2785),
.B(n_1538),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2723),
.B(n_1517),
.Y(n_3249)
);

AO21x1_ASAP7_75t_L g3250 ( 
.A1(n_2769),
.A2(n_1850),
.B(n_1847),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3023),
.B(n_3025),
.Y(n_3251)
);

OAI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3114),
.A2(n_2723),
.B(n_2910),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3101),
.B(n_2999),
.Y(n_3253)
);

OAI21xp33_ASAP7_75t_L g3254 ( 
.A1(n_3214),
.A2(n_2799),
.B(n_2763),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3071),
.B(n_3001),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3127),
.A2(n_2820),
.B(n_2881),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3049),
.Y(n_3257)
);

AOI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_3020),
.A2(n_2886),
.B(n_2882),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3165),
.B(n_2791),
.Y(n_3259)
);

BUFx12f_ASAP7_75t_L g3260 ( 
.A(n_3042),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3152),
.A2(n_2807),
.B1(n_2728),
.B2(n_2934),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3052),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3205),
.B(n_2793),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_3029),
.A2(n_2897),
.B(n_2888),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3066),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_SL g3266 ( 
.A(n_3173),
.B(n_2767),
.Y(n_3266)
);

A2O1A1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_3113),
.A2(n_3140),
.B(n_3018),
.C(n_3068),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3103),
.A2(n_2903),
.B(n_2902),
.Y(n_3268)
);

AND2x6_ASAP7_75t_SL g3269 ( 
.A(n_3019),
.B(n_1251),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3089),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3050),
.B(n_1255),
.Y(n_3271)
);

O2A1O1Ixp33_ASAP7_75t_SL g3272 ( 
.A1(n_3027),
.A2(n_2859),
.B(n_2756),
.C(n_2858),
.Y(n_3272)
);

BUFx12f_ASAP7_75t_L g3273 ( 
.A(n_3182),
.Y(n_3273)
);

AOI22xp5_ASAP7_75t_L g3274 ( 
.A1(n_3243),
.A2(n_2738),
.B1(n_2732),
.B2(n_2783),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_3105),
.A2(n_2917),
.B(n_2905),
.Y(n_3275)
);

OR2x2_ASAP7_75t_L g3276 ( 
.A(n_3139),
.B(n_2860),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_3142),
.B(n_2849),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_3107),
.B(n_3106),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3062),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_L g3280 ( 
.A(n_3221),
.B(n_732),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3064),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3026),
.A2(n_2924),
.B(n_2920),
.Y(n_3282)
);

BUFx3_ASAP7_75t_L g3283 ( 
.A(n_3079),
.Y(n_3283)
);

OR2x6_ASAP7_75t_L g3284 ( 
.A(n_3133),
.B(n_2925),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3093),
.B(n_2831),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_3173),
.B(n_2885),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3094),
.B(n_2834),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3122),
.B(n_1257),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_3243),
.A2(n_2728),
.B1(n_2918),
.B2(n_2891),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_3107),
.B(n_737),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3136),
.B(n_2930),
.Y(n_3291)
);

AOI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3018),
.A2(n_2918),
.B1(n_2774),
.B2(n_2868),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3104),
.Y(n_3293)
);

AOI22x1_ASAP7_75t_L g3294 ( 
.A1(n_3058),
.A2(n_2772),
.B1(n_2798),
.B2(n_2707),
.Y(n_3294)
);

BUFx2_ASAP7_75t_L g3295 ( 
.A(n_3100),
.Y(n_3295)
);

O2A1O1Ixp33_ASAP7_75t_SL g3296 ( 
.A1(n_3033),
.A2(n_2856),
.B(n_2852),
.C(n_2851),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3036),
.B(n_2930),
.Y(n_3297)
);

INVx3_ASAP7_75t_L g3298 ( 
.A(n_3213),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3026),
.A2(n_2933),
.B(n_3012),
.Y(n_3299)
);

CKINVDCx8_ASAP7_75t_R g3300 ( 
.A(n_3134),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_3247),
.Y(n_3301)
);

O2A1O1Ixp33_ASAP7_75t_L g3302 ( 
.A1(n_3138),
.A2(n_2869),
.B(n_2876),
.C(n_2847),
.Y(n_3302)
);

AOI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3177),
.A2(n_2774),
.B1(n_2911),
.B2(n_2846),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3091),
.A2(n_3014),
.B(n_3005),
.Y(n_3304)
);

BUFx6f_ASAP7_75t_L g3305 ( 
.A(n_3117),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_3183),
.B(n_3219),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3119),
.Y(n_3307)
);

BUFx6f_ASAP7_75t_L g3308 ( 
.A(n_3117),
.Y(n_3308)
);

NOR2xp67_ASAP7_75t_L g3309 ( 
.A(n_3075),
.B(n_2707),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3166),
.B(n_2968),
.Y(n_3310)
);

AOI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_3091),
.A2(n_3007),
.B(n_3004),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3072),
.B(n_2993),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_3111),
.B(n_1259),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3065),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_3234),
.B(n_2772),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3074),
.B(n_2995),
.Y(n_3316)
);

OR2x6_ASAP7_75t_L g3317 ( 
.A(n_3234),
.B(n_2911),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_SL g3318 ( 
.A(n_3161),
.B(n_3022),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3078),
.B(n_3006),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3132),
.Y(n_3320)
);

AO22x1_ASAP7_75t_L g3321 ( 
.A1(n_3057),
.A2(n_2838),
.B1(n_2899),
.B2(n_2894),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3083),
.B(n_3088),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3082),
.A2(n_3013),
.B(n_3009),
.Y(n_3323)
);

OAI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3147),
.A2(n_2877),
.B1(n_2788),
.B2(n_2790),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_3092),
.A2(n_2892),
.B1(n_2845),
.B2(n_2988),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_3201),
.B(n_741),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3090),
.A2(n_2911),
.B1(n_2991),
.B2(n_2825),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3170),
.B(n_1538),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3041),
.B(n_3175),
.Y(n_3329)
);

AOI21xp33_ASAP7_75t_L g3330 ( 
.A1(n_3240),
.A2(n_3242),
.B(n_3125),
.Y(n_3330)
);

BUFx12f_ASAP7_75t_L g3331 ( 
.A(n_3076),
.Y(n_3331)
);

A2O1A1Ixp33_ASAP7_75t_L g3332 ( 
.A1(n_3046),
.A2(n_3096),
.B(n_3021),
.C(n_3129),
.Y(n_3332)
);

AO32x1_ASAP7_75t_L g3333 ( 
.A1(n_3039),
.A2(n_2931),
.A3(n_2932),
.B1(n_2914),
.B2(n_2913),
.Y(n_3333)
);

OR2x2_ASAP7_75t_L g3334 ( 
.A(n_3135),
.B(n_2991),
.Y(n_3334)
);

NOR3xp33_ASAP7_75t_L g3335 ( 
.A(n_3086),
.B(n_3038),
.C(n_3096),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3175),
.B(n_1538),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3146),
.Y(n_3337)
);

AO21x1_ASAP7_75t_L g3338 ( 
.A1(n_3039),
.A2(n_2965),
.B(n_2964),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3058),
.A2(n_2825),
.B1(n_2805),
.B2(n_2804),
.Y(n_3339)
);

O2A1O1Ixp33_ASAP7_75t_SL g3340 ( 
.A1(n_3045),
.A2(n_2887),
.B(n_2970),
.C(n_2973),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3180),
.B(n_2885),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3194),
.B(n_1538),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3097),
.A2(n_3080),
.B(n_3040),
.Y(n_3343)
);

O2A1O1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_3239),
.A2(n_1265),
.B(n_1266),
.C(n_1260),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3197),
.Y(n_3345)
);

A2O1A1Ixp33_ASAP7_75t_L g3346 ( 
.A1(n_3087),
.A2(n_2989),
.B(n_2992),
.C(n_2987),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3203),
.B(n_1540),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3211),
.B(n_1540),
.Y(n_3348)
);

BUFx6f_ASAP7_75t_L g3349 ( 
.A(n_3076),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3222),
.B(n_1540),
.Y(n_3350)
);

NOR2xp33_ASAP7_75t_L g3351 ( 
.A(n_3235),
.B(n_3233),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3223),
.B(n_1540),
.Y(n_3352)
);

O2A1O1Ixp33_ASAP7_75t_L g3353 ( 
.A1(n_3095),
.A2(n_1272),
.B(n_1273),
.C(n_1269),
.Y(n_3353)
);

BUFx12f_ASAP7_75t_L g3354 ( 
.A(n_3076),
.Y(n_3354)
);

NAND2x1p5_ASAP7_75t_L g3355 ( 
.A(n_3099),
.B(n_2885),
.Y(n_3355)
);

OAI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3051),
.A2(n_3084),
.B1(n_3249),
.B2(n_3085),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_3156),
.Y(n_3357)
);

BUFx2_ASAP7_75t_L g3358 ( 
.A(n_3156),
.Y(n_3358)
);

BUFx12f_ASAP7_75t_L g3359 ( 
.A(n_3156),
.Y(n_3359)
);

A2O1A1Ixp33_ASAP7_75t_L g3360 ( 
.A1(n_3087),
.A2(n_2994),
.B(n_1853),
.C(n_1913),
.Y(n_3360)
);

BUFx12f_ASAP7_75t_L g3361 ( 
.A(n_3190),
.Y(n_3361)
);

NAND3xp33_ASAP7_75t_L g3362 ( 
.A(n_3189),
.B(n_745),
.C(n_742),
.Y(n_3362)
);

AOI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3154),
.A2(n_2928),
.B1(n_2854),
.B2(n_2952),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3056),
.A2(n_2818),
.B(n_2784),
.Y(n_3364)
);

AND2x4_ASAP7_75t_L g3365 ( 
.A(n_3225),
.B(n_2798),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3098),
.B(n_2940),
.Y(n_3366)
);

CKINVDCx5p33_ASAP7_75t_R g3367 ( 
.A(n_3216),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_3030),
.A2(n_2956),
.B1(n_2961),
.B2(n_2951),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3241),
.B(n_2975),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3128),
.B(n_2978),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3063),
.A2(n_2818),
.B(n_2875),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3070),
.A2(n_2875),
.B(n_2940),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_3225),
.B(n_2940),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3055),
.A2(n_2952),
.B1(n_2867),
.B2(n_2889),
.Y(n_3374)
);

INVx3_ASAP7_75t_L g3375 ( 
.A(n_3099),
.Y(n_3375)
);

O2A1O1Ixp33_ASAP7_75t_SL g3376 ( 
.A1(n_3047),
.A2(n_1857),
.B(n_1863),
.C(n_1852),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3069),
.Y(n_3377)
);

BUFx3_ASAP7_75t_L g3378 ( 
.A(n_3196),
.Y(n_3378)
);

BUFx6f_ASAP7_75t_L g3379 ( 
.A(n_3225),
.Y(n_3379)
);

NOR2x1p5_ASAP7_75t_SL g3380 ( 
.A(n_3130),
.B(n_2854),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3081),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_3229),
.B(n_2984),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3143),
.B(n_3000),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3108),
.A2(n_2984),
.B(n_2952),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_3153),
.B(n_746),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3150),
.B(n_3016),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_3061),
.B(n_2984),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3048),
.A2(n_2867),
.B(n_2840),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_3190),
.Y(n_3389)
);

CKINVDCx8_ASAP7_75t_R g3390 ( 
.A(n_3229),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3075),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3148),
.B(n_2854),
.Y(n_3392)
);

NAND2x1p5_ASAP7_75t_L g3393 ( 
.A(n_3121),
.B(n_2273),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3109),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_SL g3395 ( 
.A(n_3121),
.B(n_2854),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3024),
.B(n_1529),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3118),
.B(n_1531),
.Y(n_3397)
);

INVx2_ASAP7_75t_SL g3398 ( 
.A(n_3229),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3116),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_L g3400 ( 
.A(n_3123),
.B(n_752),
.Y(n_3400)
);

BUFx12f_ASAP7_75t_L g3401 ( 
.A(n_3035),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3217),
.B(n_1531),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_3164),
.B(n_2854),
.Y(n_3403)
);

OA21x2_ASAP7_75t_L g3404 ( 
.A1(n_3231),
.A2(n_2889),
.B(n_2840),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3217),
.B(n_1531),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3059),
.B(n_755),
.Y(n_3406)
);

OA22x2_ASAP7_75t_L g3407 ( 
.A1(n_3220),
.A2(n_1295),
.B1(n_1298),
.B2(n_1293),
.Y(n_3407)
);

A2O1A1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_3206),
.A2(n_1922),
.B(n_1910),
.C(n_1870),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3043),
.A2(n_2944),
.B1(n_2966),
.B2(n_2904),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_3126),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3124),
.A2(n_2904),
.B(n_2944),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3187),
.B(n_1531),
.Y(n_3412)
);

O2A1O1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3077),
.A2(n_1276),
.B(n_1277),
.C(n_1274),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3155),
.A2(n_2172),
.B1(n_2174),
.B2(n_2173),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_SL g3415 ( 
.A1(n_3192),
.A2(n_2928),
.B1(n_2921),
.B2(n_757),
.Y(n_3415)
);

O2A1O1Ixp5_ASAP7_75t_L g3416 ( 
.A1(n_3228),
.A2(n_1879),
.B(n_1882),
.C(n_1864),
.Y(n_3416)
);

O2A1O1Ixp33_ASAP7_75t_L g3417 ( 
.A1(n_3144),
.A2(n_1286),
.B(n_1288),
.C(n_1278),
.Y(n_3417)
);

A2O1A1Ixp33_ASAP7_75t_SL g3418 ( 
.A1(n_3145),
.A2(n_1290),
.B(n_1291),
.C(n_1289),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3162),
.B(n_1526),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3188),
.B(n_1526),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_3035),
.B(n_2928),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3207),
.A2(n_2928),
.B1(n_3171),
.B2(n_3191),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3172),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3060),
.A2(n_2971),
.B(n_2966),
.Y(n_3424)
);

BUFx2_ASAP7_75t_L g3425 ( 
.A(n_3171),
.Y(n_3425)
);

BUFx2_ASAP7_75t_L g3426 ( 
.A(n_3200),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3204),
.B(n_1548),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_3244),
.B(n_2928),
.Y(n_3428)
);

BUFx3_ASAP7_75t_L g3429 ( 
.A(n_3186),
.Y(n_3429)
);

AOI21x1_ASAP7_75t_L g3430 ( 
.A1(n_3250),
.A2(n_1892),
.B(n_1891),
.Y(n_3430)
);

BUFx3_ASAP7_75t_L g3431 ( 
.A(n_3215),
.Y(n_3431)
);

AND2x4_ASAP7_75t_L g3432 ( 
.A(n_3169),
.B(n_2921),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3157),
.A2(n_2971),
.B1(n_761),
.B2(n_766),
.Y(n_3433)
);

BUFx3_ASAP7_75t_L g3434 ( 
.A(n_3218),
.Y(n_3434)
);

AO21x1_ASAP7_75t_L g3435 ( 
.A1(n_3244),
.A2(n_3209),
.B(n_3237),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3248),
.B(n_1324),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3232),
.B(n_2921),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3028),
.A2(n_2928),
.B(n_2326),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_3181),
.B(n_756),
.Y(n_3439)
);

O2A1O1Ixp33_ASAP7_75t_L g3440 ( 
.A1(n_3115),
.A2(n_1308),
.B(n_1312),
.C(n_1307),
.Y(n_3440)
);

AOI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3159),
.A2(n_784),
.B1(n_796),
.B2(n_785),
.Y(n_3441)
);

OAI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3163),
.A2(n_3178),
.B1(n_3158),
.B2(n_3246),
.Y(n_3442)
);

A2O1A1Ixp33_ASAP7_75t_L g3443 ( 
.A1(n_3209),
.A2(n_1917),
.B(n_1905),
.C(n_1899),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3176),
.A2(n_2326),
.B(n_2325),
.Y(n_3444)
);

INVx3_ASAP7_75t_L g3445 ( 
.A(n_3208),
.Y(n_3445)
);

O2A1O1Ixp5_ASAP7_75t_L g3446 ( 
.A1(n_3102),
.A2(n_1901),
.B(n_1906),
.C(n_1893),
.Y(n_3446)
);

OAI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3031),
.A2(n_1916),
.B(n_1907),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3212),
.B(n_774),
.Y(n_3448)
);

HB1xp67_ASAP7_75t_L g3449 ( 
.A(n_3053),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3230),
.B(n_1548),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_3112),
.A2(n_2325),
.B(n_2278),
.Y(n_3451)
);

NOR2xp67_ASAP7_75t_L g3452 ( 
.A(n_3141),
.B(n_2275),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3236),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3179),
.B(n_1548),
.Y(n_3454)
);

NOR2xp67_ASAP7_75t_L g3455 ( 
.A(n_3067),
.B(n_2278),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3110),
.A2(n_2284),
.B(n_2282),
.Y(n_3456)
);

NOR2xp67_ASAP7_75t_SL g3457 ( 
.A(n_3073),
.B(n_1918),
.Y(n_3457)
);

AOI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3034),
.A2(n_2284),
.B(n_2282),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3037),
.A2(n_2288),
.B(n_1745),
.Y(n_3459)
);

NOR2xp33_ASAP7_75t_L g3460 ( 
.A(n_3044),
.B(n_802),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3044),
.B(n_1568),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3257),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3251),
.B(n_3053),
.Y(n_3463)
);

INVx4_ASAP7_75t_L g3464 ( 
.A(n_3331),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3276),
.B(n_3246),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_L g3466 ( 
.A1(n_3430),
.A2(n_3149),
.B(n_3210),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3295),
.Y(n_3467)
);

AND2x2_ASAP7_75t_SL g3468 ( 
.A(n_3306),
.B(n_936),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_3267),
.B(n_3160),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3322),
.B(n_3167),
.Y(n_3470)
);

OAI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3343),
.A2(n_3120),
.B(n_3145),
.Y(n_3471)
);

AND2x2_ASAP7_75t_SL g3472 ( 
.A(n_3319),
.B(n_936),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3253),
.B(n_3168),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3312),
.B(n_1325),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3279),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3255),
.B(n_1326),
.Y(n_3476)
);

NAND4xp25_ASAP7_75t_L g3477 ( 
.A(n_3326),
.B(n_1317),
.C(n_1320),
.D(n_1316),
.Y(n_3477)
);

AOI21x1_ASAP7_75t_L g3478 ( 
.A1(n_3387),
.A2(n_3238),
.B(n_3227),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3316),
.B(n_804),
.Y(n_3479)
);

OA22x2_ASAP7_75t_L g3480 ( 
.A1(n_3254),
.A2(n_808),
.B1(n_809),
.B2(n_805),
.Y(n_3480)
);

NAND3xp33_ASAP7_75t_L g3481 ( 
.A(n_3460),
.B(n_3252),
.C(n_3356),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3432),
.Y(n_3482)
);

OAI21x1_ASAP7_75t_SL g3483 ( 
.A1(n_3435),
.A2(n_3137),
.B(n_3131),
.Y(n_3483)
);

INVxp67_ASAP7_75t_L g3484 ( 
.A(n_3351),
.Y(n_3484)
);

OAI21x1_ASAP7_75t_L g3485 ( 
.A1(n_3438),
.A2(n_3174),
.B(n_3151),
.Y(n_3485)
);

OAI21x1_ASAP7_75t_L g3486 ( 
.A1(n_3371),
.A2(n_3032),
.B(n_3224),
.Y(n_3486)
);

OAI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3304),
.A2(n_3184),
.B(n_3195),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3263),
.B(n_811),
.Y(n_3488)
);

AO31x2_ASAP7_75t_L g3489 ( 
.A1(n_3338),
.A2(n_3226),
.A3(n_3193),
.B(n_3185),
.Y(n_3489)
);

OA22x2_ASAP7_75t_L g3490 ( 
.A1(n_3274),
.A2(n_818),
.B1(n_821),
.B2(n_814),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_3283),
.Y(n_3491)
);

OAI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3332),
.A2(n_3199),
.B(n_3198),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3285),
.B(n_3202),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3311),
.A2(n_3054),
.B(n_3245),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3262),
.Y(n_3495)
);

AOI211x1_ASAP7_75t_L g3496 ( 
.A1(n_3362),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_3496)
);

OAI21x1_ASAP7_75t_L g3497 ( 
.A1(n_3258),
.A2(n_2178),
.B(n_2288),
.Y(n_3497)
);

CKINVDCx11_ASAP7_75t_R g3498 ( 
.A(n_3260),
.Y(n_3498)
);

INVx3_ASAP7_75t_L g3499 ( 
.A(n_3432),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3265),
.Y(n_3500)
);

AOI21x1_ASAP7_75t_SL g3501 ( 
.A1(n_3271),
.A2(n_3313),
.B(n_3287),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3259),
.B(n_823),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3296),
.A2(n_3272),
.B(n_3256),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3264),
.A2(n_1928),
.B(n_1745),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3281),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3329),
.B(n_830),
.Y(n_3506)
);

A2O1A1Ixp33_ASAP7_75t_L g3507 ( 
.A1(n_3335),
.A2(n_832),
.B(n_833),
.C(n_831),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3270),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3426),
.B(n_835),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3310),
.B(n_836),
.Y(n_3510)
);

BUFx12f_ASAP7_75t_L g3511 ( 
.A(n_3269),
.Y(n_3511)
);

OAI22xp5_ASAP7_75t_L g3512 ( 
.A1(n_3261),
.A2(n_890),
.B1(n_903),
.B2(n_854),
.Y(n_3512)
);

OAI21x1_ASAP7_75t_L g3513 ( 
.A1(n_3458),
.A2(n_1769),
.B(n_1742),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3442),
.A2(n_3418),
.B(n_3299),
.Y(n_3514)
);

OAI21x1_ASAP7_75t_L g3515 ( 
.A1(n_3459),
.A2(n_1769),
.B(n_1742),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3314),
.Y(n_3516)
);

AOI21xp33_ASAP7_75t_L g3517 ( 
.A1(n_3407),
.A2(n_1909),
.B(n_1902),
.Y(n_3517)
);

INVx1_ASAP7_75t_SL g3518 ( 
.A(n_3301),
.Y(n_3518)
);

AND2x4_ASAP7_75t_L g3519 ( 
.A(n_3379),
.B(n_1389),
.Y(n_3519)
);

NAND2x1p5_ASAP7_75t_L g3520 ( 
.A(n_3298),
.B(n_2173),
.Y(n_3520)
);

OAI21x1_ASAP7_75t_SL g3521 ( 
.A1(n_3294),
.A2(n_1772),
.B(n_1902),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_3301),
.Y(n_3522)
);

A2O1A1Ixp33_ASAP7_75t_SL g3523 ( 
.A1(n_3406),
.A2(n_1743),
.B(n_1780),
.C(n_1738),
.Y(n_3523)
);

AO31x2_ASAP7_75t_L g3524 ( 
.A1(n_3346),
.A2(n_1909),
.A3(n_1912),
.B(n_1911),
.Y(n_3524)
);

OAI21x1_ASAP7_75t_SL g3525 ( 
.A1(n_3282),
.A2(n_1772),
.B(n_1911),
.Y(n_3525)
);

BUFx2_ASAP7_75t_L g3526 ( 
.A(n_3354),
.Y(n_3526)
);

NAND2x1p5_ASAP7_75t_L g3527 ( 
.A(n_3298),
.B(n_2174),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3293),
.Y(n_3528)
);

AND2x4_ASAP7_75t_L g3529 ( 
.A(n_3379),
.B(n_1389),
.Y(n_3529)
);

O2A1O1Ixp5_ASAP7_75t_L g3530 ( 
.A1(n_3392),
.A2(n_1914),
.B(n_1919),
.C(n_1912),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3278),
.B(n_838),
.Y(n_3531)
);

AO31x2_ASAP7_75t_L g3532 ( 
.A1(n_3360),
.A2(n_1919),
.A3(n_1924),
.B(n_1914),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3388),
.A2(n_1704),
.B(n_1696),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_3367),
.B(n_3300),
.Y(n_3534)
);

BUFx12f_ASAP7_75t_L g3535 ( 
.A(n_3301),
.Y(n_3535)
);

OR2x6_ASAP7_75t_L g3536 ( 
.A(n_3266),
.B(n_2176),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3378),
.B(n_7),
.Y(n_3537)
);

INVx4_ASAP7_75t_L g3538 ( 
.A(n_3359),
.Y(n_3538)
);

AO31x2_ASAP7_75t_L g3539 ( 
.A1(n_3364),
.A2(n_3327),
.A3(n_3424),
.B(n_3411),
.Y(n_3539)
);

AOI21x1_ASAP7_75t_L g3540 ( 
.A1(n_3321),
.A2(n_1593),
.B(n_1568),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3453),
.B(n_839),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3268),
.A2(n_1704),
.B(n_1696),
.Y(n_3542)
);

AOI21xp5_ASAP7_75t_L g3543 ( 
.A1(n_3275),
.A2(n_1704),
.B(n_1696),
.Y(n_3543)
);

INVxp67_ASAP7_75t_SL g3544 ( 
.A(n_3449),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3307),
.Y(n_3545)
);

OAI21x1_ASAP7_75t_L g3546 ( 
.A1(n_3323),
.A2(n_1934),
.B(n_1924),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3320),
.Y(n_3547)
);

AOI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3403),
.A2(n_1593),
.B(n_1568),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3337),
.B(n_842),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3345),
.Y(n_3550)
);

OAI21xp33_ASAP7_75t_L g3551 ( 
.A1(n_3400),
.A2(n_852),
.B(n_851),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3447),
.A2(n_1712),
.B(n_1704),
.Y(n_3552)
);

BUFx3_ASAP7_75t_L g3553 ( 
.A(n_3273),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3291),
.B(n_855),
.Y(n_3554)
);

BUFx2_ASAP7_75t_SL g3555 ( 
.A(n_3288),
.Y(n_3555)
);

OAI21x1_ASAP7_75t_L g3556 ( 
.A1(n_3384),
.A2(n_1936),
.B(n_1934),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3334),
.Y(n_3557)
);

OAI21x1_ASAP7_75t_SL g3558 ( 
.A1(n_3372),
.A2(n_3339),
.B(n_3302),
.Y(n_3558)
);

BUFx6f_ASAP7_75t_L g3559 ( 
.A(n_3305),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3357),
.B(n_8),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3340),
.A2(n_1712),
.B(n_1704),
.Y(n_3561)
);

A2O1A1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_3297),
.A2(n_858),
.B(n_859),
.C(n_856),
.Y(n_3562)
);

OAI21x1_ASAP7_75t_L g3563 ( 
.A1(n_3416),
.A2(n_1937),
.B(n_1936),
.Y(n_3563)
);

OAI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3289),
.A2(n_3292),
.B1(n_3277),
.B2(n_3303),
.Y(n_3564)
);

OAI21x1_ASAP7_75t_L g3565 ( 
.A1(n_3451),
.A2(n_1949),
.B(n_1937),
.Y(n_3565)
);

AO31x2_ASAP7_75t_L g3566 ( 
.A1(n_3374),
.A2(n_1957),
.A3(n_1958),
.B(n_1949),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3394),
.Y(n_3567)
);

OAI21xp33_ASAP7_75t_L g3568 ( 
.A1(n_3439),
.A2(n_868),
.B(n_863),
.Y(n_3568)
);

OA22x2_ASAP7_75t_L g3569 ( 
.A1(n_3363),
.A2(n_877),
.B1(n_882),
.B2(n_875),
.Y(n_3569)
);

O2A1O1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_3330),
.A2(n_1593),
.B(n_1643),
.C(n_1599),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_3318),
.B(n_1389),
.Y(n_3571)
);

AND2x2_ASAP7_75t_SL g3572 ( 
.A(n_3379),
.B(n_936),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3445),
.B(n_887),
.Y(n_3573)
);

NOR4xp25_ASAP7_75t_L g3574 ( 
.A(n_3440),
.B(n_12),
.C(n_10),
.D(n_11),
.Y(n_3574)
);

AOI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_3325),
.A2(n_3290),
.B1(n_3317),
.B2(n_3280),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3428),
.A2(n_1716),
.B(n_1712),
.Y(n_3576)
);

OAI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_3441),
.A2(n_893),
.B1(n_894),
.B2(n_888),
.Y(n_3577)
);

AOI21x1_ASAP7_75t_L g3578 ( 
.A1(n_3452),
.A2(n_1643),
.B(n_1599),
.Y(n_3578)
);

AND2x2_ASAP7_75t_SL g3579 ( 
.A(n_3373),
.B(n_1599),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3398),
.B(n_1389),
.Y(n_3580)
);

AO31x2_ASAP7_75t_L g3581 ( 
.A1(n_3409),
.A2(n_1958),
.A3(n_1969),
.B(n_1957),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3443),
.A2(n_1716),
.B(n_1712),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3376),
.A2(n_1716),
.B(n_1712),
.Y(n_3583)
);

OAI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3385),
.A2(n_1507),
.B(n_1643),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3358),
.B(n_12),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3395),
.A2(n_3454),
.B(n_3452),
.Y(n_3586)
);

AO22x2_ASAP7_75t_L g3587 ( 
.A1(n_3377),
.A2(n_2180),
.B1(n_2183),
.B2(n_2176),
.Y(n_3587)
);

AO31x2_ASAP7_75t_L g3588 ( 
.A1(n_3444),
.A2(n_1985),
.A3(n_1987),
.B(n_1969),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3397),
.A2(n_3456),
.B(n_3421),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3361),
.Y(n_3590)
);

BUFx12f_ASAP7_75t_L g3591 ( 
.A(n_3284),
.Y(n_3591)
);

CKINVDCx6p67_ASAP7_75t_R g3592 ( 
.A(n_3284),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3445),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3369),
.Y(n_3594)
);

OR2x2_ASAP7_75t_L g3595 ( 
.A(n_3370),
.B(n_3383),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3436),
.B(n_3386),
.Y(n_3596)
);

NAND2x1_ASAP7_75t_L g3597 ( 
.A(n_3391),
.B(n_1400),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3381),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3423),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3412),
.A2(n_1987),
.B(n_1985),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3399),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3415),
.A2(n_900),
.B1(n_901),
.B2(n_897),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3365),
.B(n_905),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3349),
.B(n_1400),
.Y(n_3604)
);

CKINVDCx5p33_ASAP7_75t_R g3605 ( 
.A(n_3410),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3342),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3347),
.A2(n_1995),
.B(n_1994),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_3448),
.A2(n_909),
.B(n_910),
.C(n_908),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3348),
.A2(n_1995),
.B(n_1994),
.Y(n_3609)
);

OAI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3433),
.A2(n_914),
.B1(n_915),
.B2(n_911),
.Y(n_3610)
);

OAI21x1_ASAP7_75t_L g3611 ( 
.A1(n_3350),
.A2(n_1999),
.B(n_1998),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3352),
.A2(n_3446),
.B(n_3391),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3349),
.B(n_1400),
.Y(n_3613)
);

OAI21x1_ASAP7_75t_SL g3614 ( 
.A1(n_3422),
.A2(n_1999),
.B(n_1998),
.Y(n_3614)
);

OAI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3324),
.A2(n_917),
.B(n_916),
.Y(n_3615)
);

AOI221x1_ASAP7_75t_L g3616 ( 
.A1(n_3328),
.A2(n_1402),
.B1(n_1400),
.B2(n_1350),
.C(n_1357),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_3349),
.Y(n_3617)
);

AO31x2_ASAP7_75t_L g3618 ( 
.A1(n_3408),
.A2(n_2183),
.A3(n_2180),
.B(n_1371),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3429),
.Y(n_3619)
);

OAI21x1_ASAP7_75t_L g3620 ( 
.A1(n_3461),
.A2(n_1743),
.B(n_1738),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3366),
.A2(n_1780),
.B(n_1743),
.Y(n_3621)
);

A2O1A1Ixp33_ASAP7_75t_L g3622 ( 
.A1(n_3417),
.A2(n_3353),
.B(n_3344),
.C(n_3380),
.Y(n_3622)
);

NAND3x1_ASAP7_75t_L g3623 ( 
.A(n_3375),
.B(n_14),
.C(n_15),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3402),
.A2(n_3405),
.B(n_3404),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3333),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3404),
.A2(n_1780),
.B(n_1402),
.Y(n_3626)
);

NAND3xp33_ASAP7_75t_SL g3627 ( 
.A(n_3413),
.B(n_923),
.C(n_919),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3431),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_3286),
.A2(n_1734),
.B(n_1716),
.Y(n_3629)
);

O2A1O1Ixp5_ASAP7_75t_L g3630 ( 
.A1(n_3457),
.A2(n_1371),
.B(n_17),
.C(n_14),
.Y(n_3630)
);

BUFx2_ASAP7_75t_L g3631 ( 
.A(n_3389),
.Y(n_3631)
);

AOI211x1_ASAP7_75t_L g3632 ( 
.A1(n_3341),
.A2(n_19),
.B(n_16),
.C(n_18),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_SL g3633 ( 
.A(n_3437),
.B(n_1402),
.Y(n_3633)
);

AOI31xp67_ASAP7_75t_L g3634 ( 
.A1(n_3396),
.A2(n_1371),
.A3(n_1807),
.B(n_1800),
.Y(n_3634)
);

AOI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_3317),
.A2(n_926),
.B1(n_928),
.B2(n_925),
.Y(n_3635)
);

INVx4_ASAP7_75t_L g3636 ( 
.A(n_3375),
.Y(n_3636)
);

OAI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_3425),
.A2(n_933),
.B1(n_938),
.B2(n_931),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3365),
.B(n_945),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3309),
.A2(n_1734),
.B(n_1716),
.Y(n_3639)
);

INVx3_ASAP7_75t_SL g3640 ( 
.A(n_3315),
.Y(n_3640)
);

INVx1_ASAP7_75t_SL g3641 ( 
.A(n_3315),
.Y(n_3641)
);

INVx1_ASAP7_75t_SL g3642 ( 
.A(n_3305),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3333),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3333),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_L g3645 ( 
.A1(n_3455),
.A2(n_1402),
.B(n_1800),
.Y(n_3645)
);

OAI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3393),
.A2(n_1807),
.B(n_1800),
.Y(n_3646)
);

AO31x2_ASAP7_75t_L g3647 ( 
.A1(n_3427),
.A2(n_1371),
.A3(n_1808),
.B(n_1807),
.Y(n_3647)
);

OAI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3390),
.A2(n_949),
.B1(n_950),
.B2(n_947),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3305),
.B(n_18),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_SL g3650 ( 
.A1(n_3450),
.A2(n_20),
.B(n_21),
.Y(n_3650)
);

BUFx2_ASAP7_75t_SL g3651 ( 
.A(n_3308),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3434),
.B(n_951),
.Y(n_3652)
);

BUFx6f_ASAP7_75t_L g3653 ( 
.A(n_3308),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_3368),
.A2(n_1371),
.B1(n_1462),
.B2(n_1443),
.Y(n_3654)
);

AOI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3401),
.A2(n_954),
.B1(n_957),
.B2(n_953),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3373),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3309),
.A2(n_1744),
.B(n_1734),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3437),
.A2(n_1744),
.B(n_1734),
.Y(n_3658)
);

HB1xp67_ASAP7_75t_L g3659 ( 
.A(n_3382),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3419),
.A2(n_963),
.B(n_962),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3382),
.A2(n_1744),
.B(n_1734),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3336),
.A2(n_1751),
.B(n_1744),
.Y(n_3662)
);

AOI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_3420),
.A2(n_1751),
.B(n_1744),
.Y(n_3663)
);

OAI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_3355),
.A2(n_967),
.B(n_964),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_3308),
.A2(n_3414),
.B(n_1760),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3267),
.B(n_1512),
.Y(n_3666)
);

OAI22xp5_ASAP7_75t_SL g3667 ( 
.A1(n_3306),
.A2(n_973),
.B1(n_25),
.B2(n_21),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_SL g3668 ( 
.A1(n_3252),
.A2(n_22),
.B(n_27),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3276),
.B(n_22),
.Y(n_3669)
);

INVx4_ASAP7_75t_L g3670 ( 
.A(n_3331),
.Y(n_3670)
);

NAND2x1_ASAP7_75t_L g3671 ( 
.A(n_3391),
.B(n_1371),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3304),
.A2(n_1760),
.B(n_1751),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3276),
.B(n_28),
.Y(n_3673)
);

AO21x2_ASAP7_75t_L g3674 ( 
.A1(n_3430),
.A2(n_1524),
.B(n_1512),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3257),
.Y(n_3675)
);

OAI21xp5_ASAP7_75t_SL g3676 ( 
.A1(n_3267),
.A2(n_29),
.B(n_31),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_SL g3677 ( 
.A1(n_3252),
.A2(n_31),
.B(n_32),
.Y(n_3677)
);

OAI21xp33_ASAP7_75t_SL g3678 ( 
.A1(n_3460),
.A2(n_33),
.B(n_34),
.Y(n_3678)
);

A2O1A1Ixp33_ASAP7_75t_L g3679 ( 
.A1(n_3267),
.A2(n_751),
.B(n_754),
.C(n_749),
.Y(n_3679)
);

BUFx3_ASAP7_75t_L g3680 ( 
.A(n_3491),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3481),
.A2(n_1443),
.B1(n_1462),
.B2(n_1807),
.Y(n_3681)
);

OR2x6_ASAP7_75t_L g3682 ( 
.A(n_3555),
.B(n_1807),
.Y(n_3682)
);

OA21x2_ASAP7_75t_L g3683 ( 
.A1(n_3625),
.A2(n_769),
.B(n_765),
.Y(n_3683)
);

INVxp67_ASAP7_75t_L g3684 ( 
.A(n_3467),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3462),
.Y(n_3685)
);

NAND2xp33_ASAP7_75t_L g3686 ( 
.A(n_3667),
.B(n_3679),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3598),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3484),
.B(n_33),
.Y(n_3688)
);

OR2x2_ASAP7_75t_L g3689 ( 
.A(n_3544),
.B(n_3462),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3495),
.Y(n_3690)
);

AND2x4_ASAP7_75t_L g3691 ( 
.A(n_3482),
.B(n_34),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3495),
.Y(n_3692)
);

AND2x4_ASAP7_75t_L g3693 ( 
.A(n_3482),
.B(n_36),
.Y(n_3693)
);

NAND2x1p5_ASAP7_75t_L g3694 ( 
.A(n_3572),
.B(n_1808),
.Y(n_3694)
);

OAI321xp33_ASAP7_75t_L g3695 ( 
.A1(n_3615),
.A2(n_1989),
.A3(n_1823),
.B1(n_1808),
.B2(n_1829),
.C(n_1827),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3463),
.B(n_3593),
.Y(n_3696)
);

O2A1O1Ixp33_ASAP7_75t_L g3697 ( 
.A1(n_3676),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_3697)
);

BUFx2_ASAP7_75t_L g3698 ( 
.A(n_3631),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3465),
.B(n_37),
.Y(n_3699)
);

AND2x6_ASAP7_75t_L g3700 ( 
.A(n_3499),
.B(n_1808),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_3498),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_L g3702 ( 
.A1(n_3468),
.A2(n_1443),
.B1(n_1462),
.B2(n_1808),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3500),
.Y(n_3703)
);

INVx3_ASAP7_75t_L g3704 ( 
.A(n_3499),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3605),
.B(n_39),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3473),
.B(n_40),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3599),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3514),
.A2(n_1760),
.B(n_1751),
.Y(n_3708)
);

A2O1A1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3507),
.A2(n_3678),
.B(n_3575),
.C(n_3551),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3500),
.Y(n_3710)
);

BUFx2_ASAP7_75t_L g3711 ( 
.A(n_3535),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3475),
.Y(n_3712)
);

BUFx2_ASAP7_75t_L g3713 ( 
.A(n_3522),
.Y(n_3713)
);

OA21x2_ASAP7_75t_L g3714 ( 
.A1(n_3625),
.A2(n_3644),
.B(n_3643),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3508),
.B(n_41),
.Y(n_3715)
);

OAI21xp33_ASAP7_75t_L g3716 ( 
.A1(n_3469),
.A2(n_777),
.B(n_775),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3505),
.Y(n_3717)
);

AND2x6_ASAP7_75t_L g3718 ( 
.A(n_3656),
.B(n_1810),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_3553),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3503),
.A2(n_1760),
.B(n_1751),
.Y(n_3720)
);

CKINVDCx5p33_ASAP7_75t_R g3721 ( 
.A(n_3511),
.Y(n_3721)
);

HB1xp67_ASAP7_75t_L g3722 ( 
.A(n_3508),
.Y(n_3722)
);

BUFx3_ASAP7_75t_L g3723 ( 
.A(n_3591),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3528),
.Y(n_3724)
);

OR2x6_ASAP7_75t_L g3725 ( 
.A(n_3651),
.B(n_1810),
.Y(n_3725)
);

A2O1A1Ixp33_ASAP7_75t_L g3726 ( 
.A1(n_3568),
.A2(n_783),
.B(n_787),
.C(n_782),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3669),
.B(n_41),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3516),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3528),
.Y(n_3729)
);

OR2x2_ASAP7_75t_SL g3730 ( 
.A(n_3619),
.B(n_42),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3675),
.B(n_42),
.Y(n_3731)
);

INVx1_ASAP7_75t_SL g3732 ( 
.A(n_3518),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3673),
.B(n_43),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3534),
.B(n_44),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3640),
.B(n_44),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3472),
.B(n_902),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_SL g3737 ( 
.A1(n_3564),
.A2(n_902),
.B1(n_791),
.B2(n_799),
.Y(n_3737)
);

BUFx2_ASAP7_75t_L g3738 ( 
.A(n_3636),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3595),
.B(n_45),
.Y(n_3739)
);

O2A1O1Ixp5_ASAP7_75t_SL g3740 ( 
.A1(n_3493),
.A2(n_3666),
.B(n_3644),
.C(n_3643),
.Y(n_3740)
);

INVx2_ASAP7_75t_SL g3741 ( 
.A(n_3592),
.Y(n_3741)
);

AOI22xp33_ASAP7_75t_L g3742 ( 
.A1(n_3480),
.A2(n_3490),
.B1(n_3557),
.B2(n_3628),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3675),
.B(n_3470),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3494),
.A2(n_1761),
.B(n_1760),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3567),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3526),
.B(n_3590),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3545),
.B(n_45),
.Y(n_3747)
);

HB1xp67_ASAP7_75t_L g3748 ( 
.A(n_3547),
.Y(n_3748)
);

INVx3_ASAP7_75t_L g3749 ( 
.A(n_3636),
.Y(n_3749)
);

INVx3_ASAP7_75t_L g3750 ( 
.A(n_3550),
.Y(n_3750)
);

NAND2x1p5_ASAP7_75t_L g3751 ( 
.A(n_3464),
.B(n_1810),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3596),
.B(n_46),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3594),
.B(n_46),
.Y(n_3753)
);

AOI22xp33_ASAP7_75t_L g3754 ( 
.A1(n_3569),
.A2(n_1443),
.B1(n_1462),
.B2(n_1810),
.Y(n_3754)
);

CKINVDCx6p67_ASAP7_75t_R g3755 ( 
.A(n_3464),
.Y(n_3755)
);

CKINVDCx20_ASAP7_75t_R g3756 ( 
.A(n_3538),
.Y(n_3756)
);

INVx4_ASAP7_75t_L g3757 ( 
.A(n_3538),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3601),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3656),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3587),
.Y(n_3760)
);

A2O1A1Ixp33_ASAP7_75t_SL g3761 ( 
.A1(n_3664),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_3761)
);

INVx4_ASAP7_75t_L g3762 ( 
.A(n_3670),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3606),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_3552),
.A2(n_1768),
.B(n_1761),
.Y(n_3764)
);

BUFx2_ASAP7_75t_L g3765 ( 
.A(n_3670),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3487),
.A2(n_1768),
.B(n_1761),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3606),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3672),
.A2(n_1768),
.B(n_1761),
.Y(n_3768)
);

INVx1_ASAP7_75t_SL g3769 ( 
.A(n_3537),
.Y(n_3769)
);

CKINVDCx5p33_ASAP7_75t_R g3770 ( 
.A(n_3559),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3512),
.A2(n_902),
.B1(n_1823),
.B2(n_1810),
.Y(n_3771)
);

INVx2_ASAP7_75t_SL g3772 ( 
.A(n_3559),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3659),
.B(n_47),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3623),
.A2(n_810),
.B1(n_816),
.B2(n_788),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3582),
.A2(n_1768),
.B(n_1761),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3539),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3539),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3558),
.A2(n_1768),
.B(n_1823),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3589),
.A2(n_1827),
.B(n_1823),
.Y(n_3779)
);

INVx3_ASAP7_75t_L g3780 ( 
.A(n_3559),
.Y(n_3780)
);

O2A1O1Ixp33_ASAP7_75t_L g3781 ( 
.A1(n_3562),
.A2(n_51),
.B(n_48),
.C(n_50),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3492),
.A2(n_1827),
.B(n_1823),
.Y(n_3782)
);

OAI21x1_ASAP7_75t_SL g3783 ( 
.A1(n_3650),
.A2(n_50),
.B(n_52),
.Y(n_3783)
);

AND2x4_ASAP7_75t_L g3784 ( 
.A(n_3641),
.B(n_52),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3474),
.B(n_53),
.Y(n_3785)
);

INVx3_ASAP7_75t_L g3786 ( 
.A(n_3653),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3587),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3560),
.B(n_54),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3585),
.B(n_56),
.Y(n_3789)
);

AOI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_3586),
.A2(n_1829),
.B(n_1827),
.Y(n_3790)
);

AOI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3571),
.A2(n_3627),
.B1(n_3579),
.B2(n_3536),
.Y(n_3791)
);

AOI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3597),
.A2(n_902),
.B(n_845),
.Y(n_3792)
);

AOI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3540),
.A2(n_902),
.B(n_869),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3476),
.Y(n_3794)
);

O2A1O1Ixp33_ASAP7_75t_SL g3795 ( 
.A1(n_3608),
.A2(n_64),
.B(n_56),
.C(n_57),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3539),
.Y(n_3796)
);

AOI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3542),
.A2(n_1829),
.B(n_1827),
.Y(n_3797)
);

OA21x2_ASAP7_75t_L g3798 ( 
.A1(n_3624),
.A2(n_870),
.B(n_825),
.Y(n_3798)
);

BUFx3_ASAP7_75t_L g3799 ( 
.A(n_3653),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3581),
.Y(n_3800)
);

BUFx6f_ASAP7_75t_L g3801 ( 
.A(n_3653),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3617),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3543),
.A2(n_1845),
.B(n_1829),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3554),
.B(n_57),
.Y(n_3804)
);

INVx1_ASAP7_75t_SL g3805 ( 
.A(n_3642),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3581),
.Y(n_3806)
);

AND2x4_ASAP7_75t_L g3807 ( 
.A(n_3580),
.B(n_64),
.Y(n_3807)
);

BUFx3_ASAP7_75t_L g3808 ( 
.A(n_3649),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_3479),
.B(n_65),
.Y(n_3809)
);

BUFx6f_ASAP7_75t_L g3810 ( 
.A(n_3536),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3581),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3496),
.A2(n_884),
.B1(n_896),
.B2(n_879),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3566),
.Y(n_3813)
);

INVx3_ASAP7_75t_L g3814 ( 
.A(n_3485),
.Y(n_3814)
);

BUFx6f_ASAP7_75t_L g3815 ( 
.A(n_3520),
.Y(n_3815)
);

OAI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3632),
.A2(n_3622),
.B1(n_3635),
.B2(n_3655),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3612),
.Y(n_3817)
);

BUFx6f_ASAP7_75t_L g3818 ( 
.A(n_3527),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3566),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3566),
.Y(n_3820)
);

AOI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3483),
.A2(n_1845),
.B(n_1829),
.Y(n_3821)
);

OR2x6_ASAP7_75t_L g3822 ( 
.A(n_3658),
.B(n_1845),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3488),
.B(n_65),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3502),
.B(n_66),
.Y(n_3824)
);

OAI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3573),
.A2(n_937),
.B1(n_942),
.B2(n_924),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3588),
.Y(n_3826)
);

NAND2x1p5_ASAP7_75t_L g3827 ( 
.A(n_3633),
.B(n_1845),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3531),
.B(n_66),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3524),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_3652),
.Y(n_3830)
);

INVx4_ASAP7_75t_SL g3831 ( 
.A(n_3580),
.Y(n_3831)
);

OAI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3574),
.A2(n_955),
.B(n_946),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3506),
.B(n_67),
.Y(n_3833)
);

OR2x2_ASAP7_75t_L g3834 ( 
.A(n_3509),
.B(n_67),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_SL g3835 ( 
.A(n_3519),
.B(n_902),
.Y(n_3835)
);

AOI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3610),
.A2(n_902),
.B1(n_1848),
.B2(n_1845),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3510),
.B(n_68),
.Y(n_3837)
);

AOI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3602),
.A2(n_3584),
.B1(n_3477),
.B2(n_3637),
.Y(n_3838)
);

BUFx4_ASAP7_75t_SL g3839 ( 
.A(n_3501),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3523),
.A2(n_1871),
.B(n_1848),
.Y(n_3840)
);

BUFx6f_ASAP7_75t_L g3841 ( 
.A(n_3519),
.Y(n_3841)
);

A2O1A1Ixp33_ASAP7_75t_SL g3842 ( 
.A1(n_3660),
.A2(n_71),
.B(n_68),
.C(n_69),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_3603),
.B(n_72),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3588),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3638),
.A2(n_3577),
.B1(n_3648),
.B2(n_3541),
.Y(n_3845)
);

INVx1_ASAP7_75t_SL g3846 ( 
.A(n_3549),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3588),
.Y(n_3847)
);

BUFx3_ASAP7_75t_L g3848 ( 
.A(n_3529),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3533),
.A2(n_1871),
.B(n_1848),
.Y(n_3849)
);

CKINVDCx11_ASAP7_75t_R g3850 ( 
.A(n_3529),
.Y(n_3850)
);

BUFx3_ASAP7_75t_L g3851 ( 
.A(n_3671),
.Y(n_3851)
);

BUFx2_ASAP7_75t_L g3852 ( 
.A(n_3647),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3524),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3524),
.Y(n_3854)
);

AND2x4_ASAP7_75t_L g3855 ( 
.A(n_3471),
.B(n_3665),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3626),
.Y(n_3856)
);

OR2x2_ASAP7_75t_SL g3857 ( 
.A(n_3668),
.B(n_72),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3621),
.B(n_3661),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3489),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3532),
.B(n_73),
.Y(n_3860)
);

BUFx2_ASAP7_75t_L g3861 ( 
.A(n_3647),
.Y(n_3861)
);

NAND3xp33_ASAP7_75t_L g3862 ( 
.A(n_3630),
.B(n_1547),
.C(n_1544),
.Y(n_3862)
);

INVx3_ASAP7_75t_L g3863 ( 
.A(n_3647),
.Y(n_3863)
);

BUFx12f_ASAP7_75t_L g3864 ( 
.A(n_3677),
.Y(n_3864)
);

BUFx6f_ASAP7_75t_L g3865 ( 
.A(n_3646),
.Y(n_3865)
);

OR2x2_ASAP7_75t_L g3866 ( 
.A(n_3532),
.B(n_3489),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3478),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3532),
.B(n_73),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3604),
.Y(n_3869)
);

O2A1O1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_3525),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_3870)
);

INVx4_ASAP7_75t_L g3871 ( 
.A(n_3674),
.Y(n_3871)
);

CKINVDCx16_ASAP7_75t_R g3872 ( 
.A(n_3613),
.Y(n_3872)
);

NOR2xp67_ASAP7_75t_SL g3873 ( 
.A(n_3629),
.B(n_1989),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3489),
.B(n_74),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3654),
.A2(n_966),
.B1(n_974),
.B2(n_958),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3620),
.B(n_77),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3517),
.A2(n_3614),
.B1(n_3663),
.B2(n_3662),
.Y(n_3877)
);

HB1xp67_ASAP7_75t_L g3878 ( 
.A(n_3618),
.Y(n_3878)
);

HB1xp67_ASAP7_75t_L g3879 ( 
.A(n_3618),
.Y(n_3879)
);

BUFx3_ASAP7_75t_L g3880 ( 
.A(n_3521),
.Y(n_3880)
);

BUFx2_ASAP7_75t_L g3881 ( 
.A(n_3618),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3561),
.A2(n_1871),
.B(n_1848),
.Y(n_3882)
);

BUFx2_ASAP7_75t_L g3883 ( 
.A(n_3466),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3486),
.B(n_78),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3607),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3576),
.A2(n_1871),
.B(n_1848),
.Y(n_3886)
);

CKINVDCx20_ASAP7_75t_R g3887 ( 
.A(n_3639),
.Y(n_3887)
);

HB1xp67_ASAP7_75t_L g3888 ( 
.A(n_3609),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3611),
.Y(n_3889)
);

AOI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_3504),
.A2(n_1877),
.B(n_1871),
.Y(n_3890)
);

CKINVDCx5p33_ASAP7_75t_R g3891 ( 
.A(n_3657),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3583),
.A2(n_1888),
.B(n_1877),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3570),
.A2(n_1547),
.B(n_1554),
.C(n_1544),
.Y(n_3893)
);

AND2x6_ASAP7_75t_L g3894 ( 
.A(n_3530),
.B(n_1877),
.Y(n_3894)
);

HB1xp67_ASAP7_75t_L g3895 ( 
.A(n_3600),
.Y(n_3895)
);

INVx3_ASAP7_75t_SL g3896 ( 
.A(n_3634),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3616),
.A2(n_1888),
.B(n_1877),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3497),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3548),
.B(n_79),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3546),
.B(n_79),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3556),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3515),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3645),
.B(n_80),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3687),
.Y(n_3904)
);

BUFx4f_ASAP7_75t_SL g3905 ( 
.A(n_3701),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3707),
.Y(n_3906)
);

AOI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3686),
.A2(n_902),
.B1(n_3563),
.B2(n_1553),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_SL g3908 ( 
.A1(n_3683),
.A2(n_3513),
.B1(n_3565),
.B2(n_1547),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3680),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3838),
.A2(n_3578),
.B1(n_85),
.B2(n_82),
.Y(n_3910)
);

OAI22xp5_ASAP7_75t_SL g3911 ( 
.A1(n_3730),
.A2(n_86),
.B1(n_82),
.B2(n_84),
.Y(n_3911)
);

CKINVDCx11_ASAP7_75t_R g3912 ( 
.A(n_3756),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3816),
.A2(n_1462),
.B1(n_1443),
.B2(n_1877),
.Y(n_3913)
);

CKINVDCx5p33_ASAP7_75t_R g3914 ( 
.A(n_3719),
.Y(n_3914)
);

INVx4_ASAP7_75t_L g3915 ( 
.A(n_3757),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3846),
.A2(n_1895),
.B1(n_1939),
.B2(n_1888),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3696),
.B(n_87),
.Y(n_3917)
);

BUFx4_ASAP7_75t_R g3918 ( 
.A(n_3723),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3759),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3697),
.A2(n_3857),
.B1(n_3709),
.B2(n_3699),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3716),
.A2(n_1895),
.B1(n_1939),
.B2(n_1888),
.Y(n_3921)
);

CKINVDCx5p33_ASAP7_75t_R g3922 ( 
.A(n_3721),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3767),
.Y(n_3923)
);

INVx6_ASAP7_75t_L g3924 ( 
.A(n_3757),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3704),
.Y(n_3925)
);

AOI22xp33_ASAP7_75t_L g3926 ( 
.A1(n_3809),
.A2(n_1895),
.B1(n_1939),
.B2(n_1888),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3722),
.Y(n_3927)
);

BUFx6f_ASAP7_75t_L g3928 ( 
.A(n_3850),
.Y(n_3928)
);

BUFx3_ASAP7_75t_L g3929 ( 
.A(n_3830),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3742),
.A2(n_1939),
.B1(n_1989),
.B2(n_1895),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3712),
.Y(n_3931)
);

INVx3_ASAP7_75t_SL g3932 ( 
.A(n_3755),
.Y(n_3932)
);

INVx6_ASAP7_75t_L g3933 ( 
.A(n_3762),
.Y(n_3933)
);

BUFx6f_ASAP7_75t_L g3934 ( 
.A(n_3801),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3748),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3685),
.Y(n_3936)
);

INVx8_ASAP7_75t_L g3937 ( 
.A(n_3682),
.Y(n_3937)
);

BUFx3_ASAP7_75t_L g3938 ( 
.A(n_3746),
.Y(n_3938)
);

INVx2_ASAP7_75t_SL g3939 ( 
.A(n_3713),
.Y(n_3939)
);

OAI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3706),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_3940)
);

INVx6_ASAP7_75t_L g3941 ( 
.A(n_3762),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_SL g3942 ( 
.A1(n_3683),
.A2(n_1547),
.B1(n_1554),
.B2(n_1544),
.Y(n_3942)
);

BUFx4f_ASAP7_75t_SL g3943 ( 
.A(n_3711),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3685),
.Y(n_3944)
);

BUFx6f_ASAP7_75t_L g3945 ( 
.A(n_3801),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3690),
.Y(n_3946)
);

INVx4_ASAP7_75t_L g3947 ( 
.A(n_3682),
.Y(n_3947)
);

OAI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3737),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3690),
.Y(n_3949)
);

OAI22xp5_ASAP7_75t_L g3950 ( 
.A1(n_3715),
.A2(n_3731),
.B1(n_3804),
.B2(n_3752),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3692),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3717),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3864),
.A2(n_1939),
.B1(n_1989),
.B2(n_1895),
.Y(n_3953)
);

INVx6_ASAP7_75t_L g3954 ( 
.A(n_3841),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_SL g3955 ( 
.A1(n_3734),
.A2(n_93),
.B(n_94),
.Y(n_3955)
);

AOI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3736),
.A2(n_1553),
.B1(n_1619),
.B2(n_1476),
.Y(n_3956)
);

CKINVDCx16_ASAP7_75t_R g3957 ( 
.A(n_3808),
.Y(n_3957)
);

INVx1_ASAP7_75t_SL g3958 ( 
.A(n_3698),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3760),
.A2(n_1989),
.B1(n_1512),
.B2(n_1530),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3787),
.A2(n_1512),
.B1(n_1530),
.B2(n_1524),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3692),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3743),
.B(n_93),
.Y(n_3962)
);

INVx1_ASAP7_75t_SL g3963 ( 
.A(n_3732),
.Y(n_3963)
);

BUFx4f_ASAP7_75t_SL g3964 ( 
.A(n_3741),
.Y(n_3964)
);

AOI22xp33_ASAP7_75t_L g3965 ( 
.A1(n_3832),
.A2(n_1512),
.B1(n_1530),
.B2(n_1524),
.Y(n_3965)
);

CKINVDCx14_ASAP7_75t_R g3966 ( 
.A(n_3705),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3791),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3728),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3794),
.A2(n_3843),
.B1(n_3868),
.B2(n_3860),
.Y(n_3969)
);

CKINVDCx11_ASAP7_75t_R g3970 ( 
.A(n_3769),
.Y(n_3970)
);

BUFx12f_ASAP7_75t_L g3971 ( 
.A(n_3834),
.Y(n_3971)
);

INVx5_ASAP7_75t_L g3972 ( 
.A(n_3700),
.Y(n_3972)
);

INVx6_ASAP7_75t_SL g3973 ( 
.A(n_3784),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3754),
.A2(n_1524),
.B1(n_1530),
.B2(n_1476),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_SL g3975 ( 
.A1(n_3798),
.A2(n_1547),
.B1(n_1554),
.B2(n_1544),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3684),
.B(n_95),
.Y(n_3976)
);

OAI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3872),
.A2(n_3845),
.B1(n_3874),
.B2(n_3887),
.Y(n_3977)
);

BUFx3_ASAP7_75t_L g3978 ( 
.A(n_3765),
.Y(n_3978)
);

INVx6_ASAP7_75t_L g3979 ( 
.A(n_3841),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3745),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3783),
.A2(n_1524),
.B1(n_1530),
.B2(n_1476),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3812),
.A2(n_1553),
.B1(n_1619),
.B2(n_1476),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3758),
.Y(n_3983)
);

INVxp67_ASAP7_75t_L g3984 ( 
.A(n_3802),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3710),
.Y(n_3985)
);

OAI22xp33_ASAP7_75t_L g3986 ( 
.A1(n_3739),
.A2(n_1554),
.B1(n_1557),
.B2(n_1544),
.Y(n_3986)
);

CKINVDCx6p67_ASAP7_75t_R g3987 ( 
.A(n_3735),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3710),
.Y(n_3988)
);

BUFx10_ASAP7_75t_L g3989 ( 
.A(n_3691),
.Y(n_3989)
);

CKINVDCx11_ASAP7_75t_R g3990 ( 
.A(n_3805),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3724),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3774),
.A2(n_1553),
.B1(n_1619),
.B2(n_1476),
.Y(n_3992)
);

INVx2_ASAP7_75t_SL g3993 ( 
.A(n_3770),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_3799),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3724),
.Y(n_3995)
);

INVx8_ASAP7_75t_L g3996 ( 
.A(n_3725),
.Y(n_3996)
);

BUFx8_ASAP7_75t_L g3997 ( 
.A(n_3788),
.Y(n_3997)
);

BUFx10_ASAP7_75t_L g3998 ( 
.A(n_3691),
.Y(n_3998)
);

CKINVDCx20_ASAP7_75t_R g3999 ( 
.A(n_3789),
.Y(n_3999)
);

OAI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3693),
.A2(n_3785),
.B1(n_3702),
.B2(n_3781),
.Y(n_4000)
);

BUFx2_ASAP7_75t_SL g4001 ( 
.A(n_3693),
.Y(n_4001)
);

OAI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3810),
.A2(n_1557),
.B1(n_1558),
.B2(n_1554),
.Y(n_4002)
);

BUFx2_ASAP7_75t_L g4003 ( 
.A(n_3738),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3729),
.Y(n_4004)
);

BUFx10_ASAP7_75t_L g4005 ( 
.A(n_3807),
.Y(n_4005)
);

BUFx3_ASAP7_75t_L g4006 ( 
.A(n_3784),
.Y(n_4006)
);

CKINVDCx20_ASAP7_75t_R g4007 ( 
.A(n_3727),
.Y(n_4007)
);

AOI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3798),
.A2(n_3823),
.B1(n_3824),
.B2(n_3828),
.Y(n_4008)
);

BUFx12f_ASAP7_75t_L g4009 ( 
.A(n_3733),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3837),
.A2(n_1619),
.B1(n_1553),
.B2(n_1558),
.Y(n_4010)
);

BUFx10_ASAP7_75t_L g4011 ( 
.A(n_3807),
.Y(n_4011)
);

OAI22xp5_ASAP7_75t_L g4012 ( 
.A1(n_3833),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_4012)
);

CKINVDCx11_ASAP7_75t_R g4013 ( 
.A(n_3801),
.Y(n_4013)
);

BUFx10_ASAP7_75t_L g4014 ( 
.A(n_3876),
.Y(n_4014)
);

AOI22xp33_ASAP7_75t_SL g4015 ( 
.A1(n_3776),
.A2(n_1557),
.B1(n_1564),
.B2(n_1558),
.Y(n_4015)
);

BUFx2_ASAP7_75t_L g4016 ( 
.A(n_3704),
.Y(n_4016)
);

BUFx2_ASAP7_75t_L g4017 ( 
.A(n_3749),
.Y(n_4017)
);

CKINVDCx6p67_ASAP7_75t_R g4018 ( 
.A(n_3688),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3796),
.A2(n_1619),
.B1(n_1553),
.B2(n_1558),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3763),
.Y(n_4020)
);

BUFx3_ASAP7_75t_L g4021 ( 
.A(n_3848),
.Y(n_4021)
);

INVx1_ASAP7_75t_SL g4022 ( 
.A(n_3689),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3729),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_3776),
.A2(n_1619),
.B1(n_1558),
.B2(n_1564),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3703),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3750),
.Y(n_4026)
);

INVx6_ASAP7_75t_L g4027 ( 
.A(n_3841),
.Y(n_4027)
);

BUFx2_ASAP7_75t_L g4028 ( 
.A(n_3749),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3750),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3747),
.A2(n_100),
.B1(n_97),
.B2(n_98),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3714),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3777),
.A2(n_1564),
.B1(n_1557),
.B2(n_1349),
.Y(n_4032)
);

OAI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3753),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_4033)
);

BUFx6f_ASAP7_75t_L g4034 ( 
.A(n_3810),
.Y(n_4034)
);

BUFx6f_ASAP7_75t_L g4035 ( 
.A(n_3810),
.Y(n_4035)
);

BUFx3_ASAP7_75t_L g4036 ( 
.A(n_3773),
.Y(n_4036)
);

OAI22x1_ASAP7_75t_L g4037 ( 
.A1(n_3839),
.A2(n_3714),
.B1(n_3817),
.B2(n_3891),
.Y(n_4037)
);

AOI21xp33_ASAP7_75t_SL g4038 ( 
.A1(n_3884),
.A2(n_101),
.B(n_102),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3777),
.Y(n_4039)
);

INVx3_ASAP7_75t_L g4040 ( 
.A(n_3780),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3867),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3859),
.Y(n_4042)
);

INVx3_ASAP7_75t_L g4043 ( 
.A(n_3780),
.Y(n_4043)
);

BUFx8_ASAP7_75t_L g4044 ( 
.A(n_3899),
.Y(n_4044)
);

INVx3_ASAP7_75t_SL g4045 ( 
.A(n_3772),
.Y(n_4045)
);

INVx2_ASAP7_75t_SL g4046 ( 
.A(n_3786),
.Y(n_4046)
);

BUFx2_ASAP7_75t_L g4047 ( 
.A(n_3786),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3813),
.Y(n_4048)
);

INVx6_ASAP7_75t_L g4049 ( 
.A(n_3831),
.Y(n_4049)
);

BUFx3_ASAP7_75t_L g4050 ( 
.A(n_3815),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3820),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3859),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_SL g4053 ( 
.A1(n_3852),
.A2(n_1564),
.B1(n_1557),
.B2(n_107),
.Y(n_4053)
);

BUFx4_ASAP7_75t_R g4054 ( 
.A(n_3851),
.Y(n_4054)
);

BUFx2_ASAP7_75t_L g4055 ( 
.A(n_3700),
.Y(n_4055)
);

AOI22xp33_ASAP7_75t_L g4056 ( 
.A1(n_3862),
.A2(n_1564),
.B1(n_1349),
.B2(n_1350),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3870),
.A2(n_111),
.B1(n_104),
.B2(n_105),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3819),
.Y(n_4058)
);

BUFx2_ASAP7_75t_L g4059 ( 
.A(n_3700),
.Y(n_4059)
);

BUFx3_ASAP7_75t_L g4060 ( 
.A(n_3815),
.Y(n_4060)
);

CKINVDCx11_ASAP7_75t_R g4061 ( 
.A(n_3831),
.Y(n_4061)
);

OAI22xp33_ASAP7_75t_L g4062 ( 
.A1(n_3695),
.A2(n_112),
.B1(n_105),
.B2(n_111),
.Y(n_4062)
);

AOI22xp33_ASAP7_75t_L g4063 ( 
.A1(n_3771),
.A2(n_1349),
.B1(n_1350),
.B2(n_1347),
.Y(n_4063)
);

BUFx2_ASAP7_75t_R g4064 ( 
.A(n_3835),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3861),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3836),
.A2(n_1349),
.B1(n_1350),
.B2(n_1347),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3866),
.Y(n_4067)
);

BUFx2_ASAP7_75t_SL g4068 ( 
.A(n_3700),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3869),
.B(n_112),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3782),
.A2(n_1357),
.B(n_1347),
.Y(n_4070)
);

INVx2_ASAP7_75t_SL g4071 ( 
.A(n_3815),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3876),
.A2(n_1357),
.B1(n_1359),
.B2(n_1347),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3895),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3881),
.A2(n_1359),
.B1(n_1360),
.B2(n_1357),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3811),
.Y(n_4075)
);

INVx1_ASAP7_75t_SL g4076 ( 
.A(n_3718),
.Y(n_4076)
);

CKINVDCx6p67_ASAP7_75t_R g4077 ( 
.A(n_3725),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3825),
.A2(n_1360),
.B1(n_1367),
.B2(n_1359),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3811),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_3681),
.A2(n_1360),
.B1(n_1367),
.B2(n_1359),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_4031),
.B(n_3740),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_SL g4082 ( 
.A1(n_4037),
.A2(n_3855),
.B(n_3880),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3977),
.A2(n_3766),
.B(n_3778),
.Y(n_4083)
);

HB1xp67_ASAP7_75t_L g4084 ( 
.A(n_3927),
.Y(n_4084)
);

OA22x2_ASAP7_75t_L g4085 ( 
.A1(n_3955),
.A2(n_3855),
.B1(n_3903),
.B2(n_3896),
.Y(n_4085)
);

AOI21xp5_ASAP7_75t_SL g4086 ( 
.A1(n_3920),
.A2(n_3900),
.B(n_3790),
.Y(n_4086)
);

OA21x2_ASAP7_75t_L g4087 ( 
.A1(n_4039),
.A2(n_3806),
.B(n_3800),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3936),
.Y(n_4088)
);

INVxp67_ASAP7_75t_L g4089 ( 
.A(n_4003),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_SL g4090 ( 
.A1(n_3920),
.A2(n_3708),
.B(n_3858),
.Y(n_4090)
);

OAI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_3955),
.A2(n_3877),
.B1(n_3694),
.B2(n_3744),
.Y(n_4091)
);

HB1xp67_ASAP7_75t_L g4092 ( 
.A(n_3923),
.Y(n_4092)
);

OA21x2_ASAP7_75t_L g4093 ( 
.A1(n_4042),
.A2(n_3883),
.B(n_3853),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_4022),
.B(n_3858),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3958),
.B(n_3814),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3958),
.B(n_3814),
.Y(n_4096)
);

O2A1O1Ixp33_ASAP7_75t_L g4097 ( 
.A1(n_3940),
.A2(n_3795),
.B(n_3842),
.C(n_3761),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3944),
.Y(n_4098)
);

NOR2x1_ASAP7_75t_SL g4099 ( 
.A(n_4068),
.B(n_4001),
.Y(n_4099)
);

OAI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_3969),
.A2(n_3726),
.B1(n_3751),
.B2(n_3822),
.Y(n_4100)
);

AND2x2_ASAP7_75t_L g4101 ( 
.A(n_3939),
.B(n_3888),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4022),
.B(n_3898),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3984),
.B(n_3898),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_4016),
.B(n_3901),
.Y(n_4104)
);

INVx5_ASAP7_75t_L g4105 ( 
.A(n_3928),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_4017),
.B(n_3889),
.Y(n_4106)
);

INVx3_ASAP7_75t_L g4107 ( 
.A(n_3925),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_3935),
.B(n_3854),
.Y(n_4108)
);

AND2x4_ASAP7_75t_L g4109 ( 
.A(n_4055),
.B(n_3863),
.Y(n_4109)
);

OA21x2_ASAP7_75t_L g4110 ( 
.A1(n_4052),
.A2(n_3853),
.B(n_3829),
.Y(n_4110)
);

INVx3_ASAP7_75t_L g4111 ( 
.A(n_3925),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3963),
.B(n_3889),
.Y(n_4112)
);

OR2x2_ASAP7_75t_L g4113 ( 
.A(n_3963),
.B(n_3829),
.Y(n_4113)
);

NOR2xp67_ASAP7_75t_L g4114 ( 
.A(n_3972),
.B(n_3863),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_4028),
.B(n_3878),
.Y(n_4115)
);

CKINVDCx20_ASAP7_75t_R g4116 ( 
.A(n_3905),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4026),
.B(n_3865),
.Y(n_4117)
);

INVxp67_ASAP7_75t_L g4118 ( 
.A(n_3929),
.Y(n_4118)
);

HB1xp67_ASAP7_75t_L g4119 ( 
.A(n_4029),
.Y(n_4119)
);

A2O1A1Ixp33_ASAP7_75t_L g4120 ( 
.A1(n_4008),
.A2(n_3893),
.B(n_3779),
.C(n_3879),
.Y(n_4120)
);

INVxp67_ASAP7_75t_SL g4121 ( 
.A(n_4065),
.Y(n_4121)
);

O2A1O1Ixp33_ASAP7_75t_L g4122 ( 
.A1(n_3940),
.A2(n_4038),
.B(n_4033),
.C(n_4012),
.Y(n_4122)
);

O2A1O1Ixp5_ASAP7_75t_L g4123 ( 
.A1(n_3917),
.A2(n_3871),
.B(n_3720),
.C(n_3764),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_3957),
.B(n_3978),
.Y(n_4124)
);

AOI21x1_ASAP7_75t_SL g4125 ( 
.A1(n_3962),
.A2(n_3873),
.B(n_3792),
.Y(n_4125)
);

NOR2xp67_ASAP7_75t_L g4126 ( 
.A(n_3972),
.B(n_3871),
.Y(n_4126)
);

NOR2xp67_ASAP7_75t_L g4127 ( 
.A(n_3972),
.B(n_3902),
.Y(n_4127)
);

HB1xp67_ASAP7_75t_L g4128 ( 
.A(n_4073),
.Y(n_4128)
);

O2A1O1Ixp5_ASAP7_75t_L g4129 ( 
.A1(n_3950),
.A2(n_3821),
.B(n_3775),
.C(n_3882),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_4020),
.B(n_3865),
.Y(n_4130)
);

AOI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_4062),
.A2(n_3822),
.B(n_3892),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3938),
.B(n_3902),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3946),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_4041),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_SL g4135 ( 
.A1(n_3928),
.A2(n_3818),
.B(n_3865),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3949),
.B(n_3718),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4036),
.B(n_4047),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3951),
.Y(n_4138)
);

OAI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_4038),
.A2(n_3818),
.B1(n_3827),
.B2(n_3768),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3961),
.Y(n_4140)
);

OA21x2_ASAP7_75t_L g4141 ( 
.A1(n_4075),
.A2(n_3844),
.B(n_3826),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_3987),
.B(n_3856),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4045),
.B(n_3885),
.Y(n_4143)
);

O2A1O1Ixp33_ASAP7_75t_L g4144 ( 
.A1(n_4033),
.A2(n_3875),
.B(n_3890),
.C(n_3849),
.Y(n_4144)
);

INVx4_ASAP7_75t_SL g4145 ( 
.A(n_3932),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_4018),
.B(n_3818),
.Y(n_4146)
);

OAI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3911),
.A2(n_3803),
.B1(n_3797),
.B2(n_3886),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3928),
.B(n_3847),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_3919),
.Y(n_4149)
);

OAI211xp5_ASAP7_75t_L g4150 ( 
.A1(n_3966),
.A2(n_3840),
.B(n_3793),
.C(n_115),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_3911),
.A2(n_3897),
.B1(n_3718),
.B2(n_3894),
.Y(n_4151)
);

OAI22xp5_ASAP7_75t_L g4152 ( 
.A1(n_3950),
.A2(n_3718),
.B1(n_3894),
.B2(n_115),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3909),
.B(n_3894),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3985),
.Y(n_4154)
);

O2A1O1Ixp5_ASAP7_75t_L g4155 ( 
.A1(n_3967),
.A2(n_3894),
.B(n_116),
.C(n_113),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_3904),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3988),
.B(n_114),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3906),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3993),
.B(n_117),
.Y(n_4159)
);

OR2x2_ASAP7_75t_L g4160 ( 
.A(n_3983),
.B(n_118),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3991),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4040),
.B(n_120),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3995),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_4040),
.B(n_121),
.Y(n_4164)
);

O2A1O1Ixp33_ASAP7_75t_L g4165 ( 
.A1(n_4030),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_4165)
);

O2A1O1Ixp33_ASAP7_75t_L g4166 ( 
.A1(n_3910),
.A2(n_125),
.B(n_122),
.C(n_124),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4004),
.Y(n_4167)
);

OR2x2_ASAP7_75t_L g4168 ( 
.A(n_4023),
.B(n_125),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_4025),
.B(n_127),
.Y(n_4169)
);

CKINVDCx9p33_ASAP7_75t_R g4170 ( 
.A(n_4054),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_4046),
.B(n_127),
.Y(n_4171)
);

OAI22xp5_ASAP7_75t_SL g4172 ( 
.A1(n_3999),
.A2(n_131),
.B1(n_128),
.B2(n_130),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_3931),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_3952),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_SL g4175 ( 
.A1(n_4059),
.A2(n_128),
.B(n_131),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_SL g4176 ( 
.A1(n_4000),
.A2(n_132),
.B(n_135),
.Y(n_4176)
);

OAI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_4057),
.A2(n_137),
.B1(n_132),
.B2(n_135),
.Y(n_4177)
);

OA21x2_ASAP7_75t_L g4178 ( 
.A1(n_4079),
.A2(n_137),
.B(n_138),
.Y(n_4178)
);

BUFx8_ASAP7_75t_SL g4179 ( 
.A(n_3922),
.Y(n_4179)
);

OR2x2_ASAP7_75t_L g4180 ( 
.A(n_4043),
.B(n_139),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_4043),
.B(n_140),
.Y(n_4181)
);

O2A1O1Ixp33_ASAP7_75t_L g4182 ( 
.A1(n_4069),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4058),
.Y(n_4183)
);

AND2x4_ASAP7_75t_L g4184 ( 
.A(n_4076),
.B(n_141),
.Y(n_4184)
);

NOR2xp67_ASAP7_75t_L g4185 ( 
.A(n_3915),
.B(n_143),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_3912),
.Y(n_4186)
);

NOR2xp67_ASAP7_75t_L g4187 ( 
.A(n_3915),
.B(n_3947),
.Y(n_4187)
);

AOI21xp5_ASAP7_75t_SL g4188 ( 
.A1(n_4006),
.A2(n_144),
.B(n_145),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3968),
.Y(n_4189)
);

AOI21x1_ASAP7_75t_SL g4190 ( 
.A1(n_3976),
.A2(n_144),
.B(n_147),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3980),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4021),
.B(n_4014),
.Y(n_4192)
);

OAI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_4053),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4067),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_4014),
.B(n_148),
.Y(n_4195)
);

NOR2xp67_ASAP7_75t_L g4196 ( 
.A(n_3947),
.B(n_150),
.Y(n_4196)
);

AOI21x1_ASAP7_75t_SL g4197 ( 
.A1(n_3918),
.A2(n_3964),
.B(n_3943),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4048),
.Y(n_4198)
);

CKINVDCx20_ASAP7_75t_R g4199 ( 
.A(n_3990),
.Y(n_4199)
);

NOR2xp33_ASAP7_75t_L g4200 ( 
.A(n_3914),
.B(n_3994),
.Y(n_4200)
);

OAI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3926),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4201)
);

BUFx3_ASAP7_75t_L g4202 ( 
.A(n_3970),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3986),
.A2(n_1367),
.B(n_1360),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4044),
.B(n_152),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3954),
.Y(n_4205)
);

O2A1O1Ixp33_ASAP7_75t_L g4206 ( 
.A1(n_3948),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_4206)
);

OAI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_4007),
.A2(n_159),
.B1(n_155),
.B2(n_156),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4077),
.A2(n_160),
.B1(n_156),
.B2(n_159),
.Y(n_4208)
);

AND2x2_ASAP7_75t_SL g4209 ( 
.A(n_4034),
.B(n_160),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4044),
.B(n_161),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_4076),
.B(n_161),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_3954),
.Y(n_4212)
);

OR2x2_ASAP7_75t_L g4213 ( 
.A(n_4071),
.B(n_4050),
.Y(n_4213)
);

O2A1O1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_3913),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_4214)
);

A2O1A1Ixp33_ASAP7_75t_L g4215 ( 
.A1(n_3942),
.A2(n_169),
.B(n_163),
.C(n_168),
.Y(n_4215)
);

BUFx4f_ASAP7_75t_SL g4216 ( 
.A(n_4116),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4183),
.Y(n_4217)
);

OAI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_4085),
.A2(n_4049),
.B1(n_3924),
.B2(n_3941),
.Y(n_4218)
);

AND2x4_ASAP7_75t_L g4219 ( 
.A(n_4124),
.B(n_4060),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4084),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_4113),
.Y(n_4221)
);

AO31x2_ASAP7_75t_L g4222 ( 
.A1(n_4081),
.A2(n_4051),
.A3(n_4070),
.B(n_3973),
.Y(n_4222)
);

NAND3xp33_ASAP7_75t_SL g4223 ( 
.A(n_4122),
.B(n_3953),
.C(n_3975),
.Y(n_4223)
);

AOI22xp33_ASAP7_75t_L g4224 ( 
.A1(n_4178),
.A2(n_3971),
.B1(n_3973),
.B2(n_3930),
.Y(n_4224)
);

OAI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_4090),
.A2(n_4049),
.B1(n_3924),
.B2(n_3941),
.Y(n_4225)
);

INVx4_ASAP7_75t_L g4226 ( 
.A(n_4105),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4092),
.Y(n_4227)
);

NAND2xp33_ASAP7_75t_R g4228 ( 
.A(n_4184),
.B(n_4061),
.Y(n_4228)
);

BUFx6f_ASAP7_75t_L g4229 ( 
.A(n_4186),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4134),
.Y(n_4230)
);

HB1xp67_ASAP7_75t_L g4231 ( 
.A(n_4128),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4109),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4088),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4137),
.B(n_4013),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4132),
.B(n_3933),
.Y(n_4235)
);

CKINVDCx5p33_ASAP7_75t_R g4236 ( 
.A(n_4179),
.Y(n_4236)
);

NOR2x1_ASAP7_75t_SL g4237 ( 
.A(n_4105),
.B(n_4009),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4098),
.Y(n_4238)
);

OR2x6_ASAP7_75t_L g4239 ( 
.A(n_4186),
.B(n_3996),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4133),
.Y(n_4240)
);

OR2x2_ASAP7_75t_L g4241 ( 
.A(n_4094),
.B(n_3937),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4138),
.Y(n_4242)
);

OAI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4086),
.A2(n_3933),
.B1(n_3937),
.B2(n_3996),
.Y(n_4243)
);

BUFx2_ASAP7_75t_L g4244 ( 
.A(n_4170),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4112),
.B(n_4102),
.Y(n_4245)
);

INVx8_ASAP7_75t_L g4246 ( 
.A(n_4105),
.Y(n_4246)
);

BUFx3_ASAP7_75t_L g4247 ( 
.A(n_4186),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4140),
.Y(n_4248)
);

HB1xp67_ASAP7_75t_L g4249 ( 
.A(n_4119),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4081),
.B(n_3989),
.Y(n_4250)
);

NAND3xp33_ASAP7_75t_SL g4251 ( 
.A(n_4083),
.B(n_3981),
.C(n_4072),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4154),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4161),
.Y(n_4253)
);

NAND2xp33_ASAP7_75t_R g4254 ( 
.A(n_4184),
.B(n_3997),
.Y(n_4254)
);

CKINVDCx5p33_ASAP7_75t_R g4255 ( 
.A(n_4199),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_4109),
.Y(n_4256)
);

OR2x6_ASAP7_75t_L g4257 ( 
.A(n_4202),
.B(n_3996),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4103),
.B(n_3989),
.Y(n_4258)
);

AOI22xp33_ASAP7_75t_L g4259 ( 
.A1(n_4178),
.A2(n_4172),
.B1(n_4100),
.B2(n_4148),
.Y(n_4259)
);

NAND4xp25_ASAP7_75t_L g4260 ( 
.A(n_4176),
.B(n_4097),
.C(n_4165),
.D(n_4182),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4099),
.B(n_4142),
.Y(n_4261)
);

CKINVDCx16_ASAP7_75t_R g4262 ( 
.A(n_4172),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_4143),
.B(n_3998),
.Y(n_4263)
);

BUFx2_ASAP7_75t_L g4264 ( 
.A(n_4145),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4108),
.Y(n_4265)
);

NAND2xp33_ASAP7_75t_R g4266 ( 
.A(n_4195),
.B(n_3997),
.Y(n_4266)
);

NOR2xp33_ASAP7_75t_R g4267 ( 
.A(n_4209),
.B(n_3998),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4163),
.B(n_4005),
.Y(n_4268)
);

NAND3xp33_ASAP7_75t_SL g4269 ( 
.A(n_4204),
.B(n_3965),
.C(n_3907),
.Y(n_4269)
);

OR2x2_ASAP7_75t_L g4270 ( 
.A(n_4089),
.B(n_4167),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4168),
.B(n_4005),
.Y(n_4271)
);

BUFx3_ASAP7_75t_L g4272 ( 
.A(n_4200),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4157),
.Y(n_4273)
);

BUFx3_ASAP7_75t_L g4274 ( 
.A(n_4159),
.Y(n_4274)
);

NAND2x1p5_ASAP7_75t_L g4275 ( 
.A(n_4196),
.B(n_4185),
.Y(n_4275)
);

XNOR2xp5_ASAP7_75t_L g4276 ( 
.A(n_4207),
.B(n_3916),
.Y(n_4276)
);

NAND2xp33_ASAP7_75t_R g4277 ( 
.A(n_4210),
.B(n_168),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4101),
.B(n_4011),
.Y(n_4278)
);

NAND2x1p5_ASAP7_75t_L g4279 ( 
.A(n_4162),
.B(n_4034),
.Y(n_4279)
);

AND2x4_ASAP7_75t_L g4280 ( 
.A(n_4187),
.B(n_3934),
.Y(n_4280)
);

AND2x4_ASAP7_75t_SL g4281 ( 
.A(n_4146),
.B(n_4011),
.Y(n_4281)
);

OR2x2_ASAP7_75t_L g4282 ( 
.A(n_4121),
.B(n_3937),
.Y(n_4282)
);

OAI221xp5_ASAP7_75t_L g4283 ( 
.A1(n_4207),
.A2(n_3908),
.B1(n_3982),
.B2(n_3959),
.C(n_3960),
.Y(n_4283)
);

INVx3_ASAP7_75t_L g4284 ( 
.A(n_4107),
.Y(n_4284)
);

BUFx6f_ASAP7_75t_L g4285 ( 
.A(n_4164),
.Y(n_4285)
);

AO31x2_ASAP7_75t_L g4286 ( 
.A1(n_4100),
.A2(n_4064),
.A3(n_4035),
.B(n_4034),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4095),
.B(n_3934),
.Y(n_4287)
);

BUFx2_ASAP7_75t_L g4288 ( 
.A(n_4145),
.Y(n_4288)
);

BUFx2_ASAP7_75t_R g4289 ( 
.A(n_4192),
.Y(n_4289)
);

CKINVDCx5p33_ASAP7_75t_R g4290 ( 
.A(n_4118),
.Y(n_4290)
);

AOI22xp33_ASAP7_75t_L g4291 ( 
.A1(n_4177),
.A2(n_4035),
.B1(n_4010),
.B2(n_4027),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4198),
.Y(n_4292)
);

AOI22xp33_ASAP7_75t_L g4293 ( 
.A1(n_4177),
.A2(n_4035),
.B1(n_4027),
.B2(n_3979),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4149),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_R g4295 ( 
.A(n_4180),
.B(n_3934),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_4093),
.Y(n_4296)
);

AOI22xp33_ASAP7_75t_L g4297 ( 
.A1(n_4193),
.A2(n_3979),
.B1(n_3921),
.B2(n_4078),
.Y(n_4297)
);

AOI221xp5_ASAP7_75t_L g4298 ( 
.A1(n_4206),
.A2(n_4066),
.B1(n_4063),
.B2(n_3907),
.C(n_4032),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4169),
.Y(n_4299)
);

INVx2_ASAP7_75t_SL g4300 ( 
.A(n_4213),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4106),
.B(n_3945),
.Y(n_4301)
);

CKINVDCx16_ASAP7_75t_R g4302 ( 
.A(n_4181),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4160),
.Y(n_4303)
);

NAND2xp33_ASAP7_75t_SL g4304 ( 
.A(n_4171),
.B(n_3945),
.Y(n_4304)
);

BUFx2_ASAP7_75t_SL g4305 ( 
.A(n_4197),
.Y(n_4305)
);

NAND2xp33_ASAP7_75t_R g4306 ( 
.A(n_4211),
.B(n_169),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4136),
.B(n_3945),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4093),
.Y(n_4308)
);

NAND3xp33_ASAP7_75t_SL g4309 ( 
.A(n_4155),
.B(n_4056),
.C(n_4015),
.Y(n_4309)
);

INVx3_ASAP7_75t_L g4310 ( 
.A(n_4107),
.Y(n_4310)
);

AOI22xp5_ASAP7_75t_L g4311 ( 
.A1(n_4150),
.A2(n_4002),
.B1(n_4074),
.B2(n_3956),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4110),
.Y(n_4312)
);

INVx6_ASAP7_75t_L g4313 ( 
.A(n_4153),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4096),
.B(n_4080),
.Y(n_4314)
);

CKINVDCx5p33_ASAP7_75t_R g4315 ( 
.A(n_4205),
.Y(n_4315)
);

AO31x2_ASAP7_75t_L g4316 ( 
.A1(n_4120),
.A2(n_4024),
.A3(n_178),
.B(n_171),
.Y(n_4316)
);

AND2x4_ASAP7_75t_L g4317 ( 
.A(n_4111),
.B(n_4115),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4104),
.B(n_171),
.Y(n_4318)
);

NOR2xp33_ASAP7_75t_R g4319 ( 
.A(n_4212),
.B(n_175),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_R g4320 ( 
.A(n_4111),
.B(n_175),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4110),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4156),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4117),
.B(n_4082),
.Y(n_4323)
);

OR2x2_ASAP7_75t_L g4324 ( 
.A(n_4130),
.B(n_180),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_4152),
.A2(n_3974),
.B1(n_3956),
.B2(n_3992),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4158),
.Y(n_4326)
);

A2O1A1Ixp33_ASAP7_75t_L g4327 ( 
.A1(n_4166),
.A2(n_4019),
.B(n_182),
.C(n_180),
.Y(n_4327)
);

CKINVDCx5p33_ASAP7_75t_R g4328 ( 
.A(n_4188),
.Y(n_4328)
);

CKINVDCx5p33_ASAP7_75t_R g4329 ( 
.A(n_4175),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4194),
.B(n_4127),
.Y(n_4330)
);

AOI22xp33_ASAP7_75t_L g4331 ( 
.A1(n_4193),
.A2(n_1374),
.B1(n_1383),
.B2(n_1367),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4189),
.Y(n_4332)
);

INVx2_ASAP7_75t_SL g4333 ( 
.A(n_4191),
.Y(n_4333)
);

INVxp67_ASAP7_75t_L g4334 ( 
.A(n_4208),
.Y(n_4334)
);

OAI21xp5_ASAP7_75t_SL g4335 ( 
.A1(n_4208),
.A2(n_181),
.B(n_183),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4173),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4091),
.B(n_181),
.Y(n_4337)
);

NAND2xp33_ASAP7_75t_R g4338 ( 
.A(n_4174),
.B(n_4087),
.Y(n_4338)
);

INVx5_ASAP7_75t_SL g4339 ( 
.A(n_4190),
.Y(n_4339)
);

INVxp67_ASAP7_75t_SL g4340 ( 
.A(n_4244),
.Y(n_4340)
);

AOI221xp5_ASAP7_75t_L g4341 ( 
.A1(n_4260),
.A2(n_4201),
.B1(n_4214),
.B2(n_4152),
.C(n_4215),
.Y(n_4341)
);

OR2x2_ASAP7_75t_L g4342 ( 
.A(n_4220),
.B(n_4091),
.Y(n_4342)
);

INVx3_ASAP7_75t_L g4343 ( 
.A(n_4226),
.Y(n_4343)
);

AND2x2_ASAP7_75t_SL g4344 ( 
.A(n_4262),
.B(n_4135),
.Y(n_4344)
);

INVx2_ASAP7_75t_SL g4345 ( 
.A(n_4246),
.Y(n_4345)
);

AO21x2_ASAP7_75t_L g4346 ( 
.A1(n_4312),
.A2(n_4321),
.B(n_4337),
.Y(n_4346)
);

OR2x2_ASAP7_75t_L g4347 ( 
.A(n_4227),
.B(n_4139),
.Y(n_4347)
);

AO21x2_ASAP7_75t_L g4348 ( 
.A1(n_4296),
.A2(n_4201),
.B(n_4203),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4259),
.A2(n_4123),
.B(n_4129),
.Y(n_4349)
);

OA21x2_ASAP7_75t_L g4350 ( 
.A1(n_4308),
.A2(n_4131),
.B(n_4126),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4333),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4217),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4230),
.Y(n_4353)
);

INVxp67_ASAP7_75t_SL g4354 ( 
.A(n_4334),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4261),
.B(n_4147),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4235),
.B(n_4147),
.Y(n_4356)
);

OAI21xp5_ASAP7_75t_L g4357 ( 
.A1(n_4335),
.A2(n_4139),
.B(n_4151),
.Y(n_4357)
);

NOR3xp33_ASAP7_75t_L g4358 ( 
.A(n_4223),
.B(n_4144),
.C(n_4151),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4232),
.B(n_4114),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4232),
.B(n_4087),
.Y(n_4360)
);

OA21x2_ASAP7_75t_L g4361 ( 
.A1(n_4250),
.A2(n_4141),
.B(n_4125),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4292),
.Y(n_4362)
);

BUFx2_ASAP7_75t_L g4363 ( 
.A(n_4264),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4294),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4233),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4238),
.Y(n_4366)
);

AOI221xp5_ASAP7_75t_L g4367 ( 
.A1(n_4276),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.C(n_189),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4240),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4256),
.B(n_4141),
.Y(n_4369)
);

HB1xp67_ASAP7_75t_L g4370 ( 
.A(n_4231),
.Y(n_4370)
);

OAI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_4329),
.A2(n_4328),
.B(n_4225),
.Y(n_4371)
);

AND2x4_ASAP7_75t_L g4372 ( 
.A(n_4256),
.B(n_187),
.Y(n_4372)
);

BUFx6f_ASAP7_75t_L g4373 ( 
.A(n_4229),
.Y(n_4373)
);

AO21x2_ASAP7_75t_L g4374 ( 
.A1(n_4318),
.A2(n_190),
.B(n_191),
.Y(n_4374)
);

OR2x6_ASAP7_75t_L g4375 ( 
.A(n_4246),
.B(n_190),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_SL g4376 ( 
.A1(n_4237),
.A2(n_192),
.B(n_193),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4317),
.B(n_195),
.Y(n_4377)
);

OA21x2_ASAP7_75t_L g4378 ( 
.A1(n_4314),
.A2(n_195),
.B(n_196),
.Y(n_4378)
);

OAI31xp33_ASAP7_75t_L g4379 ( 
.A1(n_4275),
.A2(n_199),
.A3(n_197),
.B(n_198),
.Y(n_4379)
);

BUFx4f_ASAP7_75t_SL g4380 ( 
.A(n_4229),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4242),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4322),
.Y(n_4382)
);

OA21x2_ASAP7_75t_L g4383 ( 
.A1(n_4245),
.A2(n_197),
.B(n_198),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4248),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_L g4385 ( 
.A1(n_4269),
.A2(n_203),
.B1(n_199),
.B2(n_201),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_4249),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4252),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4253),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4317),
.B(n_4323),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_4229),
.B(n_201),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4270),
.Y(n_4391)
);

OR2x2_ASAP7_75t_L g4392 ( 
.A(n_4265),
.B(n_203),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4287),
.B(n_206),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4326),
.Y(n_4394)
);

OAI21x1_ASAP7_75t_L g4395 ( 
.A1(n_4284),
.A2(n_206),
.B(n_207),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4284),
.B(n_207),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4221),
.Y(n_4397)
);

INVxp67_ASAP7_75t_SL g4398 ( 
.A(n_4306),
.Y(n_4398)
);

HB1xp67_ASAP7_75t_L g4399 ( 
.A(n_4273),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_4247),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4310),
.B(n_211),
.Y(n_4401)
);

OR2x2_ASAP7_75t_L g4402 ( 
.A(n_4299),
.B(n_212),
.Y(n_4402)
);

OAI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_4251),
.A2(n_212),
.B(n_213),
.Y(n_4403)
);

AOI21x1_ASAP7_75t_L g4404 ( 
.A1(n_4288),
.A2(n_214),
.B(n_215),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4332),
.Y(n_4405)
);

INVx3_ASAP7_75t_L g4406 ( 
.A(n_4226),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4303),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4268),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4324),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4300),
.B(n_214),
.Y(n_4410)
);

OAI321xp33_ASAP7_75t_L g4411 ( 
.A1(n_4224),
.A2(n_215),
.A3(n_216),
.B1(n_217),
.B2(n_218),
.C(n_219),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4222),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4278),
.B(n_216),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4302),
.B(n_218),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4263),
.B(n_220),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4271),
.Y(n_4416)
);

BUFx4f_ASAP7_75t_L g4417 ( 
.A(n_4239),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4222),
.Y(n_4418)
);

OA21x2_ASAP7_75t_L g4419 ( 
.A1(n_4307),
.A2(n_220),
.B(n_221),
.Y(n_4419)
);

OAI221xp5_ASAP7_75t_L g4420 ( 
.A1(n_4277),
.A2(n_223),
.B1(n_224),
.B2(n_227),
.C(n_228),
.Y(n_4420)
);

AND2x2_ASAP7_75t_L g4421 ( 
.A(n_4310),
.B(n_223),
.Y(n_4421)
);

OA21x2_ASAP7_75t_L g4422 ( 
.A1(n_4336),
.A2(n_228),
.B(n_229),
.Y(n_4422)
);

OR2x2_ASAP7_75t_L g4423 ( 
.A(n_4258),
.B(n_229),
.Y(n_4423)
);

INVx4_ASAP7_75t_L g4424 ( 
.A(n_4236),
.Y(n_4424)
);

OR2x2_ASAP7_75t_L g4425 ( 
.A(n_4282),
.B(n_230),
.Y(n_4425)
);

INVx3_ASAP7_75t_L g4426 ( 
.A(n_4313),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4281),
.B(n_230),
.Y(n_4427)
);

OR2x2_ASAP7_75t_L g4428 ( 
.A(n_4285),
.B(n_231),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4313),
.B(n_231),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4222),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4285),
.Y(n_4431)
);

OA21x2_ASAP7_75t_L g4432 ( 
.A1(n_4330),
.A2(n_232),
.B(n_233),
.Y(n_4432)
);

OR2x6_ASAP7_75t_L g4433 ( 
.A(n_4239),
.B(n_233),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4285),
.B(n_234),
.Y(n_4434)
);

OR2x6_ASAP7_75t_L g4435 ( 
.A(n_4257),
.B(n_234),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4274),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4422),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4340),
.B(n_4389),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4389),
.B(n_4237),
.Y(n_4439)
);

HB1xp67_ASAP7_75t_L g4440 ( 
.A(n_4370),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4426),
.B(n_4257),
.Y(n_4441)
);

INVxp67_ASAP7_75t_SL g4442 ( 
.A(n_4398),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4426),
.B(n_4305),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4432),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4422),
.Y(n_4445)
);

AND2x4_ASAP7_75t_SL g4446 ( 
.A(n_4426),
.B(n_4234),
.Y(n_4446)
);

INVx3_ASAP7_75t_L g4447 ( 
.A(n_4432),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4354),
.B(n_4339),
.Y(n_4448)
);

OAI222xp33_ASAP7_75t_L g4449 ( 
.A1(n_4342),
.A2(n_4338),
.B1(n_4243),
.B2(n_4286),
.C1(n_4283),
.C2(n_4293),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4399),
.B(n_4241),
.Y(n_4450)
);

OR2x2_ASAP7_75t_L g4451 ( 
.A(n_4399),
.B(n_4286),
.Y(n_4451)
);

OR2x2_ASAP7_75t_L g4452 ( 
.A(n_4407),
.B(n_4301),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4352),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4363),
.B(n_4219),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_SL g4455 ( 
.A(n_4357),
.B(n_4320),
.Y(n_4455)
);

OAI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4358),
.A2(n_4327),
.B(n_4309),
.Y(n_4456)
);

OR2x2_ASAP7_75t_L g4457 ( 
.A(n_4391),
.B(n_4286),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4422),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4355),
.B(n_4219),
.Y(n_4459)
);

OR2x2_ASAP7_75t_L g4460 ( 
.A(n_4370),
.B(n_4304),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4356),
.B(n_4289),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4409),
.B(n_4339),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4345),
.B(n_4280),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4365),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4345),
.B(n_4280),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4366),
.Y(n_4466)
);

AND2x4_ASAP7_75t_L g4467 ( 
.A(n_4343),
.B(n_4272),
.Y(n_4467)
);

INVxp67_ASAP7_75t_L g4468 ( 
.A(n_4400),
.Y(n_4468)
);

AND2x4_ASAP7_75t_L g4469 ( 
.A(n_4343),
.B(n_4290),
.Y(n_4469)
);

OR2x6_ASAP7_75t_SL g4470 ( 
.A(n_4436),
.B(n_4255),
.Y(n_4470)
);

INVx2_ASAP7_75t_L g4471 ( 
.A(n_4378),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4431),
.B(n_4218),
.Y(n_4472)
);

INVx3_ASAP7_75t_L g4473 ( 
.A(n_4432),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4368),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4381),
.Y(n_4475)
);

OR2x2_ASAP7_75t_L g4476 ( 
.A(n_4386),
.B(n_4279),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_4374),
.B(n_4267),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4384),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4374),
.B(n_4316),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4387),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4378),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4386),
.B(n_4316),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4349),
.B(n_4315),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4343),
.B(n_4316),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4373),
.B(n_4295),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4378),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4388),
.Y(n_4487)
);

OR2x2_ASAP7_75t_L g4488 ( 
.A(n_4405),
.B(n_4346),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4383),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4373),
.B(n_4319),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4373),
.B(n_4291),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4392),
.Y(n_4492)
);

OR2x2_ASAP7_75t_L g4493 ( 
.A(n_4416),
.B(n_4297),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4373),
.B(n_4228),
.Y(n_4494)
);

INVxp67_ASAP7_75t_SL g4495 ( 
.A(n_4400),
.Y(n_4495)
);

BUFx3_ASAP7_75t_L g4496 ( 
.A(n_4417),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4397),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4397),
.Y(n_4498)
);

BUFx3_ASAP7_75t_L g4499 ( 
.A(n_4417),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4383),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4406),
.B(n_4254),
.Y(n_4501)
);

BUFx12f_ASAP7_75t_L g4502 ( 
.A(n_4424),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_4344),
.B(n_4216),
.Y(n_4503)
);

OR2x2_ASAP7_75t_L g4504 ( 
.A(n_4347),
.B(n_4408),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4383),
.B(n_4331),
.Y(n_4505)
);

AOI22xp33_ASAP7_75t_L g4506 ( 
.A1(n_4346),
.A2(n_4298),
.B1(n_4325),
.B2(n_4311),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4419),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4402),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4440),
.Y(n_4509)
);

OAI221xp5_ASAP7_75t_SL g4510 ( 
.A1(n_4451),
.A2(n_4341),
.B1(n_4379),
.B2(n_4367),
.C(n_4420),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4444),
.Y(n_4511)
);

AOI22xp33_ASAP7_75t_L g4512 ( 
.A1(n_4444),
.A2(n_4348),
.B1(n_4344),
.B2(n_4350),
.Y(n_4512)
);

INVxp67_ASAP7_75t_L g4513 ( 
.A(n_4461),
.Y(n_4513)
);

AOI221xp5_ASAP7_75t_L g4514 ( 
.A1(n_4442),
.A2(n_4403),
.B1(n_4385),
.B2(n_4411),
.C(n_4348),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_R g4515 ( 
.A(n_4502),
.B(n_4380),
.Y(n_4515)
);

OAI211xp5_ASAP7_75t_SL g4516 ( 
.A1(n_4456),
.A2(n_4376),
.B(n_4423),
.C(n_4385),
.Y(n_4516)
);

NAND3xp33_ASAP7_75t_L g4517 ( 
.A(n_4506),
.B(n_4419),
.C(n_4376),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4461),
.B(n_4406),
.Y(n_4518)
);

OAI22xp5_ASAP7_75t_L g4519 ( 
.A1(n_4455),
.A2(n_4417),
.B1(n_4436),
.B2(n_4414),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4508),
.B(n_4429),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4488),
.Y(n_4521)
);

NOR2x1p5_ASAP7_75t_L g4522 ( 
.A(n_4495),
.B(n_4424),
.Y(n_4522)
);

AOI22xp33_ASAP7_75t_L g4523 ( 
.A1(n_4444),
.A2(n_4350),
.B1(n_4361),
.B2(n_4412),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_4503),
.B(n_4424),
.Y(n_4524)
);

NOR2x1_ASAP7_75t_SL g4525 ( 
.A(n_4503),
.B(n_4433),
.Y(n_4525)
);

BUFx3_ASAP7_75t_L g4526 ( 
.A(n_4470),
.Y(n_4526)
);

OAI31xp33_ASAP7_75t_SL g4527 ( 
.A1(n_4455),
.A2(n_4483),
.A3(n_4439),
.B(n_4438),
.Y(n_4527)
);

INVxp67_ASAP7_75t_L g4528 ( 
.A(n_4470),
.Y(n_4528)
);

OA21x2_ASAP7_75t_L g4529 ( 
.A1(n_4437),
.A2(n_4418),
.B(n_4412),
.Y(n_4529)
);

AO21x2_ASAP7_75t_L g4530 ( 
.A1(n_4489),
.A2(n_4430),
.B(n_4418),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_4438),
.Y(n_4531)
);

AOI22xp33_ASAP7_75t_L g4532 ( 
.A1(n_4447),
.A2(n_4350),
.B1(n_4361),
.B2(n_4353),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4447),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_4447),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_R g4535 ( 
.A1(n_4467),
.A2(n_4372),
.B(n_4380),
.Y(n_4535)
);

OAI221xp5_ASAP7_75t_L g4536 ( 
.A1(n_4473),
.A2(n_4361),
.B1(n_4371),
.B2(n_4433),
.C(n_4419),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4488),
.Y(n_4537)
);

NAND2xp33_ASAP7_75t_R g4538 ( 
.A(n_4490),
.B(n_4433),
.Y(n_4538)
);

NAND3xp33_ASAP7_75t_L g4539 ( 
.A(n_4473),
.B(n_4429),
.C(n_4406),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4459),
.B(n_4351),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4473),
.Y(n_4541)
);

HB1xp67_ASAP7_75t_L g4542 ( 
.A(n_4468),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4437),
.Y(n_4543)
);

OAI222xp33_ASAP7_75t_L g4544 ( 
.A1(n_4471),
.A2(n_4360),
.B1(n_4369),
.B2(n_4404),
.C1(n_4375),
.C2(n_4425),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4445),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4504),
.B(n_4372),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4459),
.B(n_4351),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4445),
.Y(n_4548)
);

NAND4xp75_ASAP7_75t_L g4549 ( 
.A(n_4483),
.B(n_4390),
.C(n_4427),
.D(n_4434),
.Y(n_4549)
);

AOI22xp33_ASAP7_75t_L g4550 ( 
.A1(n_4458),
.A2(n_4353),
.B1(n_4364),
.B2(n_4362),
.Y(n_4550)
);

OAI211xp5_ASAP7_75t_SL g4551 ( 
.A1(n_4448),
.A2(n_4451),
.B(n_4462),
.C(n_4460),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4453),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4458),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4531),
.B(n_4454),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4537),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4513),
.B(n_4494),
.Y(n_4556)
);

AND2x2_ASAP7_75t_SL g4557 ( 
.A(n_4527),
.B(n_4441),
.Y(n_4557)
);

OR2x2_ASAP7_75t_L g4558 ( 
.A(n_4509),
.B(n_4482),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4542),
.B(n_4454),
.Y(n_4559)
);

NAND2x1p5_ASAP7_75t_L g4560 ( 
.A(n_4522),
.B(n_4496),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4518),
.B(n_4494),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4537),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4518),
.B(n_4446),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4540),
.B(n_4493),
.Y(n_4564)
);

AOI22xp33_ASAP7_75t_L g4565 ( 
.A1(n_4517),
.A2(n_4471),
.B1(n_4486),
.B2(n_4481),
.Y(n_4565)
);

HB1xp67_ASAP7_75t_L g4566 ( 
.A(n_4511),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4543),
.Y(n_4567)
);

OR2x2_ASAP7_75t_L g4568 ( 
.A(n_4511),
.B(n_4482),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4533),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_4540),
.B(n_4507),
.Y(n_4570)
);

AND2x4_ASAP7_75t_L g4571 ( 
.A(n_4525),
.B(n_4496),
.Y(n_4571)
);

OR2x2_ASAP7_75t_L g4572 ( 
.A(n_4533),
.B(n_4464),
.Y(n_4572)
);

AND2x4_ASAP7_75t_L g4573 ( 
.A(n_4525),
.B(n_4499),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4547),
.B(n_4446),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4547),
.B(n_4501),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4534),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4526),
.B(n_4501),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4534),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4526),
.B(n_4443),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_4541),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4514),
.B(n_4507),
.Y(n_4581)
);

BUFx2_ASAP7_75t_L g4582 ( 
.A(n_4515),
.Y(n_4582)
);

OR2x2_ASAP7_75t_L g4583 ( 
.A(n_4570),
.B(n_4546),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4565),
.B(n_4545),
.Y(n_4584)
);

OR2x2_ASAP7_75t_L g4585 ( 
.A(n_4554),
.B(n_4450),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4566),
.B(n_4580),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4556),
.B(n_4545),
.Y(n_4587)
);

BUFx3_ASAP7_75t_L g4588 ( 
.A(n_4582),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4557),
.B(n_4441),
.Y(n_4589)
);

INVx2_ASAP7_75t_SL g4590 ( 
.A(n_4574),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4568),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4561),
.Y(n_4592)
);

OR2x2_ASAP7_75t_L g4593 ( 
.A(n_4559),
.B(n_4450),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4561),
.Y(n_4594)
);

OR2x2_ASAP7_75t_L g4595 ( 
.A(n_4564),
.B(n_4520),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4557),
.B(n_4441),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4568),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4556),
.B(n_4541),
.Y(n_4598)
);

HB1xp67_ASAP7_75t_L g4599 ( 
.A(n_4555),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4567),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4567),
.B(n_4553),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4575),
.B(n_4548),
.Y(n_4602)
);

NOR2xp33_ASAP7_75t_L g4603 ( 
.A(n_4582),
.B(n_4499),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4572),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4588),
.B(n_4574),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4589),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4596),
.B(n_4563),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4599),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4592),
.B(n_4575),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4599),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4586),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4594),
.B(n_4577),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4598),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4590),
.B(n_4577),
.Y(n_4614)
);

OR2x2_ASAP7_75t_L g4615 ( 
.A(n_4593),
.B(n_4558),
.Y(n_4615)
);

NAND2x1p5_ASAP7_75t_L g4616 ( 
.A(n_4603),
.B(n_4571),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4584),
.B(n_4555),
.Y(n_4617)
);

HB1xp67_ASAP7_75t_L g4618 ( 
.A(n_4586),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4602),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4609),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4609),
.Y(n_4621)
);

NOR2xp67_ASAP7_75t_SL g4622 ( 
.A(n_4618),
.B(n_4502),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4612),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4615),
.Y(n_4624)
);

OAI22xp5_ASAP7_75t_L g4625 ( 
.A1(n_4606),
.A2(n_4535),
.B1(n_4528),
.B2(n_4510),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4614),
.Y(n_4626)
);

NOR2xp33_ASAP7_75t_L g4627 ( 
.A(n_4616),
.B(n_4571),
.Y(n_4627)
);

NAND3xp33_ASAP7_75t_L g4628 ( 
.A(n_4617),
.B(n_4584),
.C(n_4605),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4624),
.Y(n_4629)
);

NOR2xp33_ASAP7_75t_L g4630 ( 
.A(n_4627),
.B(n_4571),
.Y(n_4630)
);

AOI22xp33_ASAP7_75t_L g4631 ( 
.A1(n_4628),
.A2(n_4581),
.B1(n_4543),
.B2(n_4500),
.Y(n_4631)
);

OR2x2_ASAP7_75t_L g4632 ( 
.A(n_4620),
.B(n_4602),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4623),
.B(n_4563),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4621),
.B(n_4607),
.Y(n_4634)
);

NOR2xp33_ASAP7_75t_SL g4635 ( 
.A(n_4622),
.B(n_4616),
.Y(n_4635)
);

NOR2xp33_ASAP7_75t_L g4636 ( 
.A(n_4625),
.B(n_4573),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4626),
.B(n_4613),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4624),
.B(n_4619),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4624),
.Y(n_4639)
);

OR2x2_ASAP7_75t_L g4640 ( 
.A(n_4628),
.B(n_4585),
.Y(n_4640)
);

XOR2x2_ASAP7_75t_L g4641 ( 
.A(n_4636),
.B(n_4549),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_4640),
.A2(n_4539),
.B1(n_4595),
.B2(n_4583),
.Y(n_4642)
);

OAI32xp33_ASAP7_75t_L g4643 ( 
.A1(n_4632),
.A2(n_4617),
.A3(n_4560),
.B1(n_4587),
.B2(n_4558),
.Y(n_4643)
);

AOI21xp33_ASAP7_75t_SL g4644 ( 
.A1(n_4630),
.A2(n_4573),
.B(n_4560),
.Y(n_4644)
);

OAI221xp5_ASAP7_75t_L g4645 ( 
.A1(n_4631),
.A2(n_4536),
.B1(n_4512),
.B2(n_4532),
.C(n_4523),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4634),
.Y(n_4646)
);

AOI22xp5_ASAP7_75t_L g4647 ( 
.A1(n_4629),
.A2(n_4538),
.B1(n_4573),
.B2(n_4519),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4633),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4639),
.B(n_4604),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4648),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4646),
.B(n_4591),
.Y(n_4651)
);

INVx1_ASAP7_75t_SL g4652 ( 
.A(n_4641),
.Y(n_4652)
);

NAND2xp33_ASAP7_75t_SL g4653 ( 
.A(n_4649),
.B(n_4587),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4642),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4643),
.Y(n_4655)
);

NOR3xp33_ASAP7_75t_SL g4656 ( 
.A(n_4645),
.B(n_4637),
.C(n_4638),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4650),
.B(n_4597),
.Y(n_4657)
);

INVx1_ASAP7_75t_SL g4658 ( 
.A(n_4653),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4651),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4654),
.B(n_4579),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4656),
.B(n_4579),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4655),
.B(n_4611),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4652),
.B(n_4560),
.Y(n_4663)
);

NOR2x1_ASAP7_75t_L g4664 ( 
.A(n_4657),
.B(n_4608),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4660),
.B(n_4600),
.Y(n_4665)
);

A2O1A1Ixp33_ASAP7_75t_L g4666 ( 
.A1(n_4663),
.A2(n_4647),
.B(n_4644),
.C(n_4562),
.Y(n_4666)
);

NAND3xp33_ASAP7_75t_SL g4667 ( 
.A(n_4658),
.B(n_4635),
.C(n_4610),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4661),
.Y(n_4668)
);

INVxp67_ASAP7_75t_L g4669 ( 
.A(n_4662),
.Y(n_4669)
);

NAND4xp25_ASAP7_75t_L g4670 ( 
.A(n_4658),
.B(n_4635),
.C(n_4601),
.D(n_4524),
.Y(n_4670)
);

A2O1A1Ixp33_ASAP7_75t_SL g4671 ( 
.A1(n_4659),
.A2(n_4562),
.B(n_4521),
.C(n_4569),
.Y(n_4671)
);

AND4x1_ASAP7_75t_L g4672 ( 
.A(n_4660),
.B(n_4601),
.C(n_4578),
.D(n_4576),
.Y(n_4672)
);

NOR3x1_ASAP7_75t_L g4673 ( 
.A(n_4657),
.B(n_4549),
.C(n_4572),
.Y(n_4673)
);

OAI21xp5_ASAP7_75t_SL g4674 ( 
.A1(n_4661),
.A2(n_4551),
.B(n_4544),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_4663),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4660),
.B(n_4548),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4660),
.Y(n_4677)
);

NAND4xp25_ASAP7_75t_SL g4678 ( 
.A(n_4657),
.B(n_4553),
.C(n_4552),
.D(n_4439),
.Y(n_4678)
);

NOR2xp33_ASAP7_75t_L g4679 ( 
.A(n_4669),
.B(n_4477),
.Y(n_4679)
);

OR2x2_ASAP7_75t_L g4680 ( 
.A(n_4667),
.B(n_4457),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4664),
.B(n_4530),
.Y(n_4681)
);

AOI221xp5_ASAP7_75t_SL g4682 ( 
.A1(n_4670),
.A2(n_4480),
.B1(n_4478),
.B2(n_4475),
.C(n_4474),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4677),
.B(n_4469),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4674),
.B(n_4530),
.Y(n_4684)
);

AOI21xp5_ASAP7_75t_L g4685 ( 
.A1(n_4671),
.A2(n_4469),
.B(n_4530),
.Y(n_4685)
);

NOR3xp33_ASAP7_75t_L g4686 ( 
.A(n_4668),
.B(n_4516),
.C(n_4486),
.Y(n_4686)
);

AOI22xp5_ASAP7_75t_L g4687 ( 
.A1(n_4675),
.A2(n_4490),
.B1(n_4500),
.B2(n_4489),
.Y(n_4687)
);

INVxp67_ASAP7_75t_L g4688 ( 
.A(n_4665),
.Y(n_4688)
);

AOI211xp5_ASAP7_75t_L g4689 ( 
.A1(n_4666),
.A2(n_4390),
.B(n_4449),
.C(n_4484),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_SL g4690 ( 
.A(n_4672),
.B(n_4467),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4673),
.B(n_4481),
.Y(n_4691)
);

OAI321xp33_ASAP7_75t_L g4692 ( 
.A1(n_4676),
.A2(n_4550),
.A3(n_4375),
.B1(n_4457),
.B2(n_4479),
.C(n_4505),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4678),
.Y(n_4693)
);

OR2x2_ASAP7_75t_L g4694 ( 
.A(n_4667),
.B(n_4467),
.Y(n_4694)
);

AOI21xp5_ASAP7_75t_L g4695 ( 
.A1(n_4667),
.A2(n_4469),
.B(n_4529),
.Y(n_4695)
);

OAI22xp33_ASAP7_75t_L g4696 ( 
.A1(n_4676),
.A2(n_4529),
.B1(n_4375),
.B2(n_4460),
.Y(n_4696)
);

OAI22xp33_ASAP7_75t_L g4697 ( 
.A1(n_4676),
.A2(n_4529),
.B1(n_4435),
.B2(n_4410),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_SL g4698 ( 
.A(n_4675),
.B(n_4443),
.Y(n_4698)
);

AOI22xp33_ASAP7_75t_L g4699 ( 
.A1(n_4669),
.A2(n_4484),
.B1(n_4498),
.B2(n_4497),
.Y(n_4699)
);

NOR3x1_ASAP7_75t_L g4700 ( 
.A(n_4667),
.B(n_4487),
.C(n_4466),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4669),
.B(n_4463),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4664),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4667),
.B(n_4492),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4701),
.Y(n_4704)
);

NOR4xp25_ASAP7_75t_L g4705 ( 
.A(n_4702),
.B(n_4491),
.C(n_4428),
.D(n_4472),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4680),
.A2(n_4694),
.B1(n_4703),
.B2(n_4687),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4681),
.Y(n_4707)
);

AOI211xp5_ASAP7_75t_L g4708 ( 
.A1(n_4695),
.A2(n_4484),
.B(n_4491),
.C(n_4485),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4683),
.Y(n_4709)
);

NOR3xp33_ASAP7_75t_L g4710 ( 
.A(n_4688),
.B(n_4485),
.C(n_4465),
.Y(n_4710)
);

NAND4xp25_ASAP7_75t_L g4711 ( 
.A(n_4679),
.B(n_4266),
.C(n_4465),
.D(n_4463),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4691),
.Y(n_4712)
);

NOR5xp2_ASAP7_75t_L g4713 ( 
.A(n_4693),
.B(n_4472),
.C(n_4435),
.D(n_4476),
.E(n_4377),
.Y(n_4713)
);

NAND3xp33_ASAP7_75t_L g4714 ( 
.A(n_4684),
.B(n_4435),
.C(n_4427),
.Y(n_4714)
);

NOR3xp33_ASAP7_75t_L g4715 ( 
.A(n_4698),
.B(n_4393),
.C(n_4372),
.Y(n_4715)
);

AND3x1_ASAP7_75t_L g4716 ( 
.A(n_4685),
.B(n_4377),
.C(n_4396),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_4696),
.B(n_4393),
.Y(n_4717)
);

AOI22xp33_ASAP7_75t_L g4718 ( 
.A1(n_4686),
.A2(n_4369),
.B1(n_4360),
.B2(n_4421),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4697),
.B(n_4415),
.Y(n_4719)
);

NAND4xp25_ASAP7_75t_L g4720 ( 
.A(n_4700),
.B(n_4421),
.C(n_4401),
.D(n_4396),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4690),
.B(n_4452),
.Y(n_4721)
);

OAI211xp5_ASAP7_75t_SL g4722 ( 
.A1(n_4699),
.A2(n_236),
.B(n_237),
.C(n_238),
.Y(n_4722)
);

OAI22xp33_ASAP7_75t_L g4723 ( 
.A1(n_4692),
.A2(n_4413),
.B1(n_4382),
.B2(n_4394),
.Y(n_4723)
);

NAND3xp33_ASAP7_75t_L g4724 ( 
.A(n_4689),
.B(n_4401),
.C(n_4364),
.Y(n_4724)
);

AOI221xp5_ASAP7_75t_L g4725 ( 
.A1(n_4682),
.A2(n_4362),
.B1(n_4382),
.B2(n_4394),
.C(n_4359),
.Y(n_4725)
);

NOR2xp67_ASAP7_75t_L g4726 ( 
.A(n_4694),
.B(n_236),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4701),
.Y(n_4727)
);

NOR3xp33_ASAP7_75t_L g4728 ( 
.A(n_4702),
.B(n_4395),
.C(n_237),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4685),
.B(n_4395),
.Y(n_4729)
);

NAND5xp2_ASAP7_75t_L g4730 ( 
.A(n_4679),
.B(n_4359),
.C(n_240),
.D(n_241),
.E(n_242),
.Y(n_4730)
);

O2A1O1Ixp33_ASAP7_75t_SL g4731 ( 
.A1(n_4690),
.A2(n_238),
.B(n_240),
.C(n_243),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_4730),
.B(n_244),
.Y(n_4732)
);

AOI221xp5_ASAP7_75t_L g4733 ( 
.A1(n_4706),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.C(n_247),
.Y(n_4733)
);

NOR3xp33_ASAP7_75t_SL g4734 ( 
.A(n_4712),
.B(n_246),
.C(n_249),
.Y(n_4734)
);

NAND3xp33_ASAP7_75t_SL g4735 ( 
.A(n_4709),
.B(n_249),
.C(n_250),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4715),
.B(n_250),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4705),
.B(n_251),
.Y(n_4737)
);

NAND4xp75_ASAP7_75t_L g4738 ( 
.A(n_4726),
.B(n_252),
.C(n_256),
.D(n_257),
.Y(n_4738)
);

NAND4xp25_ASAP7_75t_SL g4739 ( 
.A(n_4708),
.B(n_252),
.C(n_256),
.D(n_257),
.Y(n_4739)
);

NOR3xp33_ASAP7_75t_SL g4740 ( 
.A(n_4704),
.B(n_258),
.C(n_259),
.Y(n_4740)
);

OAI22xp5_ASAP7_75t_L g4741 ( 
.A1(n_4716),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_4741)
);

OAI211xp5_ASAP7_75t_L g4742 ( 
.A1(n_4727),
.A2(n_262),
.B(n_264),
.C(n_265),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4721),
.Y(n_4743)
);

NOR2xp33_ASAP7_75t_SL g4744 ( 
.A(n_4714),
.B(n_262),
.Y(n_4744)
);

NAND4xp25_ASAP7_75t_L g4745 ( 
.A(n_4710),
.B(n_264),
.C(n_266),
.D(n_267),
.Y(n_4745)
);

AOI221xp5_ASAP7_75t_L g4746 ( 
.A1(n_4731),
.A2(n_266),
.B1(n_268),
.B2(n_270),
.C(n_271),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4723),
.B(n_268),
.Y(n_4747)
);

AOI211xp5_ASAP7_75t_L g4748 ( 
.A1(n_4722),
.A2(n_271),
.B(n_272),
.C(n_273),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_SL g4749 ( 
.A(n_4729),
.B(n_272),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4717),
.Y(n_4750)
);

OR2x2_ASAP7_75t_L g4751 ( 
.A(n_4720),
.B(n_275),
.Y(n_4751)
);

AOI211xp5_ASAP7_75t_L g4752 ( 
.A1(n_4707),
.A2(n_276),
.B(n_277),
.C(n_281),
.Y(n_4752)
);

NAND4xp25_ASAP7_75t_L g4753 ( 
.A(n_4713),
.B(n_276),
.C(n_282),
.D(n_283),
.Y(n_4753)
);

AOI211xp5_ASAP7_75t_L g4754 ( 
.A1(n_4711),
.A2(n_284),
.B(n_285),
.C(n_286),
.Y(n_4754)
);

NOR2x1_ASAP7_75t_SL g4755 ( 
.A(n_4719),
.B(n_285),
.Y(n_4755)
);

NAND4xp25_ASAP7_75t_SL g4756 ( 
.A(n_4728),
.B(n_286),
.C(n_287),
.D(n_288),
.Y(n_4756)
);

AOI222xp33_ASAP7_75t_L g4757 ( 
.A1(n_4755),
.A2(n_4724),
.B1(n_4725),
.B2(n_4718),
.C1(n_291),
.C2(n_292),
.Y(n_4757)
);

XNOR2xp5_ASAP7_75t_L g4758 ( 
.A(n_4738),
.B(n_288),
.Y(n_4758)
);

NOR3xp33_ASAP7_75t_L g4759 ( 
.A(n_4743),
.B(n_4750),
.C(n_4737),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4753),
.B(n_289),
.Y(n_4760)
);

CKINVDCx20_ASAP7_75t_R g4761 ( 
.A(n_4732),
.Y(n_4761)
);

OAI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4749),
.A2(n_289),
.B(n_290),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4740),
.Y(n_4763)
);

OAI211xp5_ASAP7_75t_L g4764 ( 
.A1(n_4733),
.A2(n_292),
.B(n_296),
.C(n_298),
.Y(n_4764)
);

CKINVDCx20_ASAP7_75t_R g4765 ( 
.A(n_4734),
.Y(n_4765)
);

XNOR2xp5_ASAP7_75t_L g4766 ( 
.A(n_4754),
.B(n_298),
.Y(n_4766)
);

HB1xp67_ASAP7_75t_L g4767 ( 
.A(n_4741),
.Y(n_4767)
);

AOI221xp5_ASAP7_75t_L g4768 ( 
.A1(n_4739),
.A2(n_4756),
.B1(n_4746),
.B2(n_4735),
.C(n_4747),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4748),
.B(n_299),
.Y(n_4769)
);

INVx1_ASAP7_75t_SL g4770 ( 
.A(n_4751),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4736),
.Y(n_4771)
);

INVx2_ASAP7_75t_SL g4772 ( 
.A(n_4744),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4752),
.B(n_299),
.Y(n_4773)
);

NOR2xp33_ASAP7_75t_L g4774 ( 
.A(n_4745),
.B(n_4742),
.Y(n_4774)
);

XNOR2xp5_ASAP7_75t_L g4775 ( 
.A(n_4761),
.B(n_300),
.Y(n_4775)
);

NAND2xp33_ASAP7_75t_L g4776 ( 
.A(n_4760),
.B(n_301),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4758),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4765),
.Y(n_4778)
);

NOR2x1_ASAP7_75t_L g4779 ( 
.A(n_4763),
.B(n_301),
.Y(n_4779)
);

NOR2x1_ASAP7_75t_L g4780 ( 
.A(n_4771),
.B(n_302),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4766),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_4772),
.B(n_4769),
.Y(n_4782)
);

AOI22xp5_ASAP7_75t_L g4783 ( 
.A1(n_4759),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4767),
.Y(n_4784)
);

NOR2x1_ASAP7_75t_L g4785 ( 
.A(n_4773),
.B(n_303),
.Y(n_4785)
);

XOR2x2_ASAP7_75t_L g4786 ( 
.A(n_4768),
.B(n_304),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4774),
.Y(n_4787)
);

NOR3xp33_ASAP7_75t_L g4788 ( 
.A(n_4770),
.B(n_305),
.C(n_306),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4762),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4779),
.Y(n_4790)
);

XNOR2xp5_ASAP7_75t_L g4791 ( 
.A(n_4786),
.B(n_4764),
.Y(n_4791)
);

AND2x2_ASAP7_75t_SL g4792 ( 
.A(n_4776),
.B(n_4757),
.Y(n_4792)
);

XNOR2x1_ASAP7_75t_L g4793 ( 
.A(n_4784),
.B(n_307),
.Y(n_4793)
);

AND2x4_ASAP7_75t_L g4794 ( 
.A(n_4778),
.B(n_307),
.Y(n_4794)
);

AND2x4_ASAP7_75t_L g4795 ( 
.A(n_4787),
.B(n_308),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_SL g4796 ( 
.A(n_4780),
.B(n_309),
.Y(n_4796)
);

NAND3xp33_ASAP7_75t_L g4797 ( 
.A(n_4785),
.B(n_1374),
.C(n_1383),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4777),
.B(n_310),
.Y(n_4798)
);

NAND4xp25_ASAP7_75t_L g4799 ( 
.A(n_4788),
.B(n_310),
.C(n_311),
.D(n_313),
.Y(n_4799)
);

OAI211xp5_ASAP7_75t_SL g4800 ( 
.A1(n_4782),
.A2(n_311),
.B(n_314),
.C(n_315),
.Y(n_4800)
);

INVxp67_ASAP7_75t_L g4801 ( 
.A(n_4775),
.Y(n_4801)
);

AO211x2_ASAP7_75t_L g4802 ( 
.A1(n_4781),
.A2(n_316),
.B(n_317),
.C(n_318),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4790),
.Y(n_4803)
);

CKINVDCx20_ASAP7_75t_R g4804 ( 
.A(n_4801),
.Y(n_4804)
);

NAND2xp33_ASAP7_75t_L g4805 ( 
.A(n_4798),
.B(n_4783),
.Y(n_4805)
);

AOI21xp5_ASAP7_75t_L g4806 ( 
.A1(n_4793),
.A2(n_4789),
.B(n_318),
.Y(n_4806)
);

CKINVDCx5p33_ASAP7_75t_R g4807 ( 
.A(n_4791),
.Y(n_4807)
);

CKINVDCx20_ASAP7_75t_R g4808 ( 
.A(n_4796),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4795),
.Y(n_4809)
);

CKINVDCx5p33_ASAP7_75t_R g4810 ( 
.A(n_4792),
.Y(n_4810)
);

INVx1_ASAP7_75t_SL g4811 ( 
.A(n_4794),
.Y(n_4811)
);

INVx1_ASAP7_75t_SL g4812 ( 
.A(n_4797),
.Y(n_4812)
);

AOI322xp5_ASAP7_75t_L g4813 ( 
.A1(n_4804),
.A2(n_4810),
.A3(n_4803),
.B1(n_4807),
.B2(n_4811),
.C1(n_4808),
.C2(n_4809),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4805),
.A2(n_4800),
.B1(n_4799),
.B2(n_4802),
.Y(n_4814)
);

OAI211xp5_ASAP7_75t_SL g4815 ( 
.A1(n_4806),
.A2(n_316),
.B(n_321),
.C(n_323),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4812),
.Y(n_4816)
);

O2A1O1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4803),
.A2(n_321),
.B(n_323),
.C(n_324),
.Y(n_4817)
);

AOI221xp5_ASAP7_75t_L g4818 ( 
.A1(n_4810),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_4818)
);

AOI221xp5_ASAP7_75t_L g4819 ( 
.A1(n_4810),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.C(n_330),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4816),
.Y(n_4820)
);

OAI22xp5_ASAP7_75t_SL g4821 ( 
.A1(n_4814),
.A2(n_328),
.B1(n_330),
.B2(n_332),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4815),
.Y(n_4822)
);

AOI321xp33_ASAP7_75t_L g4823 ( 
.A1(n_4820),
.A2(n_4822),
.A3(n_4813),
.B1(n_4817),
.B2(n_4818),
.C(n_4819),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4821),
.B(n_336),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4824),
.B(n_336),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_SL g4826 ( 
.A(n_4823),
.B(n_1374),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4826),
.A2(n_1383),
.B(n_1374),
.Y(n_4827)
);

AOI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4825),
.A2(n_1383),
.B(n_338),
.Y(n_4828)
);

OAI22xp5_ASAP7_75t_L g4829 ( 
.A1(n_4825),
.A2(n_339),
.B1(n_1925),
.B2(n_344),
.Y(n_4829)
);

OAI22xp5_ASAP7_75t_SL g4830 ( 
.A1(n_4829),
.A2(n_1925),
.B1(n_346),
.B2(n_347),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4828),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4827),
.A2(n_1925),
.B(n_1432),
.Y(n_4832)
);

AOI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_4829),
.A2(n_1925),
.B1(n_348),
.B2(n_350),
.Y(n_4833)
);

NOR2xp67_ASAP7_75t_L g4834 ( 
.A(n_4831),
.B(n_342),
.Y(n_4834)
);

AO21x2_ASAP7_75t_L g4835 ( 
.A1(n_4832),
.A2(n_355),
.B(n_356),
.Y(n_4835)
);

INVxp67_ASAP7_75t_L g4836 ( 
.A(n_4830),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4833),
.B(n_359),
.Y(n_4837)
);

AOI22xp5_ASAP7_75t_L g4838 ( 
.A1(n_4831),
.A2(n_364),
.B1(n_366),
.B2(n_368),
.Y(n_4838)
);

OA22x2_ASAP7_75t_L g4839 ( 
.A1(n_4836),
.A2(n_373),
.B1(n_382),
.B2(n_384),
.Y(n_4839)
);

AOI22xp33_ASAP7_75t_SL g4840 ( 
.A1(n_4837),
.A2(n_385),
.B1(n_388),
.B2(n_397),
.Y(n_4840)
);

AOI22xp5_ASAP7_75t_L g4841 ( 
.A1(n_4835),
.A2(n_399),
.B1(n_401),
.B2(n_403),
.Y(n_4841)
);

AOI22xp5_ASAP7_75t_L g4842 ( 
.A1(n_4834),
.A2(n_408),
.B1(n_413),
.B2(n_415),
.Y(n_4842)
);

AOI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_4838),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_4843)
);

OAI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4836),
.A2(n_424),
.B1(n_426),
.B2(n_429),
.Y(n_4844)
);

AO22x2_ASAP7_75t_L g4845 ( 
.A1(n_4836),
.A2(n_436),
.B1(n_437),
.B2(n_442),
.Y(n_4845)
);

OAI22xp33_ASAP7_75t_L g4846 ( 
.A1(n_4836),
.A2(n_443),
.B1(n_446),
.B2(n_450),
.Y(n_4846)
);

AOI22xp5_ASAP7_75t_L g4847 ( 
.A1(n_4836),
.A2(n_451),
.B1(n_452),
.B2(n_454),
.Y(n_4847)
);

AOI22xp5_ASAP7_75t_L g4848 ( 
.A1(n_4836),
.A2(n_455),
.B1(n_461),
.B2(n_465),
.Y(n_4848)
);

AOI22xp5_ASAP7_75t_L g4849 ( 
.A1(n_4836),
.A2(n_468),
.B1(n_470),
.B2(n_472),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4839),
.Y(n_4850)
);

OA21x2_ASAP7_75t_L g4851 ( 
.A1(n_4841),
.A2(n_473),
.B(n_474),
.Y(n_4851)
);

NOR2xp33_ASAP7_75t_L g4852 ( 
.A(n_4843),
.B(n_475),
.Y(n_4852)
);

OAI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4840),
.A2(n_477),
.B(n_479),
.Y(n_4853)
);

NAND2x1p5_ASAP7_75t_L g4854 ( 
.A(n_4842),
.B(n_1407),
.Y(n_4854)
);

OAI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4844),
.A2(n_482),
.B(n_486),
.Y(n_4855)
);

OAI21x1_ASAP7_75t_L g4856 ( 
.A1(n_4849),
.A2(n_487),
.B(n_490),
.Y(n_4856)
);

AO21x2_ASAP7_75t_L g4857 ( 
.A1(n_4846),
.A2(n_492),
.B(n_494),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4850),
.B(n_4845),
.Y(n_4858)
);

BUFx2_ASAP7_75t_L g4859 ( 
.A(n_4854),
.Y(n_4859)
);

AOI21xp5_ASAP7_75t_L g4860 ( 
.A1(n_4852),
.A2(n_4848),
.B(n_4847),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4851),
.Y(n_4861)
);

HB1xp67_ASAP7_75t_L g4862 ( 
.A(n_4857),
.Y(n_4862)
);

AOI221x1_ASAP7_75t_L g4863 ( 
.A1(n_4858),
.A2(n_4855),
.B1(n_4853),
.B2(n_4856),
.C(n_503),
.Y(n_4863)
);

AOI221xp5_ASAP7_75t_L g4864 ( 
.A1(n_4861),
.A2(n_495),
.B1(n_497),
.B2(n_500),
.C(n_512),
.Y(n_4864)
);

AOI211xp5_ASAP7_75t_L g4865 ( 
.A1(n_4863),
.A2(n_4862),
.B(n_4859),
.C(n_4860),
.Y(n_4865)
);

AOI211xp5_ASAP7_75t_L g4866 ( 
.A1(n_4865),
.A2(n_4864),
.B(n_516),
.C(n_519),
.Y(n_4866)
);


endmodule