module fake_jpeg_23461_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_46),
.B1(n_34),
.B2(n_31),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_36),
.B1(n_34),
.B2(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_79),
.B1(n_55),
.B2(n_34),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_61),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_1),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_87),
.C(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_26),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_29),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_39),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_88),
.B1(n_29),
.B2(n_31),
.Y(n_115)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

OR2x4_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_51),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_66),
.B1(n_75),
.B2(n_74),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_15),
.Y(n_128)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_39),
.C(n_37),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_116),
.C(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_55),
.B1(n_53),
.B2(n_42),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_111),
.B1(n_117),
.B2(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_37),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_41),
.C(n_42),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_38),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_38),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_136),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_129),
.B1(n_141),
.B2(n_144),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_63),
.Y(n_127)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_71),
.B1(n_81),
.B2(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_31),
.B(n_29),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_138),
.B(n_143),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_80),
.C(n_61),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_80),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_149),
.C(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_145),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_140),
.B1(n_23),
.B2(n_25),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_69),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_100),
.B1(n_97),
.B2(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_1),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_78),
.B1(n_27),
.B2(n_32),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_16),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_93),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_27),
.B1(n_32),
.B2(n_69),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_94),
.B1(n_33),
.B2(n_30),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_1),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_2),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_61),
.C(n_21),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_93),
.B1(n_105),
.B2(n_101),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_167),
.B1(n_176),
.B2(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_175),
.B1(n_8),
.B2(n_4),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_118),
.B1(n_99),
.B2(n_27),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_143),
.C(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_178),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_32),
.B(n_33),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_159),
.B(n_161),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_30),
.B1(n_24),
.B2(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_33),
.B1(n_30),
.B2(n_24),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_33),
.B1(n_30),
.B2(n_21),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_24),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_148),
.B(n_24),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_128),
.C(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_192),
.C(n_206),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_125),
.B(n_128),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_191),
.B(n_201),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_148),
.C(n_112),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_196),
.B1(n_200),
.B2(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_208),
.Y(n_216)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_2),
.B1(n_3),
.B2(n_14),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_202),
.B1(n_174),
.B2(n_172),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_155),
.B1(n_179),
.B2(n_167),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_2),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_7),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_14),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_165),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_222),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_205),
.B(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_214),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_228),
.B1(n_195),
.B2(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_186),
.B(n_169),
.Y(n_222)
);

NAND4xp25_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_152),
.C(n_153),
.D(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_181),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_165),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_166),
.B1(n_172),
.B2(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

XOR2x1_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_166),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_203),
.C(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_233),
.C(n_211),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_203),
.C(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_237),
.B1(n_239),
.B2(n_244),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_189),
.B1(n_193),
.B2(n_188),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_201),
.B1(n_191),
.B2(n_190),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_230),
.A2(n_201),
.B1(n_5),
.B2(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_253),
.C(n_231),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_210),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_252),
.B1(n_233),
.B2(n_3),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_220),
.B1(n_226),
.B2(n_213),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_240),
.B(n_245),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_7),
.B(n_10),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_263),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_229),
.B1(n_220),
.B2(n_212),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_261),
.B1(n_247),
.B2(n_238),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_217),
.B(n_211),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_221),
.B1(n_5),
.B2(n_6),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_232),
.B(n_221),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_255),
.A2(n_252),
.B1(n_258),
.B2(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_274),
.B1(n_11),
.B2(n_13),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_262),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_270),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_252),
.B(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_10),
.C(n_11),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_275),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_11),
.B1(n_13),
.B2(n_252),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_250),
.C(n_256),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_284),
.B(n_273),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_282),
.Y(n_290)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_13),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_270),
.B(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_286),
.Y(n_293)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_271),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_291),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_266),
.C(n_276),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_293),
.C(n_290),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_278),
.B(n_280),
.Y(n_303)
);


endmodule