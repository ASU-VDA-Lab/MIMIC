module fake_jpeg_2722_n_697 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_697);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_697;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx3_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_62),
.Y(n_226)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_73),
.B(n_81),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_74),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_76),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_10),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_10),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_97),
.B(n_105),
.Y(n_164)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_27),
.B(n_7),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_116),
.Y(n_228)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_117),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_121),
.Y(n_234)
);

AND2x4_ASAP7_75t_SL g122 ( 
.A(n_55),
.B(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_125),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_55),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_28),
.Y(n_130)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_132),
.Y(n_231)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_32),
.B1(n_58),
.B2(n_31),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_136),
.A2(n_156),
.B1(n_159),
.B2(n_170),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_148),
.B(n_179),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_32),
.B1(n_42),
.B2(n_34),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_32),
.B1(n_58),
.B2(n_31),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_158),
.A2(n_217),
.B1(n_3),
.B2(n_4),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_55),
.B1(n_32),
.B2(n_34),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_57),
.C(n_50),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_5),
.C(n_17),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_50),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_168),
.B(n_176),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_63),
.A2(n_27),
.B1(n_54),
.B2(n_37),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_126),
.A2(n_55),
.B1(n_34),
.B2(n_41),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_172),
.A2(n_189),
.B1(n_193),
.B2(n_198),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_57),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_41),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_40),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_180),
.B(n_184),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_181),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_122),
.B(n_40),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_59),
.A2(n_49),
.B1(n_54),
.B2(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_49),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_209),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_133),
.A2(n_55),
.B1(n_42),
.B2(n_29),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_98),
.A2(n_37),
.B1(n_30),
.B2(n_29),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_12),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_206),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_91),
.A2(n_130),
.B1(n_76),
.B2(n_112),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_202),
.A2(n_204),
.B1(n_214),
.B2(n_225),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_67),
.A2(n_44),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_121),
.B(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_68),
.B(n_11),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_69),
.B(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_158),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_70),
.B(n_11),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_212),
.B(n_216),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_72),
.A2(n_44),
.B1(n_48),
.B2(n_25),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_80),
.B(n_7),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_89),
.A2(n_48),
.B1(n_56),
.B2(n_6),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_99),
.A2(n_48),
.B1(n_56),
.B2(n_6),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_0),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_104),
.A2(n_56),
.B1(n_6),
.B2(n_13),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_110),
.B(n_13),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_232),
.B(n_188),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_111),
.A2(n_5),
.B1(n_17),
.B2(n_15),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g354 ( 
.A(n_235),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_156),
.A2(n_75),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_236),
.A2(n_221),
.B1(n_191),
.B2(n_187),
.Y(n_325)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_237),
.Y(n_330)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_239),
.Y(n_348)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_240),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_162),
.A2(n_119),
.B1(n_6),
.B2(n_15),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_243),
.A2(n_251),
.B1(n_169),
.B2(n_226),
.Y(n_345)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_244),
.Y(n_333)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_245),
.Y(n_349)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_246),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_253),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_0),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_255),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_269),
.C(n_276),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_259),
.B(n_281),
.Y(n_342)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_261),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_164),
.B(n_0),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_262),
.B(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_267),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_137),
.B(n_0),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g383 ( 
.A(n_268),
.B(n_288),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_155),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_166),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_285),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_163),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_272),
.Y(n_355)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_174),
.Y(n_274)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_274),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_275),
.A2(n_277),
.B1(n_280),
.B2(n_307),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_186),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_146),
.A2(n_5),
.B1(n_15),
.B2(n_17),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_157),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_278),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_186),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_141),
.B(n_18),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_142),
.B(n_147),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_311),
.Y(n_326)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_284),
.A2(n_300),
.B1(n_318),
.B2(n_319),
.Y(n_344)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_166),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_286),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_220),
.A2(n_3),
.B1(n_4),
.B2(n_149),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_287),
.A2(n_290),
.B(n_172),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_145),
.B(n_3),
.Y(n_288)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_194),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_152),
.B(n_4),
.CI(n_153),
.CON(n_290),
.SN(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_295),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_223),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_293),
.B(n_296),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_183),
.B(n_229),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_298),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_192),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_157),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_299),
.Y(n_346)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_195),
.Y(n_298)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_201),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_135),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_302),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_175),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_303),
.B(n_309),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_177),
.B(n_222),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_197),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_306),
.B(n_310),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_219),
.A2(n_210),
.B1(n_213),
.B2(n_178),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_195),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_308),
.B(n_321),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_223),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_149),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_196),
.B(n_134),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_134),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_312),
.B(n_313),
.Y(n_381)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_139),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_196),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_314),
.B(n_317),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_139),
.A2(n_178),
.B1(n_203),
.B2(n_215),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_194),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_203),
.A2(n_204),
.B1(n_218),
.B2(n_221),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_185),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_215),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_214),
.A2(n_177),
.B1(n_187),
.B2(n_182),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_182),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_144),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_144),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_259),
.A2(n_202),
.B1(n_193),
.B2(n_233),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_323),
.A2(n_325),
.B1(n_340),
.B2(n_372),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_SL g390 ( 
.A1(n_334),
.A2(n_290),
.B(n_308),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_338),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_251),
.A2(n_159),
.B1(n_191),
.B2(n_169),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_345),
.A2(n_360),
.B1(n_367),
.B2(n_368),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_248),
.B(n_226),
.C(n_154),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_367),
.C(n_258),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_248),
.B(n_154),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_369),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_366),
.A2(n_284),
.B1(n_302),
.B2(n_306),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_279),
.B(n_194),
.C(n_201),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_262),
.B(n_201),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_279),
.A2(n_264),
.B(n_242),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_371),
.A2(n_378),
.B(n_303),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_251),
.A2(n_287),
.B1(n_280),
.B2(n_291),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_268),
.B(n_288),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_375),
.B(n_380),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_249),
.A2(n_254),
.B(n_273),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_257),
.A2(n_241),
.B1(n_236),
.B2(n_266),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_268),
.B(n_288),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_283),
.B(n_254),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_294),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_315),
.A2(n_311),
.B1(n_307),
.B2(n_290),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_386),
.A2(n_335),
.B1(n_342),
.B2(n_326),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_374),
.Y(n_438)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_390),
.A2(n_425),
.B(n_332),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_256),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_391),
.B(n_396),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_308),
.B(n_258),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_397),
.B(n_332),
.Y(n_457)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_395),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_370),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_323),
.A2(n_298),
.B(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_282),
.C(n_294),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_410),
.C(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_326),
.B(n_365),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_403),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_404),
.B(n_363),
.Y(n_464)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_379),
.A2(n_319),
.B1(n_260),
.B2(n_299),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_421),
.B1(n_426),
.B2(n_427),
.Y(n_441)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_238),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_297),
.B1(n_278),
.B2(n_321),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_412),
.A2(n_419),
.B(n_423),
.Y(n_442)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_295),
.C(n_247),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_416),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_350),
.B(n_252),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_417),
.B(n_337),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_437),
.B1(n_356),
.B2(n_355),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_434),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_327),
.A2(n_239),
.B1(n_301),
.B2(n_240),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_383),
.A2(n_235),
.B(n_274),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_424),
.A2(n_428),
.B1(n_429),
.B2(n_433),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_345),
.A2(n_271),
.B(n_246),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_325),
.A2(n_245),
.B1(n_250),
.B2(n_285),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_336),
.A2(n_267),
.B1(n_261),
.B2(n_271),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_300),
.B1(n_253),
.B2(n_289),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_340),
.A2(n_386),
.B1(n_360),
.B2(n_377),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_343),
.B(n_375),
.C(n_380),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_431),
.C(n_352),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_376),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_359),
.A2(n_368),
.B1(n_330),
.B2(n_333),
.Y(n_432)
);

AOI22x1_ASAP7_75t_L g467 ( 
.A1(n_432),
.A2(n_358),
.B1(n_348),
.B2(n_354),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_381),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_324),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_435),
.B(n_436),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_324),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_330),
.A2(n_352),
.B1(n_333),
.B2(n_374),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_468),
.C(n_471),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_388),
.B(n_356),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_461),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_443),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_437),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_472),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_451),
.A2(n_454),
.B1(n_463),
.B2(n_465),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_349),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_406),
.A2(n_346),
.B1(n_355),
.B2(n_344),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_467),
.Y(n_492)
);

AOI22x1_ASAP7_75t_SL g459 ( 
.A1(n_406),
.A2(n_341),
.B1(n_328),
.B2(n_363),
.Y(n_459)
);

AOI22x1_ASAP7_75t_SL g504 ( 
.A1(n_459),
.A2(n_426),
.B1(n_394),
.B2(n_341),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_339),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_400),
.A2(n_418),
.B1(n_403),
.B2(n_397),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_471),
.C(n_444),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_400),
.A2(n_348),
.B1(n_358),
.B2(n_324),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_331),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_392),
.B(n_331),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_475),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_351),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_432),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_392),
.B(n_351),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_403),
.A2(n_419),
.B1(n_393),
.B2(n_412),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_479),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_408),
.A2(n_348),
.B1(n_364),
.B2(n_349),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_328),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_472),
.A2(n_425),
.B1(n_416),
.B2(n_401),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_482),
.A2(n_447),
.B1(n_451),
.B2(n_465),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_423),
.B(n_415),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_484),
.A2(n_505),
.B(n_508),
.Y(n_544)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_487),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_443),
.A2(n_421),
.B(n_427),
.C(n_428),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_500),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_431),
.Y(n_490)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_490),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_387),
.C(n_399),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_491),
.B(n_493),
.C(n_510),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_404),
.C(n_422),
.Y(n_493)
);

A2O1A1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_420),
.B(n_422),
.C(n_434),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g552 ( 
.A1(n_495),
.A2(n_459),
.B(n_458),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_337),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_496),
.B(n_509),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_398),
.B1(n_409),
.B2(n_405),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_499),
.A2(n_504),
.B1(n_521),
.B2(n_441),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_456),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_501),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_402),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_502),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_456),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_512),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_442),
.A2(n_436),
.B(n_435),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_457),
.A2(n_478),
.B(n_447),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_473),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_440),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_469),
.Y(n_513)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_513),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_444),
.B(n_414),
.C(n_424),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_528)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_452),
.B(n_413),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_464),
.B(n_364),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_470),
.B(n_382),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_362),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_466),
.A2(n_439),
.B(n_467),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_519),
.A2(n_492),
.B(n_505),
.Y(n_538)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_474),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_454),
.A2(n_354),
.B1(n_407),
.B2(n_382),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_523),
.A2(n_524),
.B1(n_534),
.B2(n_538),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_498),
.A2(n_441),
.B1(n_439),
.B2(n_476),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_497),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_525),
.B(n_532),
.Y(n_563)
);

XOR2x2_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_476),
.Y(n_531)
);

XNOR2x1_ASAP7_75t_SL g575 ( 
.A(n_531),
.B(n_502),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_488),
.B(n_455),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_540),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_455),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_506),
.A2(n_473),
.B(n_462),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_481),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_542),
.B(n_553),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_545),
.B(n_483),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_506),
.A2(n_462),
.B(n_460),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_547),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_510),
.B(n_450),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_549),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_511),
.B(n_491),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_498),
.A2(n_450),
.B1(n_460),
.B2(n_479),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_550),
.A2(n_486),
.B1(n_502),
.B2(n_501),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_514),
.C(n_493),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_557),
.C(n_484),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_552),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_481),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_482),
.A2(n_492),
.B1(n_508),
.B2(n_513),
.Y(n_556)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_556),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_517),
.B(n_458),
.C(n_362),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_512),
.A2(n_503),
.B1(n_500),
.B2(n_504),
.Y(n_558)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_558),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_509),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_494),
.Y(n_567)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_564),
.B(n_566),
.C(n_571),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_551),
.B(n_527),
.C(n_528),
.Y(n_566)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_567),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_490),
.C(n_520),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_582),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_527),
.B(n_495),
.C(n_494),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_530),
.B(n_533),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_573),
.B(n_579),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_528),
.B(n_486),
.C(n_515),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_574),
.B(n_557),
.C(n_545),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_577),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_531),
.B(n_540),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_487),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_554),
.Y(n_580)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_580),
.Y(n_602)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_581),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_555),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_555),
.Y(n_583)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_583),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_584),
.A2(n_529),
.B1(n_556),
.B2(n_539),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_588),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_549),
.B(n_492),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_526),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_591),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_541),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_590),
.Y(n_595)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_526),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_522),
.B(n_548),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_535),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_562),
.A2(n_524),
.B1(n_546),
.B2(n_543),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_594),
.A2(n_611),
.B1(n_580),
.B2(n_536),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_599),
.B(n_601),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_566),
.B(n_544),
.C(n_547),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_563),
.Y(n_603)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_603),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_544),
.C(n_538),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_613),
.C(n_586),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_556),
.Y(n_605)
);

MAJx2_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_588),
.C(n_575),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_546),
.B(n_519),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_606),
.A2(n_609),
.B(n_617),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_543),
.B1(n_523),
.B2(n_550),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_608),
.A2(n_612),
.B1(n_587),
.B2(n_578),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_561),
.A2(n_556),
.B(n_521),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_568),
.A2(n_529),
.B1(n_483),
.B2(n_556),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_572),
.B(n_485),
.C(n_507),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_578),
.A2(n_489),
.B(n_560),
.Y(n_617)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_618),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_619),
.B(n_628),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_621),
.B(n_623),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_596),
.B(n_574),
.C(n_565),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_622),
.B(n_624),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_SL g623 ( 
.A(n_614),
.B(n_577),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_565),
.C(n_571),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_600),
.B(n_598),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_625),
.B(n_632),
.Y(n_644)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_626),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_600),
.Y(n_627)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_627),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_614),
.B(n_584),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_611),
.A2(n_591),
.B1(n_589),
.B2(n_587),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_630),
.A2(n_453),
.B1(n_354),
.B2(n_357),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_595),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_634),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_585),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_597),
.B(n_585),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_633),
.B(n_635),
.C(n_638),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_576),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_599),
.B(n_583),
.C(n_581),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_637),
.A2(n_612),
.B1(n_593),
.B2(n_602),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_601),
.B(n_449),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_604),
.B(n_453),
.C(n_449),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_639),
.B(n_605),
.C(n_616),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_630),
.A2(n_595),
.B(n_615),
.Y(n_643)
);

AO21x1_ASAP7_75t_L g669 ( 
.A1(n_643),
.A2(n_655),
.B(n_647),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_640),
.A2(n_610),
.B(n_606),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_646),
.B(n_648),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_647),
.B(n_654),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_626),
.A2(n_594),
.B1(n_615),
.B2(n_593),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_629),
.A2(n_617),
.B(n_608),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_650),
.B(n_628),
.Y(n_662)
);

FAx1_ASAP7_75t_SL g655 ( 
.A(n_619),
.B(n_597),
.CI(n_609),
.CON(n_655),
.SN(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_636),
.A2(n_602),
.B1(n_607),
.B2(n_616),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_656),
.A2(n_658),
.B1(n_629),
.B2(n_620),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_635),
.B(n_607),
.C(n_618),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_657),
.B(n_632),
.C(n_638),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_659),
.B(n_660),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_641),
.B(n_622),
.C(n_624),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_656),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_662),
.B(n_672),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_657),
.B(n_639),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_663),
.A2(n_664),
.B(n_665),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_642),
.B(n_631),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_642),
.B(n_621),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_649),
.A2(n_633),
.B1(n_623),
.B2(n_357),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_667),
.B(n_670),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_SL g668 ( 
.A(n_652),
.B(n_653),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_669),
.Y(n_681)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_644),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_654),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_660),
.B(n_651),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_676),
.B(n_677),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_672),
.B(n_645),
.C(n_653),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_666),
.B(n_648),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_678),
.B(n_682),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_671),
.A2(n_650),
.B(n_643),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_680),
.A2(n_669),
.B(n_662),
.Y(n_686)
);

XOR2xp5_ASAP7_75t_L g683 ( 
.A(n_677),
.B(n_668),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_684),
.Y(n_690)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_675),
.B(n_659),
.Y(n_684)
);

AOI21xp33_ASAP7_75t_L g689 ( 
.A1(n_686),
.A2(n_687),
.B(n_679),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_674),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_689),
.A2(n_691),
.B(n_687),
.Y(n_692)
);

A2O1A1O1Ixp25_ASAP7_75t_L g691 ( 
.A1(n_685),
.A2(n_674),
.B(n_673),
.C(n_681),
.D(n_682),
.Y(n_691)
);

MAJx2_ASAP7_75t_L g694 ( 
.A(n_692),
.B(n_693),
.C(n_666),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_690),
.B(n_688),
.C(n_681),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_694),
.A2(n_652),
.B(n_658),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_655),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_696),
.B(n_655),
.Y(n_697)
);


endmodule