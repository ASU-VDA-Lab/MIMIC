module fake_ariane_247_n_1133 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1133);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1133;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_931;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_608;
wire n_959;
wire n_494;
wire n_892;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_1025;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_54),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_113),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_37),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_164),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_107),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_112),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_66),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_127),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_188),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_19),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_43),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_99),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_28),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_130),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_35),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_45),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_96),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_124),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_68),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_179),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_10),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_63),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_26),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_57),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_77),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_136),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_118),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_154),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_111),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_74),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_133),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_123),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_52),
.Y(n_283)
);

BUFx2_ASAP7_75t_R g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_11),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_34),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_6),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_119),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_284),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_246),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_257),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_238),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_293),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_0),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_258),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_253),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_243),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_243),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_272),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_261),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_261),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_258),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_228),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_232),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_260),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_278),
.B1(n_285),
.B2(n_247),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_289),
.B1(n_277),
.B2(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_259),
.B(n_236),
.Y(n_351)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_222),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_341),
.Y(n_359)
);

CKINVDCx11_ASAP7_75t_R g360 ( 
.A(n_306),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_298),
.A2(n_274),
.B1(n_273),
.B2(n_223),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_312),
.B(n_226),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_294),
.B(n_236),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_236),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_298),
.A2(n_242),
.B1(n_265),
.B2(n_263),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_227),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

OAI22x1_ASAP7_75t_SL g377 ( 
.A1(n_306),
.A2(n_229),
.B1(n_231),
.B2(n_234),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_303),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_305),
.A2(n_237),
.B(n_235),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_302),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_295),
.B(n_239),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_295),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_315),
.B(n_259),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_299),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_299),
.A2(n_251),
.B1(n_241),
.B2(n_254),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_335),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

AO21x2_ASAP7_75t_L g403 ( 
.A1(n_349),
.A2(n_323),
.B(n_244),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_321),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_360),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_326),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_345),
.A2(n_332),
.B1(n_326),
.B2(n_296),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_397),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_352),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_240),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_352),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_393),
.B(n_332),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_352),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_397),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_384),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_384),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_334),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_343),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_384),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_386),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_386),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_386),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_386),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_386),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_394),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_396),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_377),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_361),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_395),
.B(n_334),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_259),
.Y(n_450)
);

BUFx6f_ASAP7_75t_SL g451 ( 
.A(n_345),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_387),
.B(n_250),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_395),
.B(n_252),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_374),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_389),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_348),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_390),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_390),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_364),
.B(n_30),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_388),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_R g463 ( 
.A(n_364),
.B(n_31),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_358),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_345),
.B(n_259),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_383),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_R g470 ( 
.A(n_364),
.B(n_32),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_382),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_372),
.Y(n_474)
);

BUFx4f_ASAP7_75t_L g475 ( 
.A(n_425),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_398),
.B(n_363),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_372),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_427),
.B(n_375),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_409),
.B(n_381),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_385),
.B1(n_365),
.B2(n_376),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_429),
.B(n_383),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_414),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_419),
.B(n_383),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_383),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_451),
.A2(n_385),
.B1(n_365),
.B2(n_376),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_428),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_415),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_435),
.B(n_366),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_413),
.B(n_366),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_367),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_366),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_436),
.B(n_366),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_450),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_413),
.B(n_366),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_378),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_462),
.B(n_385),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_451),
.B(n_458),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_448),
.B(n_368),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_454),
.B(n_365),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_405),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_454),
.B(n_365),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_439),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_471),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_370),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_440),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_401),
.B(n_404),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_411),
.B(n_362),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_432),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_365),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_422),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_420),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_467),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_443),
.B(n_379),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g541 ( 
.A(n_455),
.B(n_362),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_423),
.B(n_378),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_468),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_442),
.B(n_380),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_410),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_380),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_450),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_461),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_403),
.B(n_351),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_403),
.B(n_0),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_421),
.A2(n_270),
.B1(n_344),
.B2(n_347),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_472),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_520),
.B(n_535),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_491),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_547),
.A2(n_421),
.B1(n_444),
.B2(n_455),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_518),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_475),
.B(n_351),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_484),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_483),
.A2(n_344),
.B1(n_2),
.B2(n_3),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_540),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_463),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_477),
.B(n_470),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_521),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_353),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_544),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_1),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_512),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_542),
.B(n_353),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_507),
.A2(n_270),
.B1(n_6),
.B2(n_7),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_479),
.B(n_5),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_532),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_546),
.B(n_5),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_490),
.B(n_270),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_490),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_545),
.B(n_270),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

NAND3x1_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_9),
.C(n_11),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_539),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_497),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_510),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_542),
.B(n_540),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_505),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_519),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_523),
.B(n_12),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_517),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_543),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_529),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_517),
.B(n_13),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_538),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_552),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_514),
.Y(n_610)
);

AO22x2_ASAP7_75t_L g611 ( 
.A1(n_522),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_543),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_534),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_522),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_533),
.B(n_18),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_554),
.B(n_20),
.Y(n_617)
);

AO22x2_ASAP7_75t_L g618 ( 
.A1(n_533),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_523),
.B(n_21),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_492),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

O2A1O1Ixp5_ASAP7_75t_L g626 ( 
.A1(n_573),
.A2(n_555),
.B(n_550),
.C(n_511),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_557),
.B(n_492),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_523),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_587),
.B(n_526),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_571),
.A2(n_541),
.B(n_515),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_621),
.A2(n_622),
.B(n_565),
.Y(n_631)
);

AO21x1_ASAP7_75t_L g632 ( 
.A1(n_586),
.A2(n_551),
.B(n_502),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_556),
.A2(n_501),
.B1(n_537),
.B2(n_496),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_593),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_617),
.A2(n_494),
.B(n_480),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_621),
.A2(n_524),
.B(n_551),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_584),
.A2(n_501),
.B(n_614),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_482),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_623),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_601),
.B(n_605),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_591),
.A2(n_610),
.B(n_559),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_607),
.B(n_498),
.C(n_493),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_556),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_596),
.B(n_489),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_578),
.B(n_482),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_488),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_559),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_506),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_560),
.A2(n_500),
.B(n_489),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_486),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_596),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_570),
.A2(n_500),
.B(n_485),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_564),
.B(n_486),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_572),
.A2(n_485),
.B(n_478),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_566),
.B(n_486),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_612),
.B(n_543),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_574),
.A2(n_509),
.B1(n_485),
.B2(n_528),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_583),
.A2(n_509),
.B(n_478),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_580),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_585),
.B(n_486),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_589),
.A2(n_553),
.B1(n_528),
.B2(n_525),
.C(n_509),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_580),
.B(n_478),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_525),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_602),
.B(n_525),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_563),
.Y(n_665)
);

NOR2x1_ASAP7_75t_L g666 ( 
.A(n_579),
.B(n_528),
.Y(n_666)
);

OR2x4_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_22),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_602),
.B(n_549),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_619),
.B(n_562),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_582),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_558),
.A2(n_23),
.B(n_25),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_619),
.B(n_26),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_575),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_569),
.A2(n_36),
.B(n_33),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_581),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_609),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_622),
.A2(n_29),
.B(n_38),
.C(n_39),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_624),
.A2(n_40),
.B(n_42),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_562),
.B(n_44),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_620),
.A2(n_46),
.B(n_48),
.Y(n_680)
);

AOI33xp33_ASAP7_75t_L g681 ( 
.A1(n_603),
.A2(n_49),
.A3(n_50),
.B1(n_51),
.B2(n_53),
.B3(n_55),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_608),
.A2(n_56),
.B(n_58),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_600),
.A2(n_59),
.B(n_60),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_606),
.A2(n_61),
.B(n_62),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_581),
.A2(n_64),
.B(n_67),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_577),
.B(n_70),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_613),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_643),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_647),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_676),
.A2(n_670),
.B(n_629),
.C(n_633),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_634),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_638),
.B(n_604),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_640),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_628),
.B(n_588),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_675),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_628),
.B(n_594),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_645),
.A2(n_567),
.B(n_615),
.C(n_611),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_675),
.B(n_599),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_639),
.B(n_592),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_646),
.B(n_567),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_675),
.B(n_563),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_681),
.A2(n_618),
.B(n_615),
.C(n_611),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_672),
.A2(n_618),
.B1(n_589),
.B2(n_576),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_664),
.B(n_597),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_625),
.B(n_651),
.Y(n_705)
);

OAI21xp33_ASAP7_75t_L g706 ( 
.A1(n_671),
.A2(n_576),
.B(n_590),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_668),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_661),
.A2(n_590),
.B(n_76),
.C(n_78),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_R g709 ( 
.A(n_665),
.B(n_590),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_626),
.A2(n_590),
.B(n_79),
.C(n_80),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_625),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_659),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_659),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_625),
.B(n_75),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_630),
.A2(n_81),
.B(n_83),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_651),
.B(n_85),
.Y(n_716)
);

BUFx8_ASAP7_75t_L g717 ( 
.A(n_651),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_659),
.B(n_86),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_669),
.B(n_87),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_627),
.B(n_220),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_644),
.B(n_88),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_SL g722 ( 
.A1(n_637),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_656),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_639),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_679),
.A2(n_686),
.B1(n_667),
.B2(n_673),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_663),
.B(n_92),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_642),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.C(n_98),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_673),
.B(n_662),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_649),
.B(n_219),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_650),
.B(n_100),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_653),
.B(n_216),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_SL g735 ( 
.A1(n_682),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_636),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_677),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_631),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_657),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_655),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_660),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_654),
.B(n_108),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_685),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_635),
.A2(n_110),
.B(n_114),
.C(n_115),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_687),
.A2(n_116),
.B(n_117),
.C(n_120),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_658),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_717),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_712),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_712),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_691),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_721),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_724),
.B(n_632),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_739),
.B(n_652),
.Y(n_753)
);

BUFx4_ASAP7_75t_SL g754 ( 
.A(n_711),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_717),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_724),
.B(n_726),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_706),
.B(n_680),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_692),
.B(n_121),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_705),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_695),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_695),
.Y(n_761)
);

BUFx12f_ASAP7_75t_L g762 ( 
.A(n_716),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_713),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_696),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_688),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_689),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_713),
.B(n_701),
.Y(n_767)
);

BUFx12f_ASAP7_75t_L g768 ( 
.A(n_716),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_721),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_731),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_698),
.Y(n_771)
);

BUFx6f_ASAP7_75t_SL g772 ( 
.A(n_732),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_125),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_693),
.Y(n_775)
);

BUFx5_ASAP7_75t_L g776 ( 
.A(n_732),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_707),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_723),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_733),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_727),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_703),
.A2(n_684),
.B1(n_683),
.B2(n_674),
.Y(n_781)
);

INVx5_ASAP7_75t_L g782 ( 
.A(n_740),
.Y(n_782)
);

BUFx2_ASAP7_75t_R g783 ( 
.A(n_700),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_728),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_704),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_678),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_725),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_700),
.B(n_213),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_738),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_741),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_743),
.B(n_126),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_702),
.B(n_128),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_694),
.B(n_729),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_736),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_734),
.Y(n_796)
);

INVx6_ASAP7_75t_L g797 ( 
.A(n_699),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_719),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_720),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_742),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_746),
.B(n_708),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_714),
.B(n_129),
.Y(n_802)
);

INVx6_ASAP7_75t_SL g803 ( 
.A(n_718),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_690),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_715),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_737),
.B(n_212),
.Y(n_806)
);

NOR2x1_ASAP7_75t_R g807 ( 
.A(n_730),
.B(n_131),
.Y(n_807)
);

CKINVDCx6p67_ASAP7_75t_R g808 ( 
.A(n_722),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_744),
.B(n_132),
.Y(n_809)
);

INVx5_ASAP7_75t_SL g810 ( 
.A(n_735),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_745),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_804),
.A2(n_710),
.B(n_137),
.C(n_138),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_757),
.A2(n_134),
.B(n_139),
.Y(n_813)
);

AO32x2_ASAP7_75t_L g814 ( 
.A1(n_763),
.A2(n_140),
.A3(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_775),
.B(n_144),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_787),
.A2(n_145),
.B(n_146),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_757),
.A2(n_147),
.B(n_149),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_794),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_747),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_754),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_766),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_765),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_754),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_778),
.Y(n_824)
);

AO21x2_ASAP7_75t_L g825 ( 
.A1(n_789),
.A2(n_151),
.B(n_152),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_750),
.Y(n_826)
);

AO21x2_ASAP7_75t_L g827 ( 
.A1(n_789),
.A2(n_153),
.B(n_156),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_804),
.A2(n_157),
.B(n_158),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_777),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_781),
.A2(n_161),
.B(n_162),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_798),
.B(n_163),
.Y(n_832)
);

OA21x2_ASAP7_75t_L g833 ( 
.A1(n_787),
.A2(n_165),
.B(n_166),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_786),
.A2(n_167),
.B(n_168),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_795),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_772),
.A2(n_751),
.B1(n_774),
.B2(n_797),
.Y(n_836)
);

AOI222xp33_ASAP7_75t_SL g837 ( 
.A1(n_773),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.C1(n_174),
.C2(n_175),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_800),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_759),
.B(n_181),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_752),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_753),
.A2(n_182),
.B(n_183),
.C(n_184),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_781),
.A2(n_185),
.B(n_186),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_759),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_755),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_797),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_791),
.A2(n_189),
.B(n_190),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_764),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_811),
.A2(n_191),
.B(n_192),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_770),
.Y(n_849)
);

AO21x2_ASAP7_75t_L g850 ( 
.A1(n_791),
.A2(n_194),
.B(n_195),
.Y(n_850)
);

OAI21x1_ASAP7_75t_SL g851 ( 
.A1(n_749),
.A2(n_801),
.B(n_776),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_756),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_756),
.Y(n_853)
);

INVxp33_ASAP7_75t_L g854 ( 
.A(n_785),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_771),
.B(n_197),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_790),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_799),
.B(n_198),
.Y(n_857)
);

AO31x2_ASAP7_75t_L g858 ( 
.A1(n_786),
.A2(n_805),
.A3(n_808),
.B(n_810),
.Y(n_858)
);

OA21x2_ASAP7_75t_L g859 ( 
.A1(n_805),
.A2(n_203),
.B(n_204),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_809),
.A2(n_205),
.B(n_206),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_792),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_861)
);

AO21x2_ASAP7_75t_L g862 ( 
.A1(n_758),
.A2(n_211),
.B(n_810),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_771),
.B(n_785),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_810),
.A2(n_811),
.B(n_776),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_796),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_760),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_818),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_824),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_865),
.B(n_776),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_818),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_831),
.A2(n_788),
.B(n_776),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_865),
.B(n_776),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_824),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_861),
.A2(n_784),
.B1(n_788),
.B2(n_751),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_866),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_861),
.A2(n_788),
.B1(n_751),
.B2(n_769),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_858),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_826),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_864),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_821),
.Y(n_880)
);

INVx8_ASAP7_75t_L g881 ( 
.A(n_849),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_830),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_822),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_843),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_840),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_863),
.B(n_796),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_856),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_852),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_858),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_853),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_858),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_858),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_851),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_864),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_833),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_842),
.A2(n_817),
.B(n_813),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_864),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_833),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_833),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_859),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_866),
.B(n_769),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_816),
.A2(n_793),
.B(n_802),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_859),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_828),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_828),
.B(n_785),
.Y(n_905)
);

AOI21x1_ASAP7_75t_L g906 ( 
.A1(n_859),
.A2(n_806),
.B(n_811),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_825),
.Y(n_907)
);

CKINVDCx12_ASAP7_75t_R g908 ( 
.A(n_905),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_884),
.B(n_845),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_881),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_881),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_875),
.A2(n_823),
.B(n_820),
.C(n_847),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_884),
.B(n_854),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_874),
.A2(n_836),
.B1(n_860),
.B2(n_862),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_875),
.B(n_819),
.Y(n_915)
);

HB1xp67_ASAP7_75t_SL g916 ( 
.A(n_905),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_881),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_881),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_906),
.B(n_848),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_876),
.A2(n_836),
.B1(n_834),
.B2(n_838),
.Y(n_921)
);

NOR2x1p5_ASAP7_75t_L g922 ( 
.A(n_904),
.B(n_835),
.Y(n_922)
);

NAND2xp33_ASAP7_75t_R g923 ( 
.A(n_897),
.B(n_806),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_SL g924 ( 
.A(n_869),
.B(n_844),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_906),
.B(n_762),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_881),
.B(n_835),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_869),
.B(n_854),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_868),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_870),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_873),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_R g932 ( 
.A(n_897),
.B(n_806),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_872),
.B(n_904),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_904),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_872),
.B(n_862),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_885),
.B(n_839),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_900),
.A2(n_779),
.B1(n_768),
.B2(n_857),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_893),
.B(n_887),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_917),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_934),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_933),
.B(n_889),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_913),
.B(n_878),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_928),
.B(n_889),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_929),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_920),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_934),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_935),
.B(n_877),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_909),
.B(n_878),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_920),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_938),
.B(n_877),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_938),
.B(n_893),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_931),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_936),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_922),
.B(n_880),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_925),
.Y(n_955)
);

INVxp67_ASAP7_75t_R g956 ( 
.A(n_915),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_930),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_924),
.B(n_885),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_918),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_911),
.B(n_882),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_916),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_959),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_952),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_939),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_945),
.B(n_910),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_955),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_940),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_939),
.Y(n_968)
);

OAI211xp5_ASAP7_75t_L g969 ( 
.A1(n_945),
.A2(n_912),
.B(n_914),
.C(n_937),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_944),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_959),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_944),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_953),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_942),
.B(n_886),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_SL g975 ( 
.A1(n_961),
.A2(n_919),
.B(n_921),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_948),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_945),
.B(n_949),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_961),
.A2(n_912),
.B(n_914),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_973),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_973),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_971),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_966),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_969),
.B(n_932),
.C(n_923),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_964),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_976),
.B(n_958),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_966),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_965),
.B(n_945),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_965),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_968),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_970),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_965),
.B(n_956),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_981),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_991),
.B(n_956),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_979),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_962),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_991),
.B(n_975),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_980),
.B(n_963),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_984),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_985),
.B(n_974),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_983),
.A2(n_969),
.B1(n_837),
.B2(n_923),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_989),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_998),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_988),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_995),
.B(n_988),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_985),
.Y(n_1005)
);

NAND2x1_ASAP7_75t_SL g1006 ( 
.A(n_996),
.B(n_988),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_994),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1005),
.B(n_997),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1007),
.B(n_990),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1002),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1001),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1003),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_1004),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1006),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1006),
.B(n_1000),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_1006),
.B(n_987),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1005),
.A2(n_1000),
.B1(n_978),
.B2(n_993),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1003),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1008),
.B(n_972),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1015),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1009),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_1012),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1016),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1010),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1016),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1011),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1018),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1022),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1020),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_1023),
.B(n_1013),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1020),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1027),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1019),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_1017),
.B1(n_1014),
.B2(n_987),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1021),
.B(n_987),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1024),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_1026),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1029),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1028),
.B(n_967),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_967),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1032),
.B(n_943),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1035),
.B(n_982),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_1036),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1044),
.B(n_1037),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1044),
.B(n_1034),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_1038),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1040),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1041),
.B(n_977),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_1039),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_977),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1048),
.B(n_982),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_1046),
.B(n_977),
.Y(n_1054)
);

AOI211xp5_ASAP7_75t_SL g1055 ( 
.A1(n_1045),
.A2(n_857),
.B(n_832),
.C(n_841),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_1050),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1047),
.A2(n_986),
.B(n_954),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1049),
.B(n_986),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1045),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_1059),
.B(n_910),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1058),
.A2(n_945),
.B1(n_949),
.B2(n_812),
.C(n_829),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_1054),
.B(n_838),
.C(n_927),
.Y(n_1062)
);

AOI222xp33_ASAP7_75t_L g1063 ( 
.A1(n_1053),
.A2(n_949),
.B1(n_947),
.B2(n_898),
.C1(n_899),
.C2(n_895),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_949),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1057),
.A2(n_841),
.B(n_855),
.C(n_920),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1055),
.B1(n_949),
.B2(n_815),
.C(n_895),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1060),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_1062),
.A2(n_947),
.B1(n_958),
.B2(n_899),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1065),
.A2(n_937),
.B(n_941),
.C(n_898),
.Y(n_1069)
);

AOI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1061),
.A2(n_927),
.B(n_910),
.C(n_807),
.Y(n_1070)
);

OAI211xp5_ASAP7_75t_SL g1071 ( 
.A1(n_1063),
.A2(n_946),
.B(n_940),
.C(n_901),
.Y(n_1071)
);

OAI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1060),
.A2(n_946),
.B(n_940),
.C(n_910),
.Y(n_1072)
);

OAI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_1064),
.A2(n_932),
.B1(n_926),
.B2(n_802),
.C(n_946),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1064),
.A2(n_850),
.B(n_846),
.C(n_825),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1068),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_1067),
.A2(n_951),
.B(n_941),
.C(n_943),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1068),
.B(n_951),
.Y(n_1077)
);

OAI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1073),
.A2(n_1066),
.B1(n_1069),
.B2(n_1071),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1074),
.A2(n_803),
.B1(n_926),
.B2(n_907),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_1072),
.Y(n_1080)
);

OAI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1070),
.A2(n_926),
.B1(n_803),
.B2(n_894),
.Y(n_1081)
);

AOI221xp5_ASAP7_75t_L g1082 ( 
.A1(n_1066),
.A2(n_850),
.B1(n_846),
.B2(n_900),
.C(n_907),
.Y(n_1082)
);

OAI321xp33_ASAP7_75t_L g1083 ( 
.A1(n_1067),
.A2(n_767),
.A3(n_891),
.B1(n_950),
.B2(n_894),
.C(n_888),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1067),
.B(n_749),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_1080),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1075),
.B(n_950),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1084),
.B(n_748),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1077),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1076),
.B(n_960),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1078),
.B(n_748),
.Y(n_1090)
);

OAI221xp5_ASAP7_75t_L g1091 ( 
.A1(n_1082),
.A2(n_767),
.B1(n_879),
.B2(n_880),
.C(n_882),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1081),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1079),
.B(n_960),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1083),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_1080),
.B(n_780),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_1080),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1075),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1085),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_1088),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1096),
.A2(n_902),
.B(n_879),
.C(n_903),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1087),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1097),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1086),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1090),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1094),
.A2(n_827),
.B1(n_896),
.B2(n_894),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1095),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1099),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_SL g1108 ( 
.A1(n_1098),
.A2(n_1092),
.B(n_1091),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1104),
.A2(n_1089),
.B1(n_1093),
.B2(n_814),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1102),
.Y(n_1110)
);

XOR2x2_ASAP7_75t_L g1111 ( 
.A(n_1103),
.B(n_1089),
.Y(n_1111)
);

NOR4xp75_ASAP7_75t_SL g1112 ( 
.A(n_1101),
.B(n_1106),
.C(n_1105),
.D(n_1100),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1102),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_1110),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1107),
.A2(n_892),
.B1(n_891),
.B2(n_827),
.C(n_894),
.Y(n_1115)
);

AND4x1_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_814),
.C(n_890),
.D(n_888),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1114),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_1108),
.B1(n_1112),
.B2(n_1111),
.C(n_1115),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1118),
.A2(n_1109),
.B1(n_1116),
.B2(n_916),
.Y(n_1119)
);

NAND5xp2_ASAP7_75t_L g1120 ( 
.A(n_1119),
.B(n_793),
.C(n_814),
.D(n_783),
.E(n_807),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_814),
.B(n_879),
.C(n_903),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_955),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_902),
.B(n_871),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_R g1124 ( 
.A(n_1120),
.B(n_871),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1121),
.A2(n_894),
.B1(n_761),
.B2(n_780),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_780),
.B1(n_896),
.B2(n_761),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1123),
.A2(n_761),
.B1(n_871),
.B2(n_896),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1125),
.A2(n_896),
.B1(n_908),
.B2(n_871),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_783),
.B1(n_890),
.B2(n_782),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1127),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1128),
.A2(n_782),
.B(n_957),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_782),
.B(n_957),
.Y(n_1132)
);

AOI211xp5_ASAP7_75t_L g1133 ( 
.A1(n_1132),
.A2(n_1129),
.B(n_1131),
.C(n_883),
.Y(n_1133)
);


endmodule