module fake_aes_5154_n_31 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_2), .A2(n_8), .B(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
NAND3xp33_ASAP7_75t_L g21 ( .A(n_19), .B(n_16), .C(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_21), .B(n_17), .Y(n_25) );
AO22x2_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_16), .B1(n_15), .B2(n_18), .Y(n_26) );
OAI221xp5_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_13), .B1(n_1), .B2(n_2), .C(n_3), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_13), .Y(n_28) );
AO21x2_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_0), .B(n_4), .Y(n_29) );
NAND3xp33_ASAP7_75t_SL g30 ( .A(n_29), .B(n_27), .C(n_6), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_29), .B1(n_7), .B2(n_10), .Y(n_31) );
endmodule