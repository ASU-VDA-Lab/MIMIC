module fake_netlist_5_438_n_2127 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2127);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2127;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_116),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_16),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_62),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_114),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_97),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_73),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_44),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_80),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_74),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_109),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_74),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_57),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_56),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_49),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_118),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_14),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_83),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_176),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_152),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_192),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_34),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_76),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_68),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_159),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_110),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_101),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_128),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_87),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_70),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_44),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_81),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_66),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_28),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_93),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_34),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_71),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_82),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_172),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_132),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_162),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_148),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_42),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_23),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_122),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_29),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_188),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_190),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_77),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_135),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_61),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_29),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_158),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_111),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_54),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_9),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_96),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_65),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_160),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_100),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_21),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_85),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_69),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_75),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_98),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_121),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_149),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_46),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_38),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_63),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_168),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_103),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_45),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_187),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_70),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_179),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_136),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_115),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_22),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_89),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_163),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_182),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_45),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_99),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_126),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_16),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_14),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_119),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_38),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_51),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_18),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_154),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_47),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_26),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_41),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_169),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_138),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_76),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_24),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_107),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_33),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_189),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_78),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_191),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_24),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_130),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_4),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_31),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_43),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_86),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_129),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_13),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_58),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_65),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_17),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_54),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_27),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_94),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_153),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_33),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_112),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_43),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_134),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_0),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_5),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_39),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_72),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_177),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_175),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_9),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_72),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_145),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_36),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_142),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_52),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_36),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_21),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_62),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_61),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_40),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_31),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_32),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_228),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_283),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_239),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_283),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_201),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_208),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_241),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_269),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_200),
.B(n_0),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_199),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_201),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_202),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_283),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_203),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_283),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_272),
.B(n_2),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_272),
.B(n_2),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_283),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_283),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_274),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_302),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_252),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_302),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_302),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_236),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_252),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_302),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_330),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_360),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_302),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_205),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_200),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_200),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_206),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_207),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_213),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_243),
.B(n_3),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_215),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_305),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_232),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_233),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_258),
.B(n_3),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_230),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_242),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_245),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_248),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_267),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_375),
.B(n_4),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_267),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_305),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_267),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_281),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_254),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_255),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_281),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_281),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_256),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_349),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_214),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_257),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_216),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_262),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_214),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_349),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_306),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_335),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_349),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_265),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_229),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_229),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_263),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_335),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_310),
.B(n_5),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_235),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_310),
.B(n_8),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_264),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_222),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_275),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_249),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_345),
.B(n_8),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_249),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_279),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_270),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_270),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_384),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_278),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_393),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_403),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_405),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_345),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_407),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_465),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_469),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_394),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_411),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_435),
.B(n_333),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_476),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_425),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_428),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_429),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_396),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_416),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_481),
.B(n_277),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_434),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_R g539 ( 
.A(n_436),
.B(n_284),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_450),
.B(n_277),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_484),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_452),
.B(n_222),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_472),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_400),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_452),
.B(n_287),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_424),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_473),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_401),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_292),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_441),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_442),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_454),
.B(n_222),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_474),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_446),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_485),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_413),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_454),
.B(n_289),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_447),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_419),
.A2(n_314),
.B1(n_338),
.B2(n_342),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_448),
.Y(n_573)
);

HAxp5_ASAP7_75t_SL g574 ( 
.A(n_571),
.B(n_278),
.CON(n_574),
.SN(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_551),
.B(n_457),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_495),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_504),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_513),
.B(n_340),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_545),
.B(n_458),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_493),
.Y(n_581)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_499),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_495),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_544),
.B(n_456),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_518),
.B(n_461),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_503),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_541),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_515),
.Y(n_590)
);

INVx8_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_518),
.B(n_464),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_513),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_513),
.B(n_466),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_519),
.B(n_475),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_480),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_539),
.B(n_482),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_519),
.B(n_340),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_503),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_519),
.B(n_340),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_488),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_497),
.B(n_418),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_515),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_500),
.B(n_211),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_500),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_456),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_534),
.B(n_484),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_494),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_501),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_501),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_498),
.A2(n_445),
.B1(n_410),
.B2(n_409),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_502),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_534),
.B(n_491),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_509),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_527),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_504),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_506),
.B(n_491),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_539),
.B(n_443),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_527),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

AND2x2_ASAP7_75t_SL g628 ( 
.A(n_541),
.B(n_479),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_554),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_504),
.B(n_204),
.Y(n_630)
);

OA22x2_ASAP7_75t_L g631 ( 
.A1(n_500),
.A2(n_404),
.B1(n_398),
.B2(n_440),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_555),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_520),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_504),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_554),
.B(n_459),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_504),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_523),
.B(n_486),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_554),
.B(n_459),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_547),
.B(n_307),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_527),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_530),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_511),
.Y(n_643)
);

BUFx4f_ASAP7_75t_L g644 ( 
.A(n_511),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_460),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_547),
.B(n_324),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_511),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_402),
.B1(n_453),
.B2(n_313),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_569),
.B(n_211),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_556),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_536),
.A2(n_402),
.B1(n_313),
.B2(n_337),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_525),
.B(n_460),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_571),
.B(n_467),
.C(n_463),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_507),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_511),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_511),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_520),
.B(n_462),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_507),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_556),
.B(n_557),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_510),
.B(n_462),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_509),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_543),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_557),
.B(n_559),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g670 ( 
.A(n_528),
.B(n_422),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_512),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_512),
.B(n_468),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_516),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_538),
.B(n_552),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_559),
.B(n_468),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_516),
.B(n_471),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_517),
.B(n_471),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_537),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_517),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_514),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_548),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_537),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_560),
.B(n_561),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_561),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_521),
.B(n_489),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_548),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_537),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_564),
.B(n_430),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_548),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_522),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_505),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_521),
.B(n_198),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_508),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_528),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_508),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_526),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_546),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_553),
.A2(n_451),
.B1(n_251),
.B2(n_268),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_526),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_564),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_529),
.B(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_529),
.B(n_291),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_508),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_566),
.B(n_430),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_540),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_531),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_566),
.B(n_431),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_572),
.B(n_431),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_514),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_553),
.B(n_333),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_572),
.B(n_432),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_540),
.A2(n_211),
.B1(n_231),
.B2(n_225),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_532),
.B(n_297),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_532),
.B(n_298),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_508),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_505),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_533),
.B(n_535),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_533),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_535),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_565),
.B(n_333),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_565),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_710),
.B(n_570),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_710),
.B(n_570),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_618),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_591),
.B(n_505),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_704),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_704),
.Y(n_732)
);

NOR2x1p5_ASAP7_75t_L g733 ( 
.A(n_611),
.B(n_209),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_591),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_618),
.B(n_542),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_588),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_669),
.Y(n_737)
);

AND2x6_ASAP7_75t_SL g738 ( 
.A(n_605),
.B(n_286),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_629),
.B(n_542),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_640),
.B(n_210),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_629),
.B(n_537),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_585),
.A2(n_328),
.B1(n_304),
.B2(n_312),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_669),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_588),
.B(n_524),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_649),
.B(n_537),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_645),
.B(n_607),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_581),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_592),
.B(n_317),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_607),
.A2(n_326),
.B1(n_336),
.B2(n_344),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_645),
.B(n_204),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_685),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_575),
.B(n_212),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_609),
.B(n_217),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

NAND2x1_ASAP7_75t_L g758 ( 
.A(n_622),
.B(n_558),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_645),
.B(n_219),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_609),
.B(n_240),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_607),
.B(n_219),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_220),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_607),
.A2(n_355),
.B1(n_351),
.B2(n_359),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_656),
.B(n_221),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_688),
.B(n_524),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_653),
.A2(n_337),
.B1(n_386),
.B2(n_286),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_591),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_661),
.B(n_524),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_680),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_664),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_SL g771 ( 
.A(n_615),
.B(n_550),
.C(n_546),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_664),
.Y(n_772)
);

BUFx6f_ASAP7_75t_SL g773 ( 
.A(n_628),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_664),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_607),
.A2(n_628),
.B1(n_635),
.B2(n_610),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_593),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_636),
.A2(n_562),
.B(n_558),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_658),
.B(n_693),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_709),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_661),
.B(n_487),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_579),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_658),
.B(n_220),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_603),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_610),
.B(n_487),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_637),
.B(n_377),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_610),
.A2(n_381),
.B1(n_383),
.B2(n_322),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_696),
.B(n_623),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_624),
.B(n_223),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_693),
.B(n_226),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_694),
.B(n_226),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_620),
.B(n_218),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_694),
.B(n_237),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_593),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_591),
.B(n_550),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_603),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_587),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_451),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_635),
.A2(n_332),
.B1(n_260),
.B2(n_282),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_653),
.B(n_208),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_612),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_701),
.B(n_635),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_700),
.B(n_724),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_SL g803 ( 
.A(n_703),
.B(n_568),
.C(n_227),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_653),
.B(n_208),
.Y(n_804)
);

AO22x1_ASAP7_75t_L g805 ( 
.A1(n_582),
.A2(n_339),
.B1(n_341),
.B2(n_352),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_675),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_594),
.B(n_224),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_700),
.B(n_237),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_580),
.B(n_234),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

NOR2x1p5_ASAP7_75t_L g812 ( 
.A(n_611),
.B(n_250),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_701),
.B(n_240),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_724),
.B(n_238),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_626),
.B(n_238),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_627),
.B(n_244),
.Y(n_816)
);

NOR2x1_ASAP7_75t_L g817 ( 
.A(n_597),
.B(n_244),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_574),
.A2(n_333),
.B1(n_568),
.B2(n_218),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_715),
.B(n_725),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_701),
.B(n_240),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_721),
.B(n_339),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_632),
.B(n_259),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_648),
.B(n_247),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_654),
.B(n_686),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_687),
.B(n_705),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_680),
.B(n_240),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_584),
.B(n_240),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_612),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_SL g829 ( 
.A(n_617),
.B(n_652),
.C(n_657),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_653),
.A2(n_358),
.B1(n_341),
.B2(n_379),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_579),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_579),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_584),
.B(n_247),
.Y(n_833)
);

NOR3x1_ASAP7_75t_L g834 ( 
.A(n_620),
.B(n_354),
.C(n_352),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_695),
.B(n_84),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_617),
.B(n_266),
.C(n_261),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_709),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_638),
.B(n_253),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_674),
.B(n_354),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_638),
.B(n_490),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_595),
.B(n_240),
.Y(n_841)
);

AND2x6_ASAP7_75t_SL g842 ( 
.A(n_574),
.B(n_358),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_596),
.B(n_604),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_598),
.A2(n_288),
.B1(n_378),
.B2(n_372),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_631),
.B(n_253),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_633),
.B(n_218),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_613),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_712),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_613),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_614),
.B(n_260),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_680),
.B(n_208),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_644),
.A2(n_285),
.B(n_282),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_653),
.A2(n_379),
.B1(n_363),
.B2(n_389),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_614),
.B(n_285),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_616),
.B(n_288),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_619),
.B(n_90),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_670),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_707),
.B(n_271),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_680),
.B(n_208),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_631),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_616),
.B(n_639),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_639),
.B(n_301),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_718),
.B(n_276),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_662),
.B(n_301),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_662),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_712),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_663),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_670),
.B(n_363),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_631),
.B(n_303),
.Y(n_869)
);

AND2x6_ASAP7_75t_SL g870 ( 
.A(n_590),
.B(n_374),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_712),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_598),
.A2(n_348),
.B1(n_320),
.B2(n_322),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_619),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_713),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_663),
.B(n_303),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_713),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_691),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_719),
.B(n_280),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_671),
.B(n_311),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_653),
.A2(n_386),
.B1(n_389),
.B2(n_376),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_606),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_SL g883 ( 
.A1(n_587),
.A2(n_290),
.B1(n_294),
.B2(n_295),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_671),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_673),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_691),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_673),
.B(n_311),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_681),
.B(n_293),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_698),
.B(n_702),
.C(n_682),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_716),
.B(n_490),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_680),
.B(n_208),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_716),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_L g893 ( 
.A(n_681),
.B(n_208),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_717),
.A2(n_374),
.B1(n_376),
.B2(n_353),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_711),
.B(n_320),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_711),
.B(n_723),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_723),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_747),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_740),
.B(n_598),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_769),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_729),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_729),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_729),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_729),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_740),
.B(n_602),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_768),
.B(n_667),
.Y(n_907)
);

BUFx12f_ASAP7_75t_SL g908 ( 
.A(n_730),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_736),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_874),
.B(n_667),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_764),
.B(n_602),
.Y(n_911)
);

CKINVDCx11_ASAP7_75t_R g912 ( 
.A(n_868),
.Y(n_912)
);

AOI22x1_ASAP7_75t_L g913 ( 
.A1(n_748),
.A2(n_717),
.B1(n_602),
.B2(n_630),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_776),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_748),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_744),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_737),
.B(n_717),
.Y(n_917)
);

BUFx10_ASAP7_75t_L g918 ( 
.A(n_727),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_775),
.B(n_684),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_754),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_764),
.B(n_722),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_734),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_743),
.B(n_717),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

NOR2x1_ASAP7_75t_R g925 ( 
.A(n_767),
.B(n_682),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_772),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_769),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_754),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_771),
.B(n_714),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_727),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_756),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_756),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_746),
.B(n_684),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_807),
.B(n_706),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_794),
.B(n_714),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_783),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_726),
.B(n_225),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_SL g938 ( 
.A(n_726),
.B(n_218),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_752),
.B(n_655),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_829),
.A2(n_353),
.B1(n_225),
.B2(n_231),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_774),
.B(n_665),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_757),
.A2(n_353),
.B1(n_231),
.B2(n_316),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_783),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_807),
.B(n_825),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_819),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_795),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_776),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_825),
.B(n_647),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_769),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_779),
.B(n_684),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_745),
.A2(n_644),
.B(n_647),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_795),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_860),
.A2(n_316),
.B1(n_329),
.B2(n_370),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_821),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_819),
.A2(n_647),
.B1(n_622),
.B2(n_650),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_858),
.A2(n_622),
.B1(n_659),
.B2(n_650),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_811),
.B(n_672),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_753),
.B(n_818),
.C(n_788),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_821),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_837),
.B(n_676),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_803),
.B(n_299),
.C(n_296),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_800),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_848),
.B(n_677),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_793),
.B(n_578),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_728),
.B(n_650),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_800),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_828),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_779),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_793),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_730),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_866),
.B(n_659),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_866),
.Y(n_973)
);

OR2x2_ASAP7_75t_SL g974 ( 
.A(n_842),
.B(n_316),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_828),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_847),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_858),
.A2(n_622),
.B1(n_660),
.B2(n_659),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_796),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_847),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_849),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_849),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_787),
.B(n_684),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_865),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_781),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_821),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_730),
.B(n_630),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_882),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_863),
.B(n_578),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_865),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_867),
.Y(n_990)
);

BUFx8_ASAP7_75t_L g991 ( 
.A(n_773),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_867),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_863),
.B(n_578),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_879),
.B(n_578),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_831),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_879),
.B(n_578),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_886),
.B(n_589),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_878),
.B(n_630),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_832),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_765),
.Y(n_1002)
);

BUFx10_ASAP7_75t_L g1003 ( 
.A(n_809),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_897),
.B(n_589),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_885),
.B(n_684),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_796),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_885),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_731),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_731),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_732),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_784),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_780),
.B(n_492),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_732),
.Y(n_1013)
);

OR2x2_ASAP7_75t_SL g1014 ( 
.A(n_738),
.B(n_332),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_871),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_644),
.B(n_660),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_892),
.B(n_806),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_796),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_872),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_784),
.Y(n_1020)
);

BUFx8_ASAP7_75t_L g1021 ( 
.A(n_791),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_875),
.Y(n_1022)
);

CKINVDCx14_ASAP7_75t_R g1023 ( 
.A(n_797),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_877),
.B(n_348),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_778),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_846),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_801),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_839),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_801),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_840),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_810),
.B(n_576),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_802),
.B(n_690),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_840),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_861),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_R g1035 ( 
.A(n_797),
.B(n_300),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_857),
.A2(n_327),
.B1(n_308),
.B2(n_309),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_788),
.A2(n_660),
.B1(n_690),
.B2(n_608),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_890),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_845),
.B(n_318),
.C(n_315),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_753),
.B(n_589),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_869),
.B(n_321),
.C(n_319),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_890),
.B(n_576),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_896),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_824),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_L g1045 ( 
.A(n_852),
.B(n_690),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_888),
.B(n_589),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_888),
.B(n_589),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_741),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_839),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_755),
.B(n_608),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_856),
.B(n_367),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_735),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_755),
.B(n_739),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_870),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_839),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_835),
.B(n_367),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_761),
.A2(n_368),
.B(n_370),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_850),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_785),
.B(n_608),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_854),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_758),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_855),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_809),
.B(n_608),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_751),
.B(n_608),
.Y(n_1064)
);

AO22x1_ASAP7_75t_L g1065 ( 
.A1(n_834),
.A2(n_392),
.B1(n_323),
.B2(n_325),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_862),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_762),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_851),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_864),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_876),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_880),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_887),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_797),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_851),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_SL g1075 ( 
.A(n_883),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_759),
.B(n_833),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_859),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_895),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_893),
.B(n_331),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_782),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_815),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_816),
.Y(n_1082)
);

OR2x4_ASAP7_75t_L g1083 ( 
.A(n_822),
.B(n_492),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_838),
.Y(n_1084)
);

INVx3_ASAP7_75t_SL g1085 ( 
.A(n_749),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_789),
.B(n_634),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_894),
.B(n_577),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_817),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_823),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_822),
.B(n_790),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_792),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_943),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_913),
.A2(n_891),
.B(n_859),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1016),
.A2(n_891),
.B(n_841),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_944),
.B(n_808),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_921),
.B(n_814),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1034),
.B(n_1052),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_934),
.A2(n_760),
.B(n_777),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_911),
.A2(n_760),
.B(n_813),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_959),
.A2(n_836),
.B(n_827),
.C(n_733),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1002),
.B(n_812),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_973),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1005),
.A2(n_826),
.B(n_820),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_943),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_978),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1005),
.A2(n_826),
.B(n_820),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1045),
.A2(n_643),
.B(n_634),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_1043),
.A2(n_894),
.B(n_873),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_978),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_901),
.B(n_766),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1045),
.A2(n_643),
.B(n_634),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1043),
.B(n_742),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_986),
.B(n_805),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_916),
.B(n_889),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_909),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_937),
.A2(n_786),
.B1(n_750),
.B2(n_763),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_924),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_937),
.A2(n_844),
.B1(n_798),
.B2(n_799),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_901),
.B(n_813),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_952),
.A2(n_881),
.B(n_853),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_909),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1053),
.B(n_766),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_935),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_933),
.A2(n_881),
.B(n_853),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_987),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_899),
.A2(n_804),
.B(n_830),
.Y(n_1126)
);

INVx3_ASAP7_75t_SL g1127 ( 
.A(n_922),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_SL g1128 ( 
.A(n_924),
.B(n_690),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_973),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_906),
.A2(n_830),
.B(n_692),
.Y(n_1130)
);

OR2x6_ASAP7_75t_L g1131 ( 
.A(n_986),
.B(n_368),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1044),
.B(n_577),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_930),
.B(n_246),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1044),
.B(n_583),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_930),
.B(n_334),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_901),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1091),
.B(n_583),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_946),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_973),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_919),
.A2(n_601),
.B(n_641),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1040),
.A2(n_329),
.B1(n_378),
.B2(n_372),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_919),
.A2(n_599),
.B(n_621),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1032),
.A2(n_642),
.B(n_621),
.Y(n_1143)
);

AND3x4_ASAP7_75t_L g1144 ( 
.A(n_1055),
.B(n_273),
.C(n_246),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_946),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1006),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_SL g1147 ( 
.A1(n_982),
.A2(n_449),
.B(n_444),
.C(n_439),
.Y(n_1147)
);

AOI211x1_ASAP7_75t_L g1148 ( 
.A1(n_917),
.A2(n_432),
.B(n_444),
.C(n_439),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_924),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_988),
.A2(n_634),
.B(n_643),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1058),
.B(n_586),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_SL g1152 ( 
.A1(n_914),
.A2(n_625),
.B(n_692),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1060),
.B(n_586),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1032),
.A2(n_965),
.B(n_1064),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_963),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_940),
.A2(n_599),
.B(n_641),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_922),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1062),
.B(n_601),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_938),
.A2(n_357),
.B(n_346),
.C(n_347),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1066),
.B(n_625),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_986),
.B(n_690),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_993),
.A2(n_634),
.B(n_643),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_907),
.B(n_1026),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_907),
.B(n_433),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_901),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1012),
.B(n_433),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1013),
.A2(n_646),
.B(n_642),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1063),
.A2(n_689),
.A3(n_651),
.B(n_646),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1027),
.A2(n_683),
.B(n_668),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_905),
.Y(n_1170)
);

BUFx2_ASAP7_75t_R g1171 ( 
.A(n_971),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1013),
.A2(n_651),
.B(n_666),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1013),
.A2(n_666),
.B(n_668),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_933),
.A2(n_689),
.B(n_683),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1004),
.A2(n_679),
.B(n_562),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_939),
.A2(n_388),
.B(n_350),
.C(n_356),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1029),
.A2(n_679),
.B(n_708),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1090),
.B(n_643),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_995),
.A2(n_678),
.B(n_708),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1050),
.A2(n_563),
.B(n_558),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1072),
.B(n_678),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_910),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_972),
.A2(n_563),
.B(n_567),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1039),
.B(n_387),
.C(n_361),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1048),
.A2(n_720),
.B(n_708),
.Y(n_1185)
);

AO32x2_ASAP7_75t_L g1186 ( 
.A1(n_914),
.A2(n_246),
.A3(n_273),
.B1(n_12),
.B2(n_13),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1046),
.A2(n_437),
.A3(n_438),
.B(n_449),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1047),
.A2(n_437),
.A3(n_438),
.B(n_562),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1025),
.B(n_678),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_963),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1084),
.B(n_678),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_997),
.A2(n_1086),
.B(n_966),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_982),
.A2(n_563),
.B(n_567),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_924),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_975),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_L g1196 ( 
.A(n_902),
.B(n_678),
.Y(n_1196)
);

BUFx4f_ASAP7_75t_SL g1197 ( 
.A(n_1006),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1059),
.A2(n_720),
.B(n_708),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_939),
.A2(n_373),
.B(n_364),
.C(n_365),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_948),
.A2(n_720),
.B(n_708),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_975),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1048),
.A2(n_720),
.B(n_699),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1084),
.B(n_366),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1084),
.B(n_369),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1081),
.B(n_371),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_972),
.A2(n_567),
.B(n_208),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1017),
.A2(n_385),
.B(n_380),
.C(n_391),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_951),
.A2(n_208),
.B(n_699),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_924),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1017),
.A2(n_273),
.B(n_246),
.C(n_697),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_980),
.A2(n_141),
.B(n_95),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_905),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_999),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1041),
.B(n_720),
.C(n_699),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_898),
.A2(n_699),
.B(n_697),
.Y(n_1215)
);

INVx5_ASAP7_75t_L g1216 ( 
.A(n_905),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_980),
.A2(n_140),
.B(n_102),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_947),
.A2(n_1076),
.B1(n_1070),
.B2(n_1071),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_985),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1012),
.B(n_918),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1089),
.B(n_1081),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_980),
.A2(n_156),
.B(n_108),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_947),
.A2(n_1076),
.B1(n_1070),
.B2(n_1078),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1069),
.A2(n_699),
.B(n_697),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1076),
.A2(n_697),
.B1(n_157),
.B2(n_181),
.Y(n_1225)
);

AO32x2_ASAP7_75t_L g1226 ( 
.A1(n_900),
.A2(n_273),
.A3(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1089),
.B(n_697),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1082),
.B(n_10),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_945),
.B(n_10),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_918),
.B(n_1038),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1069),
.A2(n_180),
.B(n_178),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_981),
.A2(n_990),
.B(n_989),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1082),
.B(n_11),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_950),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1071),
.B(n_15),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_L g1236 ( 
.A(n_1011),
.Y(n_1236)
);

AOI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1030),
.A2(n_17),
.B(n_18),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1021),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_989),
.A2(n_19),
.A3(n_20),
.B(n_23),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1030),
.A2(n_1033),
.B1(n_1038),
.B2(n_1003),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_981),
.A2(n_170),
.B(n_167),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1076),
.A2(n_161),
.B1(n_137),
.B2(n_133),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1020),
.B(n_926),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_990),
.A2(n_20),
.A3(n_25),
.B(n_26),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_918),
.B(n_25),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1068),
.B(n_131),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1033),
.B(n_27),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_981),
.A2(n_127),
.B(n_124),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1000),
.A2(n_123),
.B(n_91),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1000),
.A2(n_30),
.B(n_32),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_904),
.A2(n_30),
.B(n_35),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_951),
.A2(n_37),
.B(n_40),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1078),
.B(n_37),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1037),
.A2(n_46),
.B(n_48),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_915),
.A2(n_50),
.A3(n_51),
.B(n_52),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_920),
.A2(n_50),
.B(n_53),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1232),
.A2(n_1007),
.B(n_931),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1232),
.A2(n_928),
.B(n_953),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1122),
.B(n_1213),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1097),
.B(n_1221),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1238),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1220),
.B(n_1003),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1120),
.A2(n_962),
.B(n_1087),
.C(n_1049),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1105),
.Y(n_1266)
);

AND2x2_ASAP7_75t_SL g1267 ( 
.A(n_1110),
.B(n_905),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1192),
.A2(n_983),
.B(n_994),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1104),
.B(n_917),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1193),
.A2(n_979),
.B(n_936),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1135),
.A2(n_1003),
.B1(n_1055),
.B2(n_1075),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1159),
.B(n_1135),
.C(n_1100),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1104),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1175),
.A2(n_968),
.B(n_932),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1177),
.A2(n_1057),
.B(n_957),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1243),
.B(n_926),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_976),
.B(n_992),
.Y(n_1277)
);

BUFx2_ASAP7_75t_SL g1278 ( 
.A(n_1125),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1102),
.B(n_902),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1145),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1101),
.A2(n_1035),
.B1(n_1023),
.B2(n_1073),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_L g1282 ( 
.A(n_1157),
.B(n_1115),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1138),
.B(n_923),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1195),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1163),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1180),
.A2(n_967),
.B(n_1008),
.Y(n_1286)
);

AOI221xp5_ASAP7_75t_L g1287 ( 
.A1(n_1176),
.A2(n_929),
.B1(n_1075),
.B2(n_1028),
.C(n_1065),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1085),
.B(n_960),
.C(n_955),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1194),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1138),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1126),
.A2(n_1057),
.B(n_977),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1166),
.B(n_1015),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1099),
.A2(n_1057),
.B(n_956),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1243),
.B(n_926),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1149),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1236),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1205),
.B(n_945),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1157),
.B(n_925),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1105),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1155),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1112),
.B(n_945),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1094),
.A2(n_1008),
.B(n_1010),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1155),
.B(n_923),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1250),
.A2(n_942),
.B(n_1009),
.Y(n_1304)
);

NAND3x1_ASAP7_75t_L g1305 ( 
.A(n_1229),
.B(n_1075),
.C(n_908),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1201),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1130),
.A2(n_998),
.B(n_999),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1243),
.B(n_1020),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1190),
.B(n_1042),
.Y(n_1309)
);

AO21x2_ASAP7_75t_L g1310 ( 
.A1(n_1185),
.A2(n_1024),
.B(n_1022),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1167),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1163),
.B(n_1080),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1123),
.A2(n_1049),
.B1(n_1073),
.B2(n_1083),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1094),
.A2(n_969),
.B(n_949),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1250),
.A2(n_1022),
.B(n_1015),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1137),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1116),
.A2(n_1049),
.B1(n_970),
.B2(n_1020),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1133),
.B(n_1080),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1174),
.A2(n_1143),
.B(n_1172),
.Y(n_1319)
);

AOI222xp33_ASAP7_75t_L g1320 ( 
.A1(n_1114),
.A2(n_912),
.B1(n_1021),
.B2(n_1054),
.C1(n_985),
.C2(n_991),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1102),
.B(n_903),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1173),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1174),
.A2(n_969),
.B(n_949),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1247),
.B(n_1042),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1182),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1150),
.A2(n_1056),
.B(n_1031),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1093),
.A2(n_969),
.B(n_949),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1218),
.A2(n_1019),
.B(n_927),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1176),
.A2(n_1085),
.B(n_1056),
.C(n_1051),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1164),
.B(n_1019),
.Y(n_1330)
);

INVx8_ASAP7_75t_L g1331 ( 
.A(n_1117),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1156),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1093),
.A2(n_1061),
.B(n_1031),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1098),
.A2(n_1024),
.B(n_954),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1117),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1223),
.A2(n_941),
.B(n_961),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1219),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1121),
.B(n_1083),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1109),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1162),
.A2(n_1061),
.B(n_1067),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1109),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1151),
.Y(n_1342)
);

BUFx2_ASAP7_75t_SL g1343 ( 
.A(n_1146),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1141),
.A2(n_1088),
.A3(n_927),
.B(n_900),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1153),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1161),
.B(n_986),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1158),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1160),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1156),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1107),
.A2(n_1024),
.B(n_1079),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1111),
.A2(n_1067),
.B(n_1056),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1129),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1249),
.A2(n_1067),
.B(n_1056),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1249),
.A2(n_1067),
.B(n_927),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1229),
.A2(n_1011),
.B1(n_1023),
.B2(n_1049),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1132),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1113),
.A2(n_1021),
.B1(n_1049),
.B2(n_1011),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1113),
.A2(n_1011),
.B1(n_958),
.B2(n_964),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1206),
.A2(n_900),
.B(n_1077),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1199),
.B(n_958),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1211),
.A2(n_1077),
.B(n_1068),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1211),
.A2(n_1077),
.B(n_1068),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1134),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1245),
.B(n_958),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1235),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1129),
.B(n_903),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1253),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1199),
.A2(n_1051),
.B(n_1088),
.C(n_1018),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1203),
.B(n_961),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1217),
.A2(n_1077),
.B(n_1068),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1113),
.A2(n_961),
.B1(n_964),
.B2(n_941),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1139),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1110),
.A2(n_1051),
.B(n_970),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_SL g1375 ( 
.A1(n_1246),
.A2(n_1051),
.B(n_974),
.C(n_1014),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1233),
.B(n_964),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1121),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1148),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1120),
.A2(n_941),
.B(n_1036),
.C(n_970),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1181),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1184),
.A2(n_984),
.B1(n_1001),
.B2(n_996),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1217),
.A2(n_1001),
.B(n_996),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1251),
.A2(n_974),
.A3(n_1014),
.B(n_970),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1165),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1194),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1127),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1210),
.A2(n_1001),
.A3(n_996),
.B(n_57),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1146),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1117),
.B(n_1001),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1222),
.A2(n_1001),
.B(n_996),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1161),
.B(n_1018),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1222),
.A2(n_996),
.B(n_984),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1241),
.A2(n_984),
.B(n_908),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1117),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1171),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1165),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1118),
.A2(n_984),
.B1(n_971),
.B2(n_1054),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1216),
.B(n_950),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1216),
.B(n_950),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1230),
.B(n_991),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1170),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1207),
.A2(n_991),
.B1(n_912),
.B2(n_58),
.C(n_59),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1241),
.A2(n_53),
.B(n_55),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1127),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1248),
.A2(n_60),
.B(n_67),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1248),
.A2(n_67),
.B(n_71),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1210),
.A2(n_75),
.A3(n_77),
.B(n_78),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1189),
.A2(n_79),
.B(n_1178),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1183),
.A2(n_79),
.B(n_1215),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1124),
.A2(n_1204),
.B(n_1227),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1168),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1124),
.A2(n_1103),
.B(n_1106),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1168),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1179),
.A2(n_1202),
.B(n_1224),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1216),
.B(n_1246),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1131),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1194),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1161),
.B(n_1240),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1140),
.A2(n_1142),
.B(n_1208),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1147),
.A2(n_1152),
.B(n_1169),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1252),
.A2(n_1191),
.B(n_1200),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1252),
.A2(n_1254),
.B(n_1231),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1198),
.A2(n_1119),
.B(n_1196),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1168),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1170),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1212),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1364),
.B(n_1207),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1257),
.A2(n_1285),
.B1(n_1312),
.B2(n_1355),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1402),
.A2(n_1272),
.B1(n_1404),
.B2(n_1237),
.C(n_1375),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1258),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1386),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1331),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1273),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1280),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1310),
.A2(n_1178),
.B(n_1149),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1331),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1257),
.A2(n_1144),
.B1(n_1197),
.B2(n_1131),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1386),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1364),
.B(n_1324),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1318),
.B(n_1144),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1263),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1375),
.A2(n_1242),
.B1(n_1225),
.B2(n_1108),
.C(n_1238),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1271),
.A2(n_1197),
.B1(n_1131),
.B2(n_1236),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1337),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1412),
.A2(n_1214),
.B(n_1187),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1284),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1306),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1273),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1397),
.A2(n_1234),
.B1(n_1256),
.B2(n_1186),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1290),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1263),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1276),
.B(n_1136),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1276),
.B(n_1136),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1278),
.Y(n_1454)
);

OAI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1287),
.A2(n_1119),
.B1(n_1256),
.B2(n_1212),
.C(n_1216),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1295),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1266),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1266),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1365),
.A2(n_1256),
.B1(n_1234),
.B2(n_1186),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1290),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1325),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1300),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1324),
.B(n_1186),
.Y(n_1463)
);

INVxp33_ASAP7_75t_SL g1464 ( 
.A(n_1298),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1331),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1262),
.B(n_1194),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1300),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1297),
.A2(n_1209),
.B1(n_1186),
.B2(n_1226),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1276),
.B(n_1209),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1262),
.B(n_1209),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1367),
.A2(n_1226),
.B1(n_1209),
.B2(n_1255),
.Y(n_1471)
);

O2A1O1Ixp5_ASAP7_75t_L g1472 ( 
.A1(n_1301),
.A2(n_1226),
.B(n_1187),
.C(n_1188),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1269),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1338),
.B(n_1255),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1299),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1337),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1294),
.B(n_1128),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1294),
.B(n_1168),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1377),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1371),
.A2(n_1226),
.B1(n_1255),
.B2(n_1239),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1261),
.A2(n_1255),
.B1(n_1239),
.B2(n_1244),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1267),
.A2(n_1239),
.B1(n_1244),
.B2(n_1187),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1330),
.B(n_1239),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1269),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1408),
.A2(n_1188),
.B(n_1187),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1294),
.B(n_1188),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1329),
.A2(n_1188),
.B(n_1244),
.C(n_1368),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1330),
.B(n_1244),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1308),
.B(n_1346),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1292),
.B(n_1309),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1264),
.B2(n_1357),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1261),
.A2(n_1292),
.B1(n_1376),
.B2(n_1369),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1376),
.B(n_1360),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1283),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1281),
.A2(n_1313),
.B1(n_1305),
.B2(n_1418),
.Y(n_1495)
);

AOI21xp33_ASAP7_75t_L g1496 ( 
.A1(n_1288),
.A2(n_1301),
.B(n_1336),
.Y(n_1496)
);

NAND2x1p5_ASAP7_75t_L g1497 ( 
.A(n_1335),
.B(n_1394),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1283),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1267),
.A2(n_1346),
.B1(n_1305),
.B2(n_1391),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1346),
.A2(n_1391),
.B1(n_1381),
.B2(n_1416),
.Y(n_1500)
);

BUFx12f_ASAP7_75t_L g1501 ( 
.A(n_1400),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1303),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1331),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1382),
.A2(n_1390),
.B(n_1392),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1316),
.B(n_1342),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1347),
.B2(n_1363),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1317),
.A2(n_1374),
.B(n_1394),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1356),
.B(n_1309),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1308),
.B(n_1299),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1418),
.B(n_1303),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1315),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1380),
.B(n_1308),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1384),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1310),
.A2(n_1334),
.B(n_1291),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1346),
.A2(n_1391),
.B1(n_1378),
.B2(n_1282),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1379),
.A2(n_1265),
.B(n_1403),
.C(n_1406),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1339),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1339),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1418),
.A2(n_1400),
.B1(n_1343),
.B2(n_1415),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1426),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1382),
.A2(n_1390),
.B(n_1392),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1335),
.A2(n_1394),
.B(n_1389),
.Y(n_1522)
);

AOI21xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1320),
.A2(n_1395),
.B(n_1399),
.Y(n_1523)
);

OAI222xp33_ASAP7_75t_L g1524 ( 
.A1(n_1391),
.A2(n_1398),
.B1(n_1399),
.B2(n_1415),
.C1(n_1400),
.C2(n_1296),
.Y(n_1524)
);

CKINVDCx6p67_ASAP7_75t_R g1525 ( 
.A(n_1341),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1396),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1425),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1383),
.B(n_1341),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1315),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1319),
.A2(n_1353),
.B(n_1286),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1401),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1388),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1398),
.A2(n_1399),
.B1(n_1388),
.B2(n_1296),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1315),
.Y(n_1534)
);

OAI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1379),
.A2(n_1265),
.B1(n_1410),
.B2(n_1415),
.C(n_1398),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1328),
.B(n_1279),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1332),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1417),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1383),
.B(n_1407),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1335),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1291),
.A2(n_1307),
.B1(n_1334),
.B2(n_1293),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1291),
.A2(n_1307),
.B1(n_1334),
.B2(n_1293),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1383),
.B(n_1407),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1344),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1307),
.A2(n_1293),
.B1(n_1422),
.B2(n_1328),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1417),
.B(n_1279),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1289),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1289),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1352),
.A2(n_1373),
.B1(n_1424),
.B2(n_1411),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1417),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1289),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1407),
.B(n_1387),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1422),
.A2(n_1424),
.B1(n_1413),
.B2(n_1411),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1352),
.B(n_1373),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1373),
.B(n_1289),
.Y(n_1555)
);

CKINVDCx11_ASAP7_75t_R g1556 ( 
.A(n_1289),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1385),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1407),
.B(n_1387),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1422),
.A2(n_1413),
.B1(n_1310),
.B2(n_1275),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1279),
.B(n_1366),
.C(n_1321),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1275),
.A2(n_1350),
.B1(n_1268),
.B2(n_1406),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1350),
.A2(n_1403),
.B1(n_1405),
.B2(n_1275),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1389),
.A2(n_1321),
.B1(n_1366),
.B2(n_1268),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1321),
.A2(n_1366),
.B1(n_1389),
.B2(n_1349),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1385),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1319),
.A2(n_1353),
.B(n_1286),
.Y(n_1566)
);

BUFx4f_ASAP7_75t_SL g1567 ( 
.A(n_1385),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1421),
.A2(n_1333),
.B(n_1419),
.Y(n_1568)
);

OR2x6_ASAP7_75t_L g1569 ( 
.A(n_1351),
.B(n_1359),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1350),
.A2(n_1405),
.B1(n_1351),
.B2(n_1393),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1385),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1387),
.B(n_1385),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1349),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1387),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1387),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1302),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1268),
.A2(n_1326),
.B1(n_1304),
.B2(n_1322),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_R g1578 ( 
.A(n_1304),
.B(n_1393),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1259),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1326),
.A2(n_1304),
.B1(n_1311),
.B2(n_1322),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1302),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1259),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1344),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1260),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1407),
.A2(n_1311),
.B1(n_1344),
.B2(n_1277),
.C(n_1421),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1260),
.Y(n_1586)
);

AOI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1277),
.A2(n_1340),
.B(n_1420),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_SL g1588 ( 
.A(n_1361),
.B(n_1370),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1270),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1344),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1344),
.B(n_1340),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1511),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1532),
.Y(n_1593)
);

AOI222xp33_ASAP7_75t_L g1594 ( 
.A1(n_1429),
.A2(n_1333),
.B1(n_1270),
.B2(n_1274),
.C1(n_1361),
.C2(n_1370),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1463),
.B(n_1327),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1314),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1539),
.B(n_1327),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1496),
.A2(n_1440),
.B1(n_1428),
.B2(n_1437),
.C(n_1523),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1440),
.A2(n_1274),
.B1(n_1414),
.B2(n_1423),
.C(n_1362),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1491),
.A2(n_1362),
.B1(n_1354),
.B2(n_1423),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1427),
.A2(n_1354),
.B1(n_1409),
.B2(n_1419),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1478),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1489),
.B(n_1359),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1505),
.B(n_1323),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1493),
.A2(n_1409),
.B1(n_1420),
.B2(n_1323),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1493),
.A2(n_1414),
.B1(n_1442),
.B2(n_1474),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1492),
.A2(n_1500),
.B1(n_1499),
.B2(n_1489),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1492),
.A2(n_1489),
.B1(n_1439),
.B2(n_1486),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1434),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1446),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1486),
.B(n_1478),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1543),
.B(n_1552),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1486),
.A2(n_1510),
.B1(n_1495),
.B2(n_1501),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1443),
.A2(n_1464),
.B1(n_1461),
.B2(n_1501),
.Y(n_1614)
);

OAI211xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1479),
.A2(n_1454),
.B(n_1506),
.C(n_1449),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1432),
.Y(n_1616)
);

OAI211xp5_ASAP7_75t_L g1617 ( 
.A1(n_1506),
.A2(n_1459),
.B(n_1468),
.C(n_1505),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1558),
.A2(n_1459),
.B1(n_1535),
.B2(n_1487),
.C(n_1471),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1510),
.A2(n_1519),
.B1(n_1528),
.B2(n_1444),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1483),
.B(n_1574),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1533),
.A2(n_1484),
.B1(n_1502),
.B2(n_1494),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1487),
.B(n_1516),
.C(n_1562),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1507),
.B(n_1536),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1516),
.A2(n_1514),
.B(n_1585),
.Y(n_1625)
);

OAI22x1_ASAP7_75t_L g1626 ( 
.A1(n_1575),
.A2(n_1544),
.B1(n_1583),
.B2(n_1456),
.Y(n_1626)
);

BUFx4f_ASAP7_75t_SL g1627 ( 
.A(n_1532),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1476),
.B(n_1438),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1455),
.A2(n_1470),
.B(n_1488),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1485),
.A2(n_1512),
.B1(n_1508),
.B2(n_1470),
.C(n_1518),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1466),
.B(n_1473),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1431),
.A2(n_1525),
.B1(n_1457),
.B2(n_1517),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1569),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1590),
.A2(n_1431),
.B1(n_1475),
.B2(n_1567),
.Y(n_1634)
);

OAI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1541),
.A2(n_1542),
.B(n_1471),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1498),
.A2(n_1515),
.B1(n_1509),
.B2(n_1590),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1515),
.A2(n_1509),
.B1(n_1453),
.B2(n_1452),
.Y(n_1637)
);

NAND2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1432),
.B(n_1465),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1452),
.A2(n_1453),
.B1(n_1477),
.B2(n_1536),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1475),
.A2(n_1567),
.B1(n_1456),
.B2(n_1477),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1441),
.A2(n_1451),
.B1(n_1458),
.B2(n_1469),
.Y(n_1641)
);

AOI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1524),
.A2(n_1560),
.B(n_1564),
.C(n_1447),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1536),
.A2(n_1480),
.B1(n_1546),
.B2(n_1469),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1541),
.A2(n_1542),
.B1(n_1480),
.B2(n_1545),
.C(n_1481),
.Y(n_1644)
);

AOI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1445),
.A2(n_1545),
.B(n_1554),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1513),
.A2(n_1531),
.B1(n_1520),
.B2(n_1526),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1450),
.B(n_1467),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1527),
.A2(n_1564),
.B1(n_1563),
.B2(n_1544),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1432),
.A2(n_1465),
.B1(n_1503),
.B2(n_1540),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1497),
.A2(n_1436),
.B1(n_1482),
.B2(n_1550),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1591),
.B(n_1583),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1432),
.A2(n_1465),
.B1(n_1436),
.B2(n_1538),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1460),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1548),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1556),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1465),
.A2(n_1565),
.B1(n_1547),
.B2(n_1571),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1561),
.A2(n_1559),
.B(n_1570),
.C(n_1435),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1433),
.B(n_1448),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1556),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1551),
.A2(n_1462),
.B1(n_1540),
.B2(n_1548),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1472),
.A2(n_1559),
.B1(n_1549),
.B2(n_1561),
.C(n_1577),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1497),
.A2(n_1555),
.B1(n_1569),
.B2(n_1445),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1553),
.B(n_1445),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1553),
.B(n_1569),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1557),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1522),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1587),
.A2(n_1555),
.B1(n_1588),
.B2(n_1580),
.C(n_1589),
.Y(n_1667)
);

AND2x4_ASAP7_75t_SL g1668 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1549),
.A2(n_1582),
.B1(n_1586),
.B2(n_1588),
.Y(n_1669)
);

AOI222xp33_ASAP7_75t_L g1670 ( 
.A1(n_1529),
.A2(n_1534),
.B1(n_1581),
.B2(n_1576),
.C1(n_1530),
.C2(n_1566),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1504),
.A2(n_1521),
.B1(n_1568),
.B2(n_1529),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1568),
.A2(n_1578),
.B1(n_959),
.B2(n_1429),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1578),
.B(n_1572),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_L g1674 ( 
.A(n_1429),
.B(n_959),
.C(n_726),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1507),
.A2(n_937),
.B(n_944),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1430),
.Y(n_1676)
);

AO21x2_ASAP7_75t_L g1677 ( 
.A1(n_1487),
.A2(n_1587),
.B(n_1485),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1440),
.A2(n_959),
.B1(n_726),
.B2(n_937),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1429),
.A2(n_726),
.B1(n_959),
.B2(n_818),
.C(n_938),
.Y(n_1680)
);

BUFx12f_ASAP7_75t_L g1681 ( 
.A(n_1441),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1507),
.A2(n_937),
.B(n_944),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1573),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1532),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_726),
.B2(n_818),
.C(n_1402),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1487),
.A2(n_1587),
.B(n_1485),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1430),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1490),
.B(n_1505),
.Y(n_1688)
);

OAI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1429),
.A2(n_818),
.B(n_1402),
.C(n_726),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_R g1693 ( 
.A(n_1441),
.B(n_912),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1429),
.B(n_959),
.C(n_726),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1437),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1490),
.B(n_1505),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1429),
.A2(n_938),
.B(n_959),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1429),
.A2(n_959),
.B(n_937),
.C(n_944),
.Y(n_1699)
);

BUFx4f_ASAP7_75t_SL g1700 ( 
.A(n_1532),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_1402),
.B2(n_771),
.C1(n_252),
.C2(n_305),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1430),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1537),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1487),
.A2(n_1516),
.B(n_1514),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1556),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1430),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1573),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1440),
.A2(n_959),
.B1(n_726),
.B2(n_937),
.Y(n_1708)
);

AOI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1429),
.A2(n_959),
.B(n_1272),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1495),
.A2(n_938),
.B1(n_959),
.B2(n_944),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1573),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_726),
.B2(n_818),
.C(n_1402),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1489),
.B(n_1486),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1463),
.B(n_1539),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1463),
.B(n_1539),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1532),
.A2(n_726),
.B1(n_818),
.B2(n_1144),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1437),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1430),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1572),
.B(n_1574),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1429),
.A2(n_959),
.B1(n_938),
.B2(n_937),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1572),
.B(n_1574),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1668),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1633),
.Y(n_1725)
);

OAI211xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1685),
.A2(n_1712),
.B(n_1701),
.C(n_1680),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1699),
.A2(n_1682),
.B(n_1675),
.Y(n_1727)
);

AOI222xp33_ASAP7_75t_L g1728 ( 
.A1(n_1717),
.A2(n_1689),
.B1(n_1698),
.B2(n_1695),
.C1(n_1690),
.C2(n_1692),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1595),
.B(n_1612),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1604),
.B(n_1620),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1595),
.B(n_1612),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1596),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1592),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1620),
.B(n_1715),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1603),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1736)
);

NAND2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1625),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1597),
.B(n_1663),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1597),
.B(n_1663),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1664),
.B(n_1704),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1676),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1664),
.B(n_1704),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1720),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1625),
.B(n_1673),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1625),
.B(n_1673),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1679),
.B(n_1708),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1687),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1626),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1677),
.B(n_1686),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1623),
.B(n_1667),
.Y(n_1751)
);

INVx5_ASAP7_75t_L g1752 ( 
.A(n_1624),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1677),
.B(n_1686),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1678),
.A2(n_1713),
.B1(n_1694),
.B2(n_1691),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1677),
.B(n_1686),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1670),
.B(n_1720),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1723),
.B(n_1651),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1702),
.Y(n_1758)
);

AND2x4_ASAP7_75t_SL g1759 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1759)
);

AO21x2_ASAP7_75t_L g1760 ( 
.A1(n_1657),
.A2(n_1645),
.B(n_1635),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1644),
.B(n_1671),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1706),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1626),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1648),
.B(n_1669),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1618),
.B(n_1661),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1668),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1611),
.B(n_1602),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1624),
.Y(n_1768)
);

OAI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1710),
.A2(n_1709),
.B1(n_1598),
.B2(n_1614),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1714),
.B(n_1703),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1721),
.A2(n_1722),
.B(n_1617),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1672),
.B(n_1605),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1653),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1630),
.B(n_1643),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1719),
.B(n_1629),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1631),
.B(n_1658),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1662),
.B(n_1658),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1688),
.B(n_1697),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1601),
.B(n_1600),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1624),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1647),
.Y(n_1781)
);

NAND4xp25_ASAP7_75t_L g1782 ( 
.A(n_1728),
.B(n_1674),
.C(n_1696),
.D(n_1718),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1778),
.B(n_1606),
.Y(n_1783)
);

OAI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1737),
.A2(n_1650),
.B(n_1599),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1732),
.B(n_1622),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1724),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1742),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1778),
.B(n_1711),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1778),
.B(n_1775),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1742),
.Y(n_1790)
);

NAND2xp33_ASAP7_75t_R g1791 ( 
.A(n_1765),
.B(n_1666),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1754),
.A2(n_1666),
.B1(n_1700),
.B2(n_1627),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1773),
.Y(n_1793)
);

OAI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1726),
.A2(n_1615),
.A3(n_1649),
.B(n_1638),
.Y(n_1794)
);

AOI33xp33_ASAP7_75t_L g1795 ( 
.A1(n_1765),
.A2(n_1621),
.A3(n_1634),
.B1(n_1646),
.B2(n_1619),
.B3(n_1636),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1738),
.B(n_1607),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1725),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1732),
.B(n_1738),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1732),
.B(n_1622),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1769),
.A2(n_1632),
.B1(n_1707),
.B2(n_1683),
.C(n_1642),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1775),
.B(n_1608),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1733),
.Y(n_1803)
);

INVxp67_ASAP7_75t_SL g1804 ( 
.A(n_1758),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_R g1805 ( 
.A(n_1765),
.B(n_1681),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1773),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1751),
.B(n_1660),
.C(n_1656),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1773),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1744),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1744),
.Y(n_1810)
);

AOI33xp33_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1640),
.A3(n_1641),
.B1(n_1613),
.B2(n_1652),
.B3(n_1637),
.Y(n_1811)
);

INVx4_ASAP7_75t_L g1812 ( 
.A(n_1752),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1733),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1738),
.B(n_1593),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1739),
.B(n_1594),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1748),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1733),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1776),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1726),
.A2(n_1639),
.B(n_1659),
.Y(n_1820)
);

OAI33xp33_ASAP7_75t_L g1821 ( 
.A1(n_1754),
.A2(n_1665),
.A3(n_1693),
.B1(n_1655),
.B2(n_1684),
.B3(n_1593),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1764),
.A2(n_1684),
.B1(n_1705),
.B2(n_1659),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_R g1823 ( 
.A(n_1774),
.B(n_1665),
.Y(n_1823)
);

OAI31xp33_ASAP7_75t_L g1824 ( 
.A1(n_1771),
.A2(n_1638),
.A3(n_1655),
.B(n_1628),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1770),
.Y(n_1825)
);

CKINVDCx16_ASAP7_75t_R g1826 ( 
.A(n_1767),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1747),
.A2(n_1659),
.B1(n_1705),
.B2(n_1681),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1776),
.B(n_1654),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1739),
.B(n_1654),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1781),
.B(n_1659),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1733),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1739),
.B(n_1659),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1762),
.Y(n_1833)
);

BUFx10_ASAP7_75t_L g1834 ( 
.A(n_1759),
.Y(n_1834)
);

AOI222xp33_ASAP7_75t_L g1835 ( 
.A1(n_1747),
.A2(n_1616),
.B1(n_1705),
.B2(n_1751),
.C1(n_1761),
.C2(n_1772),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1730),
.B(n_1705),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1762),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1752),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1728),
.B(n_1616),
.C(n_1705),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1771),
.A2(n_1616),
.B1(n_1761),
.B2(n_1772),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1729),
.B(n_1731),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1730),
.B(n_1745),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_1724),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1793),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1793),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1806),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1806),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1812),
.B(n_1735),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1841),
.B(n_1740),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1798),
.B(n_1842),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1841),
.B(n_1740),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1789),
.B(n_1818),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1803),
.Y(n_1853)
);

AND2x4_ASAP7_75t_SL g1854 ( 
.A(n_1834),
.B(n_1766),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1825),
.B(n_1740),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1782),
.A2(n_1761),
.B1(n_1774),
.B2(n_1772),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1798),
.B(n_1745),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1842),
.B(n_1756),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1804),
.B(n_1809),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1785),
.B(n_1745),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1808),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_SL g1862 ( 
.A(n_1801),
.B(n_1774),
.C(n_1764),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1743),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1808),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1819),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1803),
.Y(n_1866)
);

NOR2x1p5_ASAP7_75t_L g1867 ( 
.A(n_1839),
.B(n_1764),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1815),
.B(n_1743),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1815),
.B(n_1743),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1832),
.B(n_1746),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1785),
.B(n_1746),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1813),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1832),
.B(n_1746),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1799),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1826),
.B(n_1729),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1813),
.B(n_1729),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1810),
.B(n_1737),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1817),
.B(n_1731),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1812),
.B(n_1735),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1819),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1817),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1799),
.B(n_1731),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1831),
.B(n_1737),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1831),
.B(n_1737),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1829),
.B(n_1737),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_L g1886 ( 
.A(n_1812),
.B(n_1727),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1833),
.B(n_1756),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1833),
.B(n_1756),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1829),
.B(n_1755),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1837),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1838),
.B(n_1755),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1837),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1787),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1790),
.B(n_1757),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1800),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1816),
.B(n_1757),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1890),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1892),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1887),
.B(n_1888),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1887),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1854),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1852),
.B(n_1788),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1890),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1868),
.B(n_1786),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1856),
.B(n_1805),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1888),
.B(n_1814),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1892),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1854),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1854),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1886),
.A2(n_1862),
.B(n_1824),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1868),
.B(n_1786),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1893),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1893),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1893),
.Y(n_1914)
);

INVx2_ASAP7_75t_SL g1915 ( 
.A(n_1890),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1858),
.B(n_1814),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1858),
.B(n_1736),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1895),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1895),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1853),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1860),
.B(n_1736),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1895),
.Y(n_1922)
);

OAI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1856),
.A2(n_1840),
.B(n_1784),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1860),
.B(n_1828),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1894),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1852),
.B(n_1836),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1871),
.B(n_1797),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1876),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1886),
.B(n_1823),
.Y(n_1929)
);

AOI21xp33_ASAP7_75t_L g1930 ( 
.A1(n_1859),
.A2(n_1791),
.B(n_1835),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1859),
.B(n_1783),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1868),
.B(n_1843),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1894),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1848),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1871),
.B(n_1797),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1896),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1853),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1857),
.B(n_1734),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1896),
.B(n_1830),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1923),
.A2(n_1867),
.B1(n_1862),
.B2(n_1760),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1899),
.B(n_1916),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1898),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1907),
.Y(n_1943)
);

NOR2x1_ASAP7_75t_L g1944 ( 
.A(n_1929),
.B(n_1867),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1912),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1901),
.B(n_1869),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1905),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_L g1948 ( 
.A(n_1929),
.B(n_1822),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1901),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1869),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1899),
.B(n_1869),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1913),
.Y(n_1952)
);

AOI21xp33_ASAP7_75t_L g1953 ( 
.A1(n_1910),
.A2(n_1760),
.B(n_1802),
.Y(n_1953)
);

INVx4_ASAP7_75t_L g1954 ( 
.A(n_1908),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1909),
.B(n_1875),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1931),
.B(n_1870),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1916),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1914),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1918),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1919),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1922),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1909),
.B(n_1875),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1915),
.Y(n_1963)
);

INVxp67_ASAP7_75t_SL g1964 ( 
.A(n_1904),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_SL g1965 ( 
.A(n_1934),
.B(n_1820),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1904),
.B(n_1875),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1930),
.B(n_1870),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1906),
.B(n_1874),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1902),
.B(n_1870),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1926),
.A2(n_1821),
.B(n_1794),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1900),
.B(n_1873),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1917),
.B(n_1933),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1897),
.Y(n_1973)
);

OAI31xp33_ASAP7_75t_L g1974 ( 
.A1(n_1917),
.A2(n_1792),
.A3(n_1807),
.B(n_1891),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1906),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1911),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1915),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1925),
.B(n_1873),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1897),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1911),
.B(n_1849),
.Y(n_1980)
);

OAI33xp33_ASAP7_75t_L g1981 ( 
.A1(n_1936),
.A2(n_1847),
.A3(n_1861),
.B1(n_1865),
.B2(n_1864),
.B3(n_1880),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1903),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1921),
.B(n_1874),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1939),
.B(n_1873),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1942),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1942),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1943),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1972),
.B(n_1921),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_L g1989 ( 
.A(n_1953),
.B(n_1811),
.C(n_1795),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1945),
.Y(n_1990)
);

A2O1A1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1944),
.A2(n_1784),
.B(n_1827),
.C(n_1750),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1945),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1970),
.B(n_1932),
.Y(n_1993)
);

XNOR2x2_ASAP7_75t_L g1994 ( 
.A(n_1948),
.B(n_1932),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1967),
.B(n_1924),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1949),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1940),
.B(n_1889),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1974),
.A2(n_1947),
.B(n_1981),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1947),
.A2(n_1965),
.B1(n_1760),
.B2(n_1750),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1952),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1955),
.B(n_1889),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1955),
.B(n_1889),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1965),
.A2(n_1760),
.B1(n_1755),
.B2(n_1753),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1957),
.B(n_1924),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1952),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1964),
.B(n_1849),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1958),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1954),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1949),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1976),
.A2(n_1760),
.B1(n_1753),
.B2(n_1750),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1956),
.B(n_1938),
.Y(n_2011)
);

OAI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1975),
.A2(n_1934),
.B1(n_1877),
.B2(n_1891),
.C(n_1928),
.Y(n_2012)
);

NAND3xp33_ASAP7_75t_L g2013 ( 
.A(n_1954),
.B(n_1753),
.C(n_1779),
.Y(n_2013)
);

OA21x2_ASAP7_75t_L g2014 ( 
.A1(n_1973),
.A2(n_1920),
.B(n_1937),
.Y(n_2014)
);

O2A1O1Ixp33_ASAP7_75t_SL g2015 ( 
.A1(n_1963),
.A2(n_1928),
.B(n_1935),
.C(n_1927),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1958),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1954),
.A2(n_1938),
.B1(n_1857),
.B2(n_1882),
.Y(n_2017)
);

AOI21xp33_ASAP7_75t_L g2018 ( 
.A1(n_1960),
.A2(n_1961),
.B(n_1968),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1959),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1959),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1966),
.B(n_1934),
.Y(n_2021)
);

OAI321xp33_ASAP7_75t_L g2022 ( 
.A1(n_1998),
.A2(n_1962),
.A3(n_1941),
.B1(n_1968),
.B2(n_1971),
.C(n_1950),
.Y(n_2022)
);

OAI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_2003),
.A2(n_1983),
.B1(n_1941),
.B2(n_1951),
.Y(n_2023)
);

OAI221xp5_ASAP7_75t_SL g2024 ( 
.A1(n_1999),
.A2(n_1962),
.B1(n_1983),
.B2(n_1951),
.C(n_1946),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1989),
.B(n_1966),
.Y(n_2025)
);

BUFx3_ASAP7_75t_L g2026 ( 
.A(n_2008),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2019),
.Y(n_2027)
);

OAI32xp33_ASAP7_75t_L g2028 ( 
.A1(n_1994),
.A2(n_1977),
.A3(n_1946),
.B1(n_1950),
.B2(n_1935),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2009),
.B(n_1996),
.Y(n_2029)
);

NAND2x1_ASAP7_75t_L g2030 ( 
.A(n_2008),
.B(n_1980),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1999),
.A2(n_1969),
.B1(n_1980),
.B2(n_1984),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2019),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_SL g2033 ( 
.A1(n_1991),
.A2(n_1838),
.B(n_1982),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1985),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1986),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1989),
.A2(n_1891),
.B1(n_1779),
.B2(n_1879),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1990),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1992),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1993),
.B(n_1978),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1996),
.B(n_1849),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2018),
.A2(n_1979),
.B1(n_1973),
.B2(n_1982),
.C(n_1779),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2013),
.A2(n_1848),
.B1(n_1879),
.B2(n_1838),
.Y(n_2042)
);

NAND4xp25_ASAP7_75t_SL g2043 ( 
.A(n_1991),
.B(n_1927),
.C(n_1855),
.D(n_1863),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2000),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1987),
.B(n_1851),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2021),
.B(n_1851),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2005),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_2004),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2029),
.B(n_1995),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_2022),
.A2(n_2015),
.B(n_1997),
.Y(n_2050)
);

XNOR2x2_ASAP7_75t_L g2051 ( 
.A(n_2025),
.B(n_2010),
.Y(n_2051)
);

OAI21xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2039),
.A2(n_2012),
.B(n_2021),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2048),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2027),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2032),
.Y(n_2055)
);

NAND4xp75_ASAP7_75t_L g2056 ( 
.A(n_2029),
.B(n_2020),
.C(n_2016),
.D(n_2007),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2039),
.B(n_2001),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2026),
.B(n_2002),
.Y(n_2058)
);

INVxp67_ASAP7_75t_SL g2059 ( 
.A(n_2026),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2034),
.Y(n_2060)
);

INVxp67_ASAP7_75t_L g2061 ( 
.A(n_2035),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2037),
.B(n_1988),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2030),
.Y(n_2063)
);

NOR2x1_ASAP7_75t_L g2064 ( 
.A(n_2030),
.B(n_2014),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2038),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2044),
.B(n_2015),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_2047),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_2046),
.B(n_2006),
.Y(n_2068)
);

NAND3xp33_ASAP7_75t_L g2069 ( 
.A(n_2050),
.B(n_2041),
.C(n_2024),
.Y(n_2069)
);

AND3x2_ASAP7_75t_L g2070 ( 
.A(n_2059),
.B(n_2033),
.C(n_2028),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2059),
.B(n_2053),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2067),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_L g2073 ( 
.A(n_2056),
.B(n_2033),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2052),
.A2(n_2043),
.B1(n_2068),
.B2(n_2058),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_SL g2075 ( 
.A(n_2051),
.B(n_2036),
.C(n_2031),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_2063),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2049),
.B(n_2046),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2057),
.B(n_2023),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2067),
.B(n_2040),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2068),
.B(n_2045),
.Y(n_2080)
);

NOR3x1_ASAP7_75t_L g2081 ( 
.A(n_2075),
.B(n_2055),
.C(n_2054),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_L g2082 ( 
.A(n_2070),
.B(n_2066),
.C(n_2061),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2069),
.A2(n_2062),
.B1(n_2064),
.B2(n_2063),
.C(n_2061),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2071),
.B(n_2072),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_SL g2085 ( 
.A(n_2073),
.B(n_2060),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2074),
.A2(n_2042),
.B1(n_2068),
.B2(n_2017),
.Y(n_2086)
);

A2O1A1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_2078),
.A2(n_2065),
.B(n_2011),
.C(n_1848),
.Y(n_2087)
);

AOI211x1_ASAP7_75t_L g2088 ( 
.A1(n_2077),
.A2(n_1855),
.B(n_1863),
.C(n_1885),
.Y(n_2088)
);

AOI211xp5_ASAP7_75t_L g2089 ( 
.A1(n_2079),
.A2(n_1879),
.B(n_1848),
.C(n_1877),
.Y(n_2089)
);

O2A1O1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_2076),
.A2(n_2014),
.B(n_1763),
.C(n_1749),
.Y(n_2090)
);

AOI221xp5_ASAP7_75t_SL g2091 ( 
.A1(n_2076),
.A2(n_1903),
.B1(n_1937),
.B2(n_1920),
.C(n_1863),
.Y(n_2091)
);

NOR2x1_ASAP7_75t_L g2092 ( 
.A(n_2082),
.B(n_2080),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2084),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2083),
.A2(n_2014),
.B(n_1741),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2085),
.Y(n_2095)
);

NAND4xp25_ASAP7_75t_SL g2096 ( 
.A(n_2087),
.B(n_1877),
.C(n_1855),
.D(n_1885),
.Y(n_2096)
);

AOI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_2086),
.A2(n_1763),
.B1(n_1749),
.B2(n_1885),
.C(n_1848),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2081),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2088),
.B(n_2089),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2095),
.B(n_2091),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_R g2101 ( 
.A(n_2093),
.B(n_2090),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2092),
.B(n_1851),
.Y(n_2102)
);

AND2x2_ASAP7_75t_SL g2103 ( 
.A(n_2098),
.B(n_2099),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2097),
.B(n_1876),
.Y(n_2104)
);

NAND4xp75_ASAP7_75t_L g2105 ( 
.A(n_2094),
.B(n_1796),
.C(n_1884),
.D(n_1883),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2096),
.B(n_1879),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2103),
.B(n_1883),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2102),
.Y(n_2108)
);

NOR2x1_ASAP7_75t_L g2109 ( 
.A(n_2100),
.B(n_1843),
.Y(n_2109)
);

NOR4xp25_ASAP7_75t_L g2110 ( 
.A(n_2101),
.B(n_1847),
.C(n_1844),
.D(n_1861),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2104),
.A2(n_1850),
.B1(n_1879),
.B2(n_1882),
.Y(n_2111)
);

NAND5xp2_ASAP7_75t_L g2112 ( 
.A(n_2105),
.B(n_1796),
.C(n_1780),
.D(n_1768),
.E(n_1777),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2112),
.B(n_2106),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2109),
.B(n_2106),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2108),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_2110),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2114),
.B(n_2107),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2117),
.A2(n_2113),
.B1(n_2115),
.B2(n_2116),
.Y(n_2118)
);

AOI221xp5_ASAP7_75t_R g2119 ( 
.A1(n_2118),
.A2(n_2116),
.B1(n_2111),
.B2(n_1766),
.C(n_1866),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_2118),
.Y(n_2120)
);

XOR2xp5_ASAP7_75t_L g2121 ( 
.A(n_2120),
.B(n_2119),
.Y(n_2121)
);

OAI22x1_ASAP7_75t_L g2122 ( 
.A1(n_2120),
.A2(n_1752),
.B1(n_1866),
.B2(n_1853),
.Y(n_2122)
);

AOI222xp33_ASAP7_75t_L g2123 ( 
.A1(n_2122),
.A2(n_1864),
.B1(n_1846),
.B2(n_1844),
.C1(n_1845),
.C2(n_1865),
.Y(n_2123)
);

AOI221xp5_ASAP7_75t_L g2124 ( 
.A1(n_2121),
.A2(n_1846),
.B1(n_1880),
.B2(n_1845),
.C(n_1881),
.Y(n_2124)
);

AOI322xp5_ASAP7_75t_L g2125 ( 
.A1(n_2124),
.A2(n_1780),
.A3(n_1768),
.B1(n_1884),
.B2(n_1883),
.C1(n_1878),
.C2(n_1876),
.Y(n_2125)
);

AOI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2125),
.A2(n_2123),
.B1(n_1881),
.B2(n_1758),
.C(n_1872),
.Y(n_2126)
);

AOI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2126),
.A2(n_1850),
.B(n_1884),
.C(n_1872),
.Y(n_2127)
);


endmodule