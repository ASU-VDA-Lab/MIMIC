module fake_jpeg_7993_n_257 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_46),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_23),
.B1(n_34),
.B2(n_20),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_66),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_27),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_45),
.B1(n_36),
.B2(n_46),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_92),
.B1(n_28),
.B2(n_31),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_78),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_59),
.B1(n_51),
.B2(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_82),
.B1(n_21),
.B2(n_31),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_85),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_51),
.B1(n_50),
.B2(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_65),
.B1(n_57),
.B2(n_62),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_36),
.B1(n_21),
.B2(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_36),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_25),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_37),
.C(n_40),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_105),
.B1(n_107),
.B2(n_71),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_40),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_65),
.B1(n_29),
.B2(n_26),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_53),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_25),
.B(n_35),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_22),
.B(n_24),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_91),
.B1(n_85),
.B2(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_128),
.Y(n_158)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_141),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_98),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_139),
.B(n_22),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_131),
.B1(n_135),
.B2(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_71),
.B1(n_79),
.B2(n_86),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_140),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_79),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_83),
.B1(n_70),
.B2(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_83),
.B1(n_70),
.B2(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_26),
.B1(n_18),
.B2(n_37),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_113),
.B1(n_112),
.B2(n_18),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_64),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_0),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_110),
.B(n_103),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_144),
.B(n_104),
.Y(n_154)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_139),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_97),
.C(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_124),
.C(n_138),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_134),
.B1(n_136),
.B2(n_25),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_113),
.B1(n_118),
.B2(n_112),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_35),
.B1(n_25),
.B2(n_32),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_64),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_35),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_60),
.A3(n_32),
.B1(n_35),
.B2(n_25),
.C1(n_24),
.C2(n_22),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_183),
.C(n_186),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_188),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_132),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_147),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_32),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_156),
.B1(n_168),
.B2(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_35),
.B1(n_32),
.B2(n_25),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_165),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_199),
.B1(n_202),
.B2(n_207),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_152),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_208),
.B(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_157),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_201),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_153),
.C(n_155),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_206),
.B(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_159),
.C(n_145),
.Y(n_205)
);

OAI321xp33_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_154),
.A3(n_145),
.B1(n_157),
.B2(n_161),
.C(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_158),
.B(n_183),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_190),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_221),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_5),
.B(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_184),
.B1(n_189),
.B2(n_171),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_222),
.B(n_213),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_188),
.B1(n_146),
.B2(n_186),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_220),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_151),
.B(n_35),
.C(n_4),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_198),
.B(n_200),
.C(n_7),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_231),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_230),
.B(n_8),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_197),
.C(n_205),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.C(n_232),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_197),
.C(n_194),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_22),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_22),
.C(n_7),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_215),
.Y(n_235)
);

OAI321xp33_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_236),
.A3(n_240),
.B1(n_219),
.B2(n_9),
.C(n_10),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_211),
.B1(n_209),
.B2(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_224),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_6),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_226),
.C(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_245),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_219),
.B(n_22),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_246),
.B(n_236),
.Y(n_247)
);

AOI31xp33_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_11),
.A3(n_12),
.B(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_8),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_8),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_237),
.B(n_233),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_13),
.C(n_14),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_12),
.B(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_253),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_252),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_15),
.Y(n_257)
);


endmodule