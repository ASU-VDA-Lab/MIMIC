module fake_netlist_6_1360_n_1104 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_113, n_39, n_63, n_223, n_270, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1104);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_270;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1104;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_886;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_901;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_683;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_569;
wire n_1092;
wire n_441;
wire n_1060;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_127),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_211),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_83),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_186),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_46),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_222),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_193),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_14),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_112),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_66),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_130),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_250),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_50),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_203),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_216),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_137),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_106),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_90),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_260),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_199),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_172),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_4),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_105),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_114),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_34),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_230),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_86),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_158),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_142),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_163),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_141),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_138),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_177),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_40),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_30),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_241),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_212),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_4),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_15),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_68),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_116),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_104),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_98),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_225),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_16),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_52),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_280),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_280),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_0),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_334),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_0),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_1),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_282),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_283),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_1),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_284),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_286),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_287),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_289),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_291),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_292),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_308),
.B(n_2),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_296),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_318),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_318),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_293),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_2),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_326),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_354),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_357),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_362),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_344),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_372),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_306),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_374),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_347),
.B(n_288),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_344),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_326),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_367),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_316),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_375),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_345),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_379),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_345),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_340),
.B(n_306),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_364),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_380),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_299),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_294),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_430),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_428),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_300),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_327),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

BUFx4f_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_301),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_412),
.B(n_340),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_319),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_429),
.A2(n_340),
.B1(n_342),
.B2(n_333),
.Y(n_454)
);

BUFx8_ASAP7_75t_SL g455 ( 
.A(n_402),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_303),
.Y(n_456)
);

BUFx8_ASAP7_75t_SL g457 ( 
.A(n_402),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_409),
.B(n_304),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_409),
.B(n_319),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_340),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_410),
.A2(n_307),
.B1(n_310),
.B2(n_305),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_313),
.B1(n_314),
.B2(n_311),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_392),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_433),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_320),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_428),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_416),
.B(n_324),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_391),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_416),
.B(n_328),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_390),
.B(n_329),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_331),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_395),
.B(n_337),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_415),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_341),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_414),
.B(n_383),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_420),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_410),
.B(n_343),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_394),
.B(n_384),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_3),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_450),
.B(n_424),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_470),
.B(n_431),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_450),
.B(n_424),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_405),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_439),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_441),
.B(n_399),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_470),
.B(n_431),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_444),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_456),
.B(n_411),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_417),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_444),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_471),
.B(n_418),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_445),
.A2(n_419),
.B(n_384),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_446),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_471),
.B(n_400),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_502),
.B(n_400),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_502),
.B(n_400),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_477),
.B(n_39),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_459),
.A2(n_425),
.B1(n_439),
.B2(n_435),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_500),
.B(n_41),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_448),
.B(n_477),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_449),
.B(n_43),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_479),
.B(n_439),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_44),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_47),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_448),
.B(n_432),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_454),
.A2(n_432),
.B1(n_435),
.B2(n_413),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_466),
.B(n_437),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_48),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_478),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_466),
.B(n_454),
.Y(n_543)
);

AOI221xp5_ASAP7_75t_L g544 ( 
.A1(n_501),
.A2(n_483),
.B1(n_463),
.B2(n_451),
.C(n_467),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_453),
.A2(n_437),
.B1(n_6),
.B2(n_3),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_462),
.Y(n_546)
);

AND2x6_ASAP7_75t_SL g547 ( 
.A(n_497),
.B(n_5),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_486),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_481),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_49),
.Y(n_550)
);

BUFx5_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_486),
.B(n_5),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_486),
.B(n_6),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_499),
.B(n_51),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_7),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_493),
.B(n_53),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_476),
.B(n_54),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_55),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_504),
.B(n_7),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_464),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_440),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_458),
.B(n_8),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_501),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_564)
);

AND2x6_ASAP7_75t_SL g565 ( 
.A(n_464),
.B(n_9),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_482),
.B(n_56),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_484),
.B(n_57),
.Y(n_567)
);

NAND2x1_ASAP7_75t_L g568 ( 
.A(n_469),
.B(n_58),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_488),
.B(n_59),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_495),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_473),
.B(n_13),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_SL g574 ( 
.A(n_544),
.B(n_472),
.C(n_503),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_551),
.B(n_473),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_507),
.A2(n_490),
.B(n_483),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_512),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_512),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_510),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_517),
.B(n_465),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_543),
.A2(n_562),
.B1(n_515),
.B2(n_507),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_520),
.B(n_465),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_513),
.A2(n_548),
.B1(n_524),
.B2(n_532),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_475),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_513),
.A2(n_529),
.B1(n_508),
.B2(n_506),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_523),
.A2(n_464),
.B1(n_475),
.B2(n_492),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_551),
.B(n_492),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_496),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_559),
.A2(n_489),
.B(n_469),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_540),
.B(n_461),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_522),
.A2(n_494),
.B(n_460),
.C(n_480),
.Y(n_593)
);

AOI21xp33_ASAP7_75t_L g594 ( 
.A1(n_573),
.A2(n_494),
.B(n_480),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_533),
.A2(n_489),
.B(n_469),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_559),
.A2(n_494),
.B(n_460),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_551),
.A2(n_461),
.B1(n_485),
.B2(n_480),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_559),
.A2(n_494),
.B(n_460),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_534),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_551),
.B(n_461),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_510),
.B(n_485),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_558),
.A2(n_61),
.B(n_60),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_559),
.A2(n_63),
.B(n_62),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_546),
.B(n_485),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_514),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_67),
.B(n_64),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_539),
.B(n_455),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_570),
.A2(n_70),
.B(n_69),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_564),
.B(n_487),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_510),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_556),
.A2(n_72),
.B(n_71),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_514),
.B(n_487),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_538),
.B(n_487),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_13),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_558),
.A2(n_74),
.B(n_73),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_567),
.A2(n_76),
.B(n_75),
.Y(n_617)
);

AND3x4_ASAP7_75t_L g618 ( 
.A(n_534),
.B(n_457),
.C(n_455),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_567),
.A2(n_78),
.B(n_77),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_80),
.B(n_79),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_560),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_557),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_552),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_527),
.B(n_17),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_527),
.B(n_18),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_571),
.A2(n_82),
.B(n_81),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_519),
.B(n_18),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_530),
.B(n_526),
.C(n_525),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_535),
.A2(n_87),
.B(n_85),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_536),
.A2(n_89),
.B(n_88),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_531),
.A2(n_92),
.B(n_91),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_550),
.A2(n_94),
.B(n_93),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_553),
.A2(n_173),
.B1(n_277),
.B2(n_276),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_578),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_528),
.B(n_521),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_585),
.B(n_509),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_595),
.A2(n_566),
.B(n_541),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_561),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_589),
.A2(n_531),
.B(n_541),
.Y(n_641)
);

O2A1O1Ixp5_ASAP7_75t_L g642 ( 
.A1(n_584),
.A2(n_554),
.B(n_568),
.C(n_563),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_605),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_608),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_627),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_575),
.A2(n_518),
.B(n_549),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_581),
.B(n_545),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_600),
.B(n_537),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_579),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_591),
.A2(n_572),
.B(n_96),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_613),
.B(n_565),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_586),
.A2(n_97),
.B(n_95),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_577),
.B(n_19),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_583),
.A2(n_100),
.B(n_99),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_608),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_608),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_614),
.B(n_19),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_20),
.Y(n_658)
);

AOI21xp33_ASAP7_75t_L g659 ( 
.A1(n_592),
.A2(n_20),
.B(n_21),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g660 ( 
.A1(n_587),
.A2(n_178),
.B(n_274),
.C(n_273),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_634),
.Y(n_661)
);

AO31x2_ASAP7_75t_L g662 ( 
.A1(n_593),
.A2(n_21),
.A3(n_22),
.B(n_23),
.Y(n_662)
);

CKINVDCx8_ASAP7_75t_R g663 ( 
.A(n_622),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_576),
.A2(n_102),
.B(n_101),
.Y(n_664)
);

OAI21x1_ASAP7_75t_SL g665 ( 
.A1(n_617),
.A2(n_107),
.B(n_103),
.Y(n_665)
);

BUFx4_ASAP7_75t_R g666 ( 
.A(n_618),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_576),
.A2(n_109),
.B(n_108),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_596),
.A2(n_111),
.B(n_110),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_597),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_457),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_SL g673 ( 
.A(n_629),
.B(n_547),
.C(n_22),
.Y(n_673)
);

OAI21x1_ASAP7_75t_SL g674 ( 
.A1(n_617),
.A2(n_115),
.B(n_113),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_615),
.A2(n_623),
.A3(n_624),
.B(n_625),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_598),
.A2(n_118),
.B(n_117),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_588),
.A2(n_120),
.B(n_119),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_611),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_612),
.A2(n_122),
.B(n_121),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_632),
.A2(n_124),
.B(n_123),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_601),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_632),
.A2(n_189),
.B(n_271),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_602),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_616),
.A2(n_620),
.B(n_619),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_626),
.A2(n_187),
.B(n_270),
.Y(n_685)
);

NOR2x1_ASAP7_75t_L g686 ( 
.A(n_604),
.B(n_125),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_610),
.B(n_23),
.Y(n_687)
);

NAND2x1_ASAP7_75t_L g688 ( 
.A(n_590),
.B(n_126),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_610),
.B(n_24),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_607),
.B(n_128),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_594),
.A2(n_191),
.B(n_269),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_635),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_630),
.A2(n_190),
.B(n_268),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_691),
.B(n_601),
.Y(n_695)
);

INVx3_ASAP7_75t_SL g696 ( 
.A(n_668),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_672),
.A2(n_633),
.B1(n_631),
.B2(n_609),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_663),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_691),
.B(n_603),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_644),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_SL g701 ( 
.A1(n_680),
.A2(n_693),
.B(n_682),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_638),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_644),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_690),
.A2(n_606),
.B1(n_25),
.B2(n_26),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_668),
.Y(n_705)
);

O2A1O1Ixp5_ASAP7_75t_L g706 ( 
.A1(n_639),
.A2(n_685),
.B(n_642),
.C(n_660),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_646),
.A2(n_185),
.B(n_267),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_671),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_651),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_647),
.B(n_667),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_678),
.B(n_27),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_668),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_653),
.B(n_27),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_636),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_644),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_658),
.B(n_28),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_SL g717 ( 
.A1(n_692),
.A2(n_194),
.B(n_266),
.C(n_265),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_645),
.B(n_28),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_648),
.B(n_29),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_681),
.B(n_640),
.Y(n_722)
);

AOI221xp5_ASAP7_75t_L g723 ( 
.A1(n_673),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_687),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_636),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_661),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_667),
.B(n_33),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_640),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_684),
.A2(n_196),
.B(n_264),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_689),
.B(n_657),
.Y(n_730)
);

AOI21x1_ASAP7_75t_L g731 ( 
.A1(n_641),
.A2(n_195),
.B(n_263),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_643),
.B(n_34),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_686),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_733)
);

AND2x2_ASAP7_75t_SL g734 ( 
.A(n_656),
.B(n_35),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_655),
.B(n_272),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_649),
.B(n_36),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_656),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_649),
.B(n_37),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_659),
.A2(n_38),
.B1(n_129),
.B2(n_131),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_666),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_688),
.B(n_132),
.Y(n_742)
);

CKINVDCx11_ASAP7_75t_R g743 ( 
.A(n_665),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_133),
.Y(n_744)
);

BUFx8_ASAP7_75t_L g745 ( 
.A(n_662),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_675),
.B(n_134),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_683),
.A2(n_201),
.B(n_135),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_675),
.B(n_637),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_677),
.B(n_38),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_714),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_725),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_710),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_726),
.Y(n_754)
);

INVx6_ASAP7_75t_L g755 ( 
.A(n_737),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_701),
.A2(n_669),
.B1(n_664),
.B2(n_654),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_734),
.A2(n_674),
.B1(n_650),
.B2(n_652),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_746),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_721),
.A2(n_662),
.B1(n_679),
.B2(n_676),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_737),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_698),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_702),
.A2(n_694),
.B1(n_675),
.B2(n_140),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_718),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_736),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_738),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_695),
.B(n_699),
.Y(n_766)
);

NOR2x1_ASAP7_75t_R g767 ( 
.A(n_728),
.B(n_262),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_708),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_706),
.A2(n_136),
.B(n_139),
.Y(n_769)
);

AOI21x1_ASAP7_75t_L g770 ( 
.A1(n_730),
.A2(n_143),
.B(n_144),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_723),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_771)
);

BUFx8_ASAP7_75t_L g772 ( 
.A(n_705),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_716),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_724),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_709),
.A2(n_261),
.B1(n_155),
.B2(n_156),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_696),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_741),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_704),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_SL g780 ( 
.A1(n_713),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_720),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_695),
.B(n_164),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_722),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_722),
.A2(n_169),
.B1(n_170),
.B2(n_174),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_733),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_712),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_732),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_719),
.B(n_181),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_739),
.A2(n_259),
.B1(n_183),
.B2(n_184),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_737),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_SL g791 ( 
.A1(n_735),
.A2(n_182),
.B1(n_192),
.B2(n_197),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_735),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_746),
.Y(n_794)
);

NOR2x1_ASAP7_75t_L g795 ( 
.A(n_711),
.B(n_198),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_743),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_700),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_748),
.A2(n_200),
.B(n_202),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_731),
.A2(n_204),
.B(n_205),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_745),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_700),
.B(n_209),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_703),
.B(n_210),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_749),
.A2(n_258),
.B1(n_214),
.B2(n_217),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_703),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_697),
.A2(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_703),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_715),
.Y(n_807)
);

OAI22x1_ASAP7_75t_L g808 ( 
.A1(n_699),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_715),
.Y(n_809)
);

OA21x2_ASAP7_75t_L g810 ( 
.A1(n_731),
.A2(n_226),
.B(n_227),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_756),
.A2(n_717),
.B(n_729),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_753),
.B(n_773),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_750),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_751),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_751),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_781),
.Y(n_816)
);

INVxp33_ASAP7_75t_SL g817 ( 
.A(n_761),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_750),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_782),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_769),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_769),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_762),
.A2(n_747),
.B(n_707),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_782),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_778),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

AO21x2_ASAP7_75t_L g827 ( 
.A1(n_798),
.A2(n_745),
.B(n_744),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_771),
.A2(n_742),
.B(n_715),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_758),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_764),
.B(n_229),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_752),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_798),
.A2(n_770),
.B(n_805),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_765),
.B(n_787),
.Y(n_834)
);

AND2x4_ASAP7_75t_SL g835 ( 
.A(n_794),
.B(n_231),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_799),
.A2(n_810),
.B(n_766),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_799),
.Y(n_837)
);

HB1xp67_ASAP7_75t_SL g838 ( 
.A(n_772),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_799),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_755),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_810),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_810),
.Y(n_842)
);

OA21x2_ASAP7_75t_L g843 ( 
.A1(n_771),
.A2(n_232),
.B(n_233),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_766),
.B(n_234),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_803),
.A2(n_235),
.B(n_236),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_803),
.A2(n_237),
.B(n_240),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_793),
.B(n_257),
.Y(n_847)
);

OA21x2_ASAP7_75t_L g848 ( 
.A1(n_789),
.A2(n_242),
.B(n_246),
.Y(n_848)
);

OAI21xp33_ASAP7_75t_SL g849 ( 
.A1(n_789),
.A2(n_247),
.B(n_248),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_759),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_755),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_800),
.B(n_249),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_768),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_778),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_759),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_757),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_800),
.B(n_802),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_757),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_808),
.A2(n_251),
.B(n_252),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_782),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_797),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_807),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_814),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_819),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_850),
.B(n_780),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_826),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_836),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_861),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_850),
.B(n_780),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_855),
.B(n_809),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_814),
.Y(n_871)
);

NAND4xp25_ASAP7_75t_SL g872 ( 
.A(n_852),
.B(n_776),
.C(n_775),
.D(n_795),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_815),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_815),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_826),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_830),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_855),
.B(n_791),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_852),
.A2(n_776),
.B1(n_775),
.B2(n_785),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_861),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_856),
.B(n_806),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_837),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_818),
.Y(n_883)
);

INVx5_ASAP7_75t_SL g884 ( 
.A(n_827),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_818),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_813),
.B(n_790),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_817),
.B(n_786),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_860),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_856),
.B(n_858),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_813),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_858),
.B(n_862),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_862),
.B(n_804),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_837),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_834),
.B(n_788),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_834),
.B(n_790),
.Y(n_895)
);

AND2x4_ASAP7_75t_SL g896 ( 
.A(n_819),
.B(n_763),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_860),
.B(n_760),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_839),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_860),
.B(n_760),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_839),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_819),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_820),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_832),
.B(n_801),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_820),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_841),
.B(n_792),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_820),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_812),
.B(n_792),
.Y(n_908)
);

CKINVDCx14_ASAP7_75t_R g909 ( 
.A(n_853),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_841),
.B(n_796),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_819),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_823),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_879),
.A2(n_857),
.B(n_828),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_897),
.B(n_823),
.Y(n_914)
);

NAND2x1_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_823),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_888),
.B(n_842),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_872),
.B(n_849),
.C(n_823),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_865),
.A2(n_843),
.B1(n_848),
.B2(n_849),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_842),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_865),
.A2(n_843),
.B1(n_848),
.B2(n_857),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_889),
.B(n_821),
.Y(n_921)
);

AND2x2_ASAP7_75t_SL g922 ( 
.A(n_896),
.B(n_848),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_SL g923 ( 
.A1(n_869),
.A2(n_878),
.B(n_896),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_864),
.B(n_851),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_863),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_898),
.B(n_831),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_898),
.B(n_831),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_900),
.B(n_844),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_910),
.B(n_774),
.C(n_848),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_SL g930 ( 
.A1(n_869),
.A2(n_843),
.B1(n_845),
.B2(n_846),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_910),
.B(n_900),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_889),
.B(n_844),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_904),
.B(n_840),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_903),
.A2(n_825),
.B(n_821),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_866),
.B(n_854),
.Y(n_935)
);

AND4x1_ASAP7_75t_L g936 ( 
.A(n_887),
.B(n_829),
.C(n_838),
.D(n_847),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_875),
.B(n_824),
.Y(n_937)
);

OAI221xp5_ASAP7_75t_L g938 ( 
.A1(n_878),
.A2(n_779),
.B1(n_843),
.B2(n_763),
.C(n_777),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_891),
.A2(n_859),
.B(n_847),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_904),
.B(n_784),
.C(n_783),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_891),
.B(n_840),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_864),
.B(n_859),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_931),
.B(n_876),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_921),
.B(n_877),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_926),
.B(n_880),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_935),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_934),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_937),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_921),
.B(n_884),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_916),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_925),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_934),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_916),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_922),
.B(n_884),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_922),
.B(n_884),
.Y(n_955)
);

AND2x4_ASAP7_75t_SL g956 ( 
.A(n_917),
.B(n_894),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_919),
.B(n_884),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_927),
.B(n_870),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_919),
.B(n_873),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_934),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_933),
.B(n_870),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_924),
.B(n_902),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_914),
.B(n_884),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_915),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_928),
.B(n_868),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_923),
.B(n_906),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_941),
.B(n_873),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_951),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_948),
.B(n_909),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_959),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_946),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_948),
.B(n_913),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_964),
.B(n_942),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_951),
.B(n_871),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_945),
.B(n_932),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_962),
.B(n_902),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_959),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_967),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_953),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_966),
.B(n_902),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_958),
.B(n_863),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_874),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_966),
.B(n_911),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_968),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_938),
.B(n_942),
.C(n_939),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_974),
.Y(n_986)
);

AOI21xp33_ASAP7_75t_L g987 ( 
.A1(n_972),
.A2(n_956),
.B(n_964),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_980),
.B(n_948),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_970),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_974),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_973),
.B(n_954),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_963),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_978),
.B(n_965),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_982),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_971),
.B(n_963),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_989),
.B(n_977),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_992),
.B(n_976),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_991),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_976),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_984),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_SL g1001 ( 
.A(n_991),
.B(n_920),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_984),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_985),
.B1(n_920),
.B2(n_956),
.Y(n_1004)
);

OA21x2_ASAP7_75t_L g1005 ( 
.A1(n_998),
.A2(n_987),
.B(n_989),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_1003),
.Y(n_1006)
);

AOI22x1_ASAP7_75t_L g1007 ( 
.A1(n_998),
.A2(n_994),
.B1(n_990),
.B2(n_986),
.Y(n_1007)
);

OAI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_996),
.A2(n_993),
.B1(n_969),
.B2(n_946),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_1006),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1007),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1005),
.B(n_997),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1008),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_1002),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_1009),
.A2(n_1012),
.B(n_1010),
.Y(n_1014)
);

AOI322xp5_ASAP7_75t_L g1015 ( 
.A1(n_1013),
.A2(n_1001),
.A3(n_1000),
.B1(n_999),
.B2(n_918),
.C1(n_995),
.C2(n_979),
.Y(n_1015)
);

AOI211xp5_ASAP7_75t_L g1016 ( 
.A1(n_1011),
.A2(n_985),
.B(n_929),
.C(n_777),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_1009),
.B(n_754),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_754),
.C(n_767),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_936),
.C(n_930),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1009),
.B(n_982),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1017),
.A2(n_955),
.B1(n_954),
.B2(n_881),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1020),
.Y(n_1022)
);

OAI211xp5_ASAP7_75t_SL g1023 ( 
.A1(n_1014),
.A2(n_918),
.B(n_975),
.C(n_961),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1019),
.B(n_960),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1018),
.B(n_979),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_1015),
.B(n_981),
.Y(n_1026)
);

OAI321xp33_ASAP7_75t_L g1027 ( 
.A1(n_1026),
.A2(n_1016),
.A3(n_955),
.B1(n_940),
.B2(n_908),
.C(n_851),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1024),
.A2(n_960),
.B(n_950),
.C(n_947),
.Y(n_1028)
);

OAI211xp5_ASAP7_75t_SL g1029 ( 
.A1(n_1022),
.A2(n_908),
.B(n_953),
.C(n_886),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_1025),
.B(n_881),
.C(n_892),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_892),
.C(n_867),
.Y(n_1031)
);

NAND4xp25_ASAP7_75t_SL g1032 ( 
.A(n_1023),
.B(n_957),
.C(n_949),
.D(n_965),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_1022),
.B(n_846),
.C(n_845),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_943),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_1028),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1034),
.Y(n_1036)
);

NOR2x2_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_952),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1030),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1032),
.A2(n_957),
.B1(n_949),
.B2(n_896),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1029),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1033),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_SL g1044 ( 
.A(n_1034),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1032),
.A2(n_755),
.B1(n_912),
.B2(n_895),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1034),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1034),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_1036),
.B(n_943),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1043),
.B(n_944),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_944),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_1035),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_864),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_1047),
.B(n_867),
.C(n_947),
.Y(n_1053)
);

AOI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_1041),
.A2(n_1040),
.B1(n_1038),
.B2(n_1042),
.C(n_1037),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1045),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1039),
.A2(n_952),
.B1(n_912),
.B2(n_911),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1044),
.B(n_864),
.Y(n_1057)
);

NAND2x1_ASAP7_75t_L g1058 ( 
.A(n_1038),
.B(n_894),
.Y(n_1058)
);

AOI32xp33_ASAP7_75t_L g1059 ( 
.A1(n_1035),
.A2(n_835),
.A3(n_911),
.B1(n_906),
.B2(n_895),
.Y(n_1059)
);

NOR4xp25_ASAP7_75t_L g1060 ( 
.A(n_1036),
.B(n_871),
.C(n_874),
.D(n_886),
.Y(n_1060)
);

AND3x4_ASAP7_75t_L g1061 ( 
.A(n_1044),
.B(n_864),
.C(n_905),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1038),
.B(n_864),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1036),
.B(n_867),
.C(n_883),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1044),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1036),
.B(n_867),
.C(n_883),
.Y(n_1065)
);

NOR3x2_ASAP7_75t_L g1066 ( 
.A(n_1044),
.B(n_835),
.C(n_255),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

XNOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1064),
.B(n_254),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_1058),
.Y(n_1069)
);

NAND4xp75_ASAP7_75t_L g1070 ( 
.A(n_1054),
.B(n_822),
.C(n_256),
.D(n_885),
.Y(n_1070)
);

NAND4xp25_ASAP7_75t_SL g1071 ( 
.A(n_1059),
.B(n_885),
.C(n_890),
.D(n_835),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_1051),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1048),
.Y(n_1073)
);

XNOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1055),
.B(n_822),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1049),
.Y(n_1075)
);

NAND4xp75_ASAP7_75t_L g1076 ( 
.A(n_1062),
.B(n_822),
.C(n_890),
.D(n_907),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1050),
.B(n_867),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1052),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1057),
.Y(n_1079)
);

OA22x2_ASAP7_75t_L g1080 ( 
.A1(n_1069),
.A2(n_1056),
.B1(n_1061),
.B2(n_1053),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1072),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_1075),
.B(n_1065),
.Y(n_1082)
);

XNOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1068),
.B(n_1063),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1073),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_1067),
.Y(n_1085)
);

XNOR2xp5_ASAP7_75t_L g1086 ( 
.A(n_1070),
.B(n_1060),
.Y(n_1086)
);

AND4x1_ASAP7_75t_L g1087 ( 
.A(n_1081),
.B(n_1079),
.C(n_1078),
.D(n_1077),
.Y(n_1087)
);

OAI211xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1085),
.A2(n_1074),
.B(n_1071),
.C(n_1076),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1084),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1086),
.B(n_1076),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_1083),
.B(n_1080),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1089),
.B(n_1082),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1091),
.B(n_1087),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1092),
.A2(n_1088),
.B1(n_867),
.B2(n_907),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1094),
.A2(n_811),
.B(n_827),
.Y(n_1096)
);

XNOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1093),
.B(n_836),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1095),
.B(n_811),
.Y(n_1098)
);

AOI222xp33_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_1097),
.B1(n_1096),
.B2(n_882),
.C1(n_901),
.C2(n_893),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1097),
.A2(n_827),
.B(n_833),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1096),
.A2(n_822),
.B(n_882),
.Y(n_1101)
);

AOI222xp33_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_901),
.B1(n_899),
.B2(n_893),
.C1(n_882),
.C2(n_905),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1100),
.B1(n_1099),
.B2(n_907),
.C(n_905),
.Y(n_1103)
);

AOI211xp5_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_899),
.B(n_893),
.C(n_901),
.Y(n_1104)
);


endmodule