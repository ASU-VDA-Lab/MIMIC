module fake_netlist_1_1887_n_877 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_877);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_877;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_769;
wire n_725;
wire n_624;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g104 ( .A(n_94), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_91), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_16), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_7), .B(n_77), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_51), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_74), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_103), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_16), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_67), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_22), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_60), .Y(n_119) );
NOR2xp67_ASAP7_75t_L g120 ( .A(n_72), .B(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_34), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_8), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_21), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_25), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_52), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_42), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_96), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_8), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_65), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_25), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_40), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_35), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
BUFx10_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_6), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_97), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_0), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
INVxp33_ASAP7_75t_L g141 ( .A(n_44), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_57), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_131), .B(n_0), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_126), .B(n_1), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_106), .B(n_1), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_106), .B(n_2), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
BUFx8_ASAP7_75t_SL g150 ( .A(n_118), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_130), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_132), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_130), .B(n_3), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_104), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_109), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_108), .B(n_4), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_108), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
XOR2xp5_ASAP7_75t_L g162 ( .A(n_114), .B(n_5), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_136), .B(n_9), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_113), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_117), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_165), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
OAI22xp33_ASAP7_75t_L g170 ( .A1(n_146), .A2(n_124), .B1(n_122), .B2(n_123), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_153), .B(n_115), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_158), .B(n_115), .Y(n_172) );
XOR2xp5_ASAP7_75t_R g173 ( .A(n_150), .B(n_10), .Y(n_173) );
BUFx8_ASAP7_75t_SL g174 ( .A(n_151), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_153), .A2(n_113), .B1(n_124), .B2(n_122), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_158), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_158), .B(n_110), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_153), .A2(n_123), .B1(n_110), .B2(n_139), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_160), .A2(n_131), .B1(n_107), .B2(n_141), .Y(n_181) );
AND2x6_ASAP7_75t_L g182 ( .A(n_158), .B(n_121), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_149), .B(n_121), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_146), .A2(n_107), .B1(n_116), .B2(n_139), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_151), .B(n_136), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_155), .A2(n_137), .B1(n_139), .B2(n_116), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_156), .B(n_136), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_156), .B(n_125), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_143), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_157), .B(n_105), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_143), .B(n_137), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
INVx5_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_145), .A2(n_137), .B1(n_139), .B2(n_116), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_144), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_163), .B(n_125), .Y(n_207) );
BUFx10_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_147), .A2(n_137), .B1(n_139), .B2(n_116), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g212 ( .A(n_147), .B(n_129), .C(n_140), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_148), .B(n_111), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_205), .B(n_148), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_178), .B(n_127), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_201), .Y(n_217) );
NAND2xp33_ASAP7_75t_L g218 ( .A(n_171), .B(n_127), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_178), .A2(n_159), .B(n_133), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_194), .B(n_159), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_174), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_199), .A2(n_164), .B1(n_160), .B2(n_152), .Y(n_222) );
AOI21x1_ASAP7_75t_L g223 ( .A1(n_187), .A2(n_133), .B(n_129), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_194), .B(n_162), .Y(n_224) );
BUFx5_ASAP7_75t_L g225 ( .A(n_171), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_197), .B(n_162), .Y(n_227) );
AND2x6_ASAP7_75t_SL g228 ( .A(n_173), .B(n_164), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_186), .B(n_112), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_201), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_213), .B(n_128), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_192), .B(n_134), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_187), .B(n_140), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_171), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_171), .A2(n_152), .B1(n_119), .B2(n_138), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_206), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_193), .B(n_142), .Y(n_241) );
NAND2xp33_ASAP7_75t_L g242 ( .A(n_171), .B(n_137), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_191), .B(n_120), .Y(n_243) );
NAND2x1_ASAP7_75t_L g244 ( .A(n_171), .B(n_137), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_171), .A2(n_116), .B1(n_139), .B2(n_165), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_193), .B(n_165), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_193), .B(n_165), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_191), .B(n_161), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_195), .B(n_26), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_193), .B(n_161), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_172), .B(n_161), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_171), .A2(n_166), .B1(n_12), .B2(n_13), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_176), .B(n_27), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_176), .B(n_53), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_200), .B(n_166), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_212), .A2(n_166), .B(n_54), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_172), .B(n_166), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_207), .B(n_175), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_179), .A2(n_166), .B1(n_12), .B2(n_13), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_170), .B(n_55), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_181), .B(n_11), .Y(n_263) );
AOI22xp5_ASAP7_75t_SL g264 ( .A1(n_181), .A2(n_14), .B1(n_15), .B2(n_17), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_212), .B(n_56), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_184), .B(n_14), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_184), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_185), .A2(n_17), .B(n_18), .C(n_19), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_SL g269 ( .A1(n_265), .A2(n_211), .B(n_204), .C(n_190), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_215), .B(n_182), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_252), .A2(n_219), .B(n_216), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_267), .A2(n_182), .B1(n_209), .B2(n_202), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_216), .A2(n_209), .B(n_214), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_214), .B(n_202), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_220), .B(n_182), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_268), .A2(n_189), .B(n_196), .C(n_167), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_260), .B(n_182), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_214), .B(n_202), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_266), .A2(n_182), .B(n_189), .C(n_196), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_224), .B(n_182), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_246), .B(n_182), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_227), .B(n_182), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_226), .A2(n_189), .B(n_196), .C(n_198), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_253), .A2(n_210), .B(n_167), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_259), .A2(n_210), .B(n_167), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_241), .B(n_19), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_251), .A2(n_210), .B(n_180), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_218), .A2(n_208), .B1(n_189), .B2(n_196), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_229), .B(n_20), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_221), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_231), .B(n_20), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_225), .B(n_208), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_225), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_249), .A2(n_183), .B(n_198), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_249), .A2(n_183), .B(n_198), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_221), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_225), .B(n_208), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_222), .B(n_173), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_264), .A2(n_188), .B(n_180), .C(n_183), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_239), .A2(n_238), .B1(n_263), .B2(n_235), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_257), .A2(n_188), .B(n_180), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_218), .A2(n_208), .B1(n_188), .B2(n_169), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_257), .A2(n_169), .B(n_203), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_230), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_234), .A2(n_169), .B(n_22), .C(n_23), .Y(n_308) );
AOI21x1_ASAP7_75t_L g309 ( .A1(n_223), .A2(n_169), .B(n_203), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_232), .B(n_21), .Y(n_310) );
NAND3xp33_ASAP7_75t_L g311 ( .A(n_242), .B(n_245), .C(n_254), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_309), .A2(n_271), .B(n_258), .Y(n_312) );
AO32x2_ASAP7_75t_L g313 ( .A1(n_303), .A2(n_261), .A3(n_243), .B1(n_236), .B2(n_242), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_225), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_277), .A2(n_236), .B(n_238), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_296), .B(n_233), .Y(n_316) );
NAND3x1_ASAP7_75t_L g317 ( .A(n_290), .B(n_228), .C(n_250), .Y(n_317) );
AO31x2_ASAP7_75t_L g318 ( .A1(n_276), .A2(n_255), .A3(n_256), .B(n_240), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_244), .B(n_243), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_299), .B(n_225), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_298), .A2(n_238), .B(n_240), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_275), .A2(n_230), .B(n_237), .Y(n_323) );
O2A1O1Ixp5_ASAP7_75t_L g324 ( .A1(n_310), .A2(n_237), .B(n_225), .C(n_169), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_270), .A2(n_225), .B(n_169), .Y(n_326) );
AOI221x1_ASAP7_75t_L g327 ( .A1(n_302), .A2(n_23), .B1(n_24), .B2(n_28), .C(n_29), .Y(n_327) );
BUFx8_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_280), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_302), .A2(n_203), .B(n_168), .C(n_32), .Y(n_330) );
BUFx8_ASAP7_75t_SL g331 ( .A(n_282), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_307), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_304), .A2(n_30), .B(n_31), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_276), .A2(n_33), .B(n_36), .C(n_37), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
BUFx4_ASAP7_75t_SL g336 ( .A(n_295), .Y(n_336) );
NOR2xp67_ASAP7_75t_SL g337 ( .A(n_295), .B(n_203), .Y(n_337) );
AOI211x1_ASAP7_75t_L g338 ( .A1(n_287), .A2(n_38), .B(n_39), .C(n_41), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_284), .A2(n_43), .B(n_45), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_335), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_332), .B(n_291), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_316), .B(n_291), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_312), .A2(n_285), .B(n_288), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_329), .B(n_281), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_336), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_329), .B(n_308), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_320), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_312), .A2(n_308), .B(n_279), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_317), .B(n_283), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_322), .A2(n_306), .B(n_272), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_278), .B(n_274), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_315), .A2(n_269), .B(n_300), .Y(n_353) );
AO21x2_ASAP7_75t_L g354 ( .A1(n_330), .A2(n_311), .B(n_269), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_323), .B(n_300), .Y(n_355) );
INVx5_ASAP7_75t_L g356 ( .A(n_331), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_317), .B(n_273), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_324), .A2(n_294), .B(n_305), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_338), .B(n_289), .C(n_294), .Y(n_363) );
CKINVDCx11_ASAP7_75t_R g364 ( .A(n_328), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_203), .B(n_168), .Y(n_366) );
AOI21x1_ASAP7_75t_L g367 ( .A1(n_327), .A2(n_46), .B(n_47), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_334), .A2(n_203), .B(n_168), .C(n_50), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_344), .A2(n_322), .B(n_339), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_340), .B(n_318), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_359), .B(n_313), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_345), .B(n_328), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_362), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_367), .A2(n_339), .B(n_333), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_359), .B(n_313), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_349), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_360), .B(n_313), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_340), .B(n_318), .Y(n_380) );
BUFx4f_ASAP7_75t_L g381 ( .A(n_360), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_341), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_357), .Y(n_383) );
AOI21xp33_ASAP7_75t_SL g384 ( .A1(n_365), .A2(n_350), .B(n_346), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
AO21x2_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_333), .B(n_318), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_367), .A2(n_318), .B(n_313), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_343), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_354), .B(n_318), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_354), .B(n_313), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_352), .A2(n_321), .B(n_337), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_48), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_356), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_366), .B(n_348), .Y(n_407) );
BUFx2_ASAP7_75t_SL g408 ( .A(n_356), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_348), .B(n_49), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_364), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_353), .A2(n_331), .B(n_59), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_340), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_358), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_360), .Y(n_415) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_403), .B(n_58), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_382), .B(n_61), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_379), .B(n_62), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_371), .B(n_63), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_411), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_375), .A2(n_66), .B(n_68), .Y(n_423) );
INVx4_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_391), .B(n_69), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_414), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_379), .B(n_70), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_414), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_413), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_414), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_373), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_413), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_371), .B(n_75), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_391), .B(n_78), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_391), .B(n_80), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_374), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_374), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_374), .Y(n_443) );
NAND2x1p5_ASAP7_75t_SL g444 ( .A(n_405), .B(n_81), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_389), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_388), .B(n_85), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_371), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_389), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_377), .B(n_86), .Y(n_452) );
OR2x6_ASAP7_75t_L g453 ( .A(n_408), .B(n_87), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_379), .B(n_89), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_377), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_393), .B(n_90), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_376), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_377), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_394), .B(n_93), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_376), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_388), .B(n_95), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_388), .B(n_99), .Y(n_465) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_400), .B(n_100), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_381), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_397), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_394), .B(n_101), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_390), .B(n_102), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_376), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_397), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_370), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_376), .Y(n_474) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_415), .B(n_168), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_390), .B(n_168), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_370), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_370), .B(n_168), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_372), .B(n_168), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_397), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_405), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_380), .B(n_203), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_380), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_380), .B(n_399), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_378), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_387), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_378), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_387), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_399), .B(n_383), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_384), .A2(n_372), .B(n_410), .C(n_412), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_378), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_387), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_378), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_384), .B(n_409), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_420), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_484), .B(n_410), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_484), .B(n_385), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
OAI21xp5_ASAP7_75t_SL g503 ( .A1(n_490), .A2(n_409), .B(n_403), .Y(n_503) );
NOR2x1p5_ASAP7_75t_L g504 ( .A(n_494), .B(n_405), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_478), .B(n_385), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_478), .B(n_385), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_456), .B(n_411), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_449), .B(n_384), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_426), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_449), .B(n_399), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_424), .A2(n_411), .B1(n_412), .B2(n_409), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_455), .B(n_383), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_455), .B(n_415), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_424), .A2(n_412), .B1(n_409), .B2(n_401), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_426), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g517 ( .A1(n_462), .A2(n_412), .B(n_401), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_430), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_460), .B(n_415), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_460), .B(n_482), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_489), .B(n_398), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_430), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_489), .B(n_398), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_473), .B(n_415), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_450), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_473), .B(n_398), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_477), .B(n_409), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_422), .B(n_409), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_477), .B(n_398), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_483), .B(n_396), .Y(n_530) );
INVx5_ASAP7_75t_L g531 ( .A(n_453), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_461), .B(n_405), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_483), .B(n_401), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_481), .B(n_396), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_481), .B(n_396), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_433), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_461), .B(n_408), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_433), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_461), .B(n_408), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_453), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_486), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_486), .B(n_397), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_420), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_488), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_420), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_488), .B(n_397), .Y(n_546) );
OR2x6_ASAP7_75t_L g547 ( .A(n_453), .B(n_404), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_434), .B(n_406), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_432), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_432), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_432), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_492), .B(n_395), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_442), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_475), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_482), .B(n_381), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_421), .B(n_381), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_442), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_434), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_421), .B(n_412), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_453), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_442), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_443), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_439), .Y(n_564) );
INVx3_ASAP7_75t_L g565 ( .A(n_429), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_443), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_429), .B(n_395), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_436), .B(n_381), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_475), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_453), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_439), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_424), .A2(n_412), .B1(n_381), .B2(n_404), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_443), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_428), .Y(n_574) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_416), .B(n_404), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_428), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_466), .B(n_395), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_436), .B(n_386), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_441), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_452), .B(n_406), .Y(n_580) );
INVx5_ASAP7_75t_L g581 ( .A(n_424), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_459), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_441), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_448), .B(n_406), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_429), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_452), .B(n_386), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_459), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_469), .B(n_386), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_467), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g591 ( .A(n_467), .B(n_395), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_469), .B(n_386), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_467), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_470), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_464), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_419), .B(n_386), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_459), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_448), .B(n_386), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_419), .B(n_392), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_497), .B(n_493), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_582), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_502), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_521), .B(n_493), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_496), .B(n_491), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_491), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_531), .B(n_467), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_520), .B(n_491), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_503), .B(n_479), .C(n_417), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_499), .B(n_487), .Y(n_612) );
OAI33xp33_ASAP7_75t_L g613 ( .A1(n_500), .A2(n_458), .A3(n_438), .B1(n_437), .B2(n_425), .B3(n_476), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_507), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_588), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_523), .B(n_487), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_504), .B(n_472), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_510), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_523), .B(n_487), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_530), .B(n_485), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_531), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_530), .B(n_485), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_498), .B(n_454), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_597), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_509), .B(n_485), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_516), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_511), .B(n_471), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_531), .B(n_466), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_513), .B(n_471), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_518), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_597), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_578), .B(n_474), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_531), .B(n_416), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_581), .Y(n_634) );
INVx4_ASAP7_75t_L g635 ( .A(n_581), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_522), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_474), .Y(n_637) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_550), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_526), .B(n_463), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_529), .B(n_542), .Y(n_640) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_550), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_585), .B(n_463), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_505), .B(n_445), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_506), .B(n_445), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_536), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_542), .B(n_480), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_525), .B(n_427), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_556), .B(n_427), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_495), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_538), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_534), .B(n_445), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_446), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_514), .B(n_446), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_533), .B(n_446), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_508), .B(n_419), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_541), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_594), .B(n_419), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_480), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_544), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_519), .B(n_457), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_551), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_549), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_542), .B(n_480), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_546), .B(n_480), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_551), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_559), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_548), .B(n_454), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
NOR2xp67_ASAP7_75t_L g669 ( .A(n_581), .B(n_472), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_537), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_527), .B(n_457), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_546), .B(n_429), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_524), .B(n_451), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_546), .B(n_468), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_548), .B(n_571), .Y(n_675) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_558), .Y(n_676) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_558), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_580), .B(n_427), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_528), .B(n_427), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_569), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_532), .B(n_451), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_495), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_553), .B(n_472), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_574), .Y(n_684) );
NOR2x1p5_ASAP7_75t_SL g685 ( .A(n_539), .B(n_457), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_553), .B(n_468), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_553), .B(n_468), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_576), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_581), .B(n_512), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_569), .B(n_423), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_543), .B(n_468), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_528), .B(n_454), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_543), .B(n_545), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_545), .B(n_472), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_552), .B(n_451), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_579), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_583), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_593), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_575), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_552), .B(n_454), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_575), .B(n_465), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_532), .B(n_476), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_540), .A2(n_416), .B(n_465), .C(n_464), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_614), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_618), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_626), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_661), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_600), .Y(n_708) );
AND3x2_ASAP7_75t_L g709 ( .A(n_701), .B(n_570), .C(n_561), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_602), .B(n_610), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_640), .B(n_547), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g712 ( .A1(n_703), .A2(n_512), .A3(n_515), .B(n_572), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_630), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_635), .B(n_515), .C(n_517), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_640), .B(n_547), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_636), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_645), .Y(n_717) );
INVxp33_ASAP7_75t_L g718 ( .A(n_635), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_604), .B(n_547), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_611), .A2(n_572), .B1(n_590), .B2(n_595), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_620), .B(n_592), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_670), .B(n_590), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_675), .B(n_589), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_698), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_650), .Y(n_725) );
INVxp67_ASAP7_75t_L g726 ( .A(n_625), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_699), .A2(n_560), .B1(n_568), .B2(n_557), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_632), .B(n_598), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_632), .B(n_587), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_703), .A2(n_577), .B(n_555), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_656), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_605), .B(n_584), .Y(n_732) );
INVxp67_ASAP7_75t_L g733 ( .A(n_606), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_622), .B(n_605), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_659), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_662), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_666), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_629), .B(n_622), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_668), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_637), .B(n_573), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_661), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_612), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_613), .A2(n_555), .B1(n_596), .B2(n_599), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_684), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_655), .B(n_586), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_637), .B(n_554), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_643), .B(n_554), .Y(n_747) );
NAND4xp25_ASAP7_75t_L g748 ( .A(n_689), .B(n_447), .C(n_591), .D(n_577), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_639), .B(n_573), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_648), .B(n_586), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_685), .A2(n_464), .B(n_465), .C(n_565), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_644), .B(n_562), .Y(n_752) );
INVx1_ASAP7_75t_SL g753 ( .A(n_634), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_665), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_635), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_647), .B(n_586), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_688), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_696), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_697), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_607), .B(n_566), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_617), .B(n_565), .Y(n_761) );
AOI32xp33_ASAP7_75t_L g762 ( .A1(n_634), .A2(n_464), .A3(n_465), .B1(n_565), .B2(n_567), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_665), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_607), .B(n_567), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_639), .B(n_566), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_616), .B(n_563), .Y(n_766) );
INVx1_ASAP7_75t_SL g767 ( .A(n_693), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_621), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_616), .B(n_567), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_619), .B(n_563), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_654), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_642), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_660), .Y(n_773) );
INVx1_ASAP7_75t_SL g774 ( .A(n_693), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_619), .Y(n_775) );
OR2x6_ASAP7_75t_L g776 ( .A(n_633), .B(n_608), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_627), .B(n_562), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_742), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_705), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_706), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_726), .B(n_677), .Y(n_781) );
A2O1A1Ixp33_ASAP7_75t_L g782 ( .A1(n_712), .A2(n_633), .B(n_669), .C(n_608), .Y(n_782) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_720), .A2(n_617), .B(n_683), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_713), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_772), .B(n_638), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_708), .A2(n_617), .B(n_683), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_776), .A2(n_628), .B(n_676), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_776), .A2(n_621), .B1(n_680), .B2(n_692), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_773), .B(n_641), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_753), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g791 ( .A1(n_776), .A2(n_621), .B1(n_680), .B2(n_679), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_716), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_717), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_727), .A2(n_708), .B1(n_719), .B2(n_723), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_771), .A2(n_672), .B1(n_663), .B2(n_674), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_755), .A2(n_680), .B1(n_623), .B2(n_663), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_725), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_SL g798 ( .A1(n_712), .A2(n_631), .B(n_682), .C(n_649), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_767), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_730), .A2(n_628), .B(n_690), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_733), .B(n_658), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_731), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_704), .A2(n_678), .B1(n_667), .B2(n_657), .C(n_658), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_735), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_736), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_764), .B(n_674), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g807 ( .A1(n_737), .A2(n_700), .B1(n_695), .B2(n_686), .C1(n_687), .C2(n_682), .Y(n_807) );
AOI222xp33_ASAP7_75t_L g808 ( .A1(n_724), .A2(n_686), .B1(n_687), .B2(n_664), .C1(n_672), .C2(n_700), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_739), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_724), .A2(n_702), .B(n_681), .Y(n_810) );
AOI32xp33_ASAP7_75t_L g811 ( .A1(n_718), .A2(n_664), .A3(n_646), .B1(n_691), .B2(n_694), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_743), .B(n_651), .Y(n_812) );
INVx1_ASAP7_75t_SL g813 ( .A(n_753), .Y(n_813) );
OAI211xp5_ASAP7_75t_SL g814 ( .A1(n_762), .A2(n_652), .B(n_671), .C(n_653), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_755), .A2(n_646), .B1(n_673), .B2(n_609), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_744), .Y(n_816) );
OA21x2_ASAP7_75t_L g817 ( .A1(n_754), .A2(n_609), .B(n_649), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_767), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_757), .Y(n_819) );
OAI322xp33_ASAP7_75t_L g820 ( .A1(n_812), .A2(n_732), .A3(n_774), .B1(n_721), .B2(n_710), .C1(n_728), .C2(n_758), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_782), .A2(n_768), .B1(n_774), .B2(n_751), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_785), .Y(n_822) );
OAI211xp5_ASAP7_75t_SL g823 ( .A1(n_783), .A2(n_714), .B(n_768), .C(n_759), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_817), .Y(n_824) );
OAI21xp33_ASAP7_75t_L g825 ( .A1(n_814), .A2(n_711), .B(n_715), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_789), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_788), .A2(n_714), .B1(n_707), .B2(n_763), .C(n_741), .Y(n_827) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_811), .A2(n_748), .B1(n_729), .B2(n_777), .C(n_765), .Y(n_828) );
OAI21xp33_ASAP7_75t_L g829 ( .A1(n_794), .A2(n_722), .B(n_748), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_791), .A2(n_775), .B1(n_749), .B2(n_746), .C(n_740), .Y(n_830) );
AOI322xp5_ASAP7_75t_L g831 ( .A1(n_786), .A2(n_734), .A3(n_769), .B1(n_750), .B2(n_745), .C1(n_770), .C2(n_756), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_787), .A2(n_738), .B1(n_760), .B2(n_766), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_807), .B(n_761), .Y(n_833) );
AOI21xp33_ASAP7_75t_L g834 ( .A1(n_798), .A2(n_761), .B(n_646), .Y(n_834) );
AOI322xp5_ASAP7_75t_L g835 ( .A1(n_803), .A2(n_796), .A3(n_801), .B1(n_813), .B2(n_790), .C1(n_795), .C2(n_781), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_807), .A2(n_709), .B1(n_747), .B2(n_752), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_778), .B(n_694), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_800), .A2(n_695), .B(n_601), .Y(n_838) );
OAI21xp33_ASAP7_75t_SL g839 ( .A1(n_808), .A2(n_691), .B(n_624), .Y(n_839) );
OAI21xp5_ASAP7_75t_SL g840 ( .A1(n_790), .A2(n_813), .B(n_815), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_799), .B(n_631), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_SL g842 ( .A1(n_810), .A2(n_444), .B(n_615), .C(n_603), .Y(n_842) );
OAI21xp33_ASAP7_75t_SL g843 ( .A1(n_818), .A2(n_624), .B(n_615), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_779), .A2(n_603), .B1(n_601), .B2(n_444), .C(n_423), .Y(n_844) );
AOI211xp5_ASAP7_75t_L g845 ( .A1(n_780), .A2(n_392), .B(n_375), .C(n_444), .Y(n_845) );
AOI21xp33_ASAP7_75t_SL g846 ( .A1(n_817), .A2(n_423), .B(n_407), .Y(n_846) );
O2A1O1Ixp33_ASAP7_75t_L g847 ( .A1(n_784), .A2(n_407), .B(n_402), .C(n_369), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_792), .Y(n_848) );
OAI211xp5_ASAP7_75t_SL g849 ( .A1(n_793), .A2(n_407), .B(n_392), .C(n_402), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g850 ( .A(n_797), .B(n_392), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_802), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_804), .A2(n_375), .B(n_407), .C(n_402), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g853 ( .A(n_805), .B(n_375), .C(n_407), .Y(n_853) );
AOI211xp5_ASAP7_75t_SL g854 ( .A1(n_809), .A2(n_407), .B(n_402), .C(n_369), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_835), .B(n_827), .C(n_829), .D(n_840), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_820), .A2(n_840), .B1(n_823), .B2(n_821), .C(n_839), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_822), .B(n_826), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_825), .B(n_828), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_851), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_838), .B(n_831), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_855), .A2(n_836), .B(n_833), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_858), .B(n_830), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_857), .Y(n_863) );
NOR3xp33_ASAP7_75t_L g864 ( .A(n_856), .B(n_834), .C(n_832), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_863), .Y(n_865) );
NOR4xp25_ASAP7_75t_L g866 ( .A(n_862), .B(n_860), .C(n_824), .D(n_843), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_864), .B(n_842), .C(n_844), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_865), .B(n_861), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_866), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_869), .B(n_867), .Y(n_870) );
AOI21x1_ASAP7_75t_L g871 ( .A1(n_868), .A2(n_859), .B(n_848), .Y(n_871) );
AOI211xp5_ASAP7_75t_L g872 ( .A1(n_870), .A2(n_846), .B(n_845), .C(n_853), .Y(n_872) );
OAI22xp5_ASAP7_75t_SL g873 ( .A1(n_871), .A2(n_819), .B1(n_816), .B2(n_837), .Y(n_873) );
AOI211xp5_ASAP7_75t_L g874 ( .A1(n_873), .A2(n_872), .B(n_847), .C(n_849), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_874), .A2(n_854), .B(n_841), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_875), .A2(n_850), .B1(n_849), .B2(n_852), .C(n_806), .Y(n_876) );
AOI21xp33_ASAP7_75t_SL g877 ( .A1(n_876), .A2(n_402), .B(n_369), .Y(n_877) );
endmodule