module fake_jpeg_1550_n_205 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_205);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_22),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_75),
.B1(n_70),
.B2(n_76),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_88),
.B1(n_78),
.B2(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_62),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx9p33_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_92),
.B1(n_56),
.B2(n_54),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_52),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_48),
.C(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

OR2x4_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_51),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_48),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_110),
.Y(n_111)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_64),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_84),
.C(n_60),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_119),
.C(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_69),
.B1(n_65),
.B2(n_53),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_61),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_59),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_0),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_54),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_44),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_50),
.B1(n_92),
.B2(n_67),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_138),
.B1(n_127),
.B2(n_6),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_140),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_0),
.B(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_6),
.B(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_145),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_25),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_150),
.C(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_24),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_26),
.C(n_43),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_139),
.B(n_153),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_168),
.B(n_13),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_143),
.B1(n_148),
.B2(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_8),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_20),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_31),
.C(n_42),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.C(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.C(n_154),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_18),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_160),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_21),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_159),
.B(n_170),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_191),
.C(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_165),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_157),
.B(n_167),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_164),
.C(n_155),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_158),
.B(n_164),
.Y(n_198)
);

OAI31xp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.A3(n_196),
.B(n_34),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_27),
.C(n_29),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_32),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_37),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_197),
.B(n_39),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_204),
.A2(n_38),
.B(n_41),
.Y(n_205)
);


endmodule