module fake_netlist_6_4605_n_533 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_533);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_533;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_229;
wire n_305;
wire n_532;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_88),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_24),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_85),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_18),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_29),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_17),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_63),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_25),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_38),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_70),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_111),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_67),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_87),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_10),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_78),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_3),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_58),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_36),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_0),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_52),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_75),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_113),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_106),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_53),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_128),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_137),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_11),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_80),
.B(n_73),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_86),
.Y(n_235)
);

OAI22x1_ASAP7_75t_SL g236 ( 
.A1(n_232),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_182),
.A2(n_1),
.B(n_6),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_169),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_8),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_164),
.A2(n_9),
.B(n_14),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_15),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_231),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_19),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_190),
.A2(n_20),
.B(n_21),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_193),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_255)
);

CKINVDCx6p67_ASAP7_75t_R g256 ( 
.A(n_208),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_200),
.A2(n_28),
.B(n_30),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_163),
.B(n_31),
.Y(n_261)
);

XNOR2x2_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_32),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_33),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_154),
.B(n_34),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_188),
.B(n_44),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_219),
.C(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_189),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_225),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_251),
.B(n_159),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_179),
.B1(n_201),
.B2(n_157),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_195),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_197),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_251),
.B(n_179),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_246),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_201),
.B1(n_153),
.B2(n_186),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_158),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_160),
.Y(n_298)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_248),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_241),
.B(n_222),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_256),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_267),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_249),
.B(n_161),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_263),
.A2(n_187),
.B1(n_155),
.B2(n_156),
.Y(n_310)
);

OAI22x1_ASAP7_75t_L g311 ( 
.A1(n_249),
.A2(n_152),
.B1(n_165),
.B2(n_166),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_273),
.A2(n_212),
.B1(n_167),
.B2(n_168),
.Y(n_314)
);

BUFx4f_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_250),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_293),
.B(n_250),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_293),
.B(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_239),
.B1(n_262),
.B2(n_248),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_294),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_255),
.B1(n_265),
.B2(n_272),
.Y(n_323)
);

CKINVDCx11_ASAP7_75t_R g324 ( 
.A(n_295),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_310),
.B(n_162),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_199),
.B1(n_174),
.B2(n_178),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_240),
.B(n_238),
.C(n_253),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_248),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_259),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_199),
.B1(n_181),
.B2(n_183),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_238),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_247),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_240),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_276),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_279),
.B(n_170),
.Y(n_340)
);

OAI221xp5_ASAP7_75t_L g341 ( 
.A1(n_314),
.A2(n_269),
.B1(n_266),
.B2(n_274),
.C(n_253),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_315),
.B(n_234),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_287),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_280),
.B(n_191),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_275),
.A2(n_239),
.B1(n_236),
.B2(n_257),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

NOR3x1_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_214),
.C(n_173),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_287),
.B(n_274),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_287),
.A2(n_239),
.B1(n_257),
.B2(n_252),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_266),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_305),
.B(n_234),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_287),
.B(n_283),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_308),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_315),
.A2(n_192),
.B1(n_194),
.B2(n_207),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_287),
.B(n_245),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_223),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_317),
.B(n_307),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_319),
.B(n_307),
.Y(n_363)
);

O2A1O1Ixp5_ASAP7_75t_L g364 ( 
.A1(n_360),
.A2(n_281),
.B(n_303),
.C(n_312),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_321),
.A2(n_300),
.B1(n_257),
.B2(n_252),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_330),
.Y(n_366)
);

O2A1O1Ixp5_ASAP7_75t_SL g367 ( 
.A1(n_325),
.A2(n_281),
.B(n_176),
.C(n_213),
.Y(n_367)
);

AOI22x1_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_171),
.B1(n_177),
.B2(n_185),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_300),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_278),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_252),
.B(n_302),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_318),
.B(n_224),
.Y(n_373)
);

CKINVDCx11_ASAP7_75t_R g374 ( 
.A(n_324),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_334),
.A2(n_245),
.B(n_209),
.C(n_217),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_309),
.B(n_290),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_300),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_300),
.B1(n_230),
.B2(n_220),
.Y(n_379)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_218),
.B1(n_300),
.B2(n_299),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_361),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_299),
.B(n_46),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_331),
.B(n_328),
.C(n_348),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_341),
.B(n_326),
.C(n_360),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_320),
.A2(n_299),
.B1(n_47),
.B2(n_48),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_333),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_45),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_49),
.Y(n_388)
);

AO32x1_ASAP7_75t_L g389 ( 
.A1(n_349),
.A2(n_50),
.A3(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_356),
.B1(n_355),
.B2(n_345),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_353),
.A2(n_56),
.B(n_57),
.C(n_60),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_61),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_336),
.A2(n_64),
.B(n_65),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_71),
.B(n_74),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_76),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_337),
.B(n_89),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_329),
.B(n_337),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_337),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_SL g403 ( 
.A(n_369),
.B(n_337),
.Y(n_403)
);

NOR4xp25_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_90),
.C(n_92),
.D(n_93),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_94),
.B(n_96),
.C(n_99),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_377),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_100),
.Y(n_407)
);

AO31x2_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_104),
.A3(n_105),
.B(n_109),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_119),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_121),
.B(n_126),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_384),
.A2(n_129),
.B(n_130),
.C(n_131),
.Y(n_412)
);

AOI221xp5_ASAP7_75t_SL g413 ( 
.A1(n_370),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.C(n_140),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_141),
.Y(n_414)
);

AOI221xp5_ASAP7_75t_SL g415 ( 
.A1(n_387),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.C(n_151),
.Y(n_415)
);

AO31x2_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_378),
.A3(n_376),
.B(n_396),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

O2A1O1Ixp33_ASAP7_75t_SL g418 ( 
.A1(n_391),
.A2(n_362),
.B(n_363),
.C(n_388),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_381),
.B(n_390),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_379),
.C(n_386),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_380),
.A2(n_386),
.B1(n_400),
.B2(n_398),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_SL g423 ( 
.A1(n_394),
.A2(n_385),
.B(n_395),
.C(n_389),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_293),
.B1(n_365),
.B2(n_284),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_389),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_389),
.A2(n_365),
.B(n_363),
.Y(n_426)
);

AO31x2_ASAP7_75t_L g427 ( 
.A1(n_375),
.A2(n_370),
.A3(n_383),
.B(n_372),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_382),
.A2(n_372),
.B(n_364),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_374),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_406),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_407),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_405),
.A2(n_412),
.B(n_414),
.C(n_410),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_420),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_411),
.B(n_426),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_402),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_427),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_427),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g439 ( 
.A1(n_425),
.A2(n_415),
.B(n_413),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_401),
.B(n_403),
.C(n_404),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_423),
.B(n_429),
.Y(n_442)
);

BUFx6f_ASAP7_75t_SL g443 ( 
.A(n_421),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_366),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_293),
.B1(n_424),
.B2(n_319),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_438),
.Y(n_448)
);

AO21x2_ASAP7_75t_L g449 ( 
.A1(n_439),
.A2(n_440),
.B(n_435),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_446),
.B(n_436),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_445),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_432),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_444),
.B(n_433),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_434),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

NAND2x1_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_442),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_443),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_452),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_448),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_459),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

NAND2x1_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_451),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_460),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_456),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_450),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_452),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_463),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_472),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_457),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_470),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_475),
.B(n_454),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_457),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_458),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_458),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_458),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_477),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_484),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_474),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_467),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_467),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_490),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_474),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_500),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_497),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_502),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_483),
.B1(n_489),
.B2(n_503),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_502),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_505),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_506),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_489),
.B(n_462),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_498),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_512),
.B(n_501),
.C(n_499),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_511),
.A2(n_494),
.B1(n_492),
.B2(n_496),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_513),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_488),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_460),
.C(n_469),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

NOR2x1_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_460),
.Y(n_520)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_469),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_518),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_522),
.Y(n_524)
);

XOR2x1_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_523),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_524),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_487),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);

AOI221xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_485),
.B1(n_476),
.B2(n_461),
.C(n_449),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_461),
.B1(n_468),
.B2(n_495),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_530),
.B(n_461),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_495),
.B(n_484),
.Y(n_533)
);


endmodule