module fake_jpeg_8902_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_8),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_54),
.Y(n_78)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_66),
.B1(n_33),
.B2(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_69),
.A2(n_46),
.B1(n_24),
.B2(n_32),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_19),
.B(n_61),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_88),
.B2(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_30),
.B1(n_33),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_89),
.B1(n_24),
.B2(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_83),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_21),
.Y(n_111)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_15),
.B(n_14),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_30),
.B1(n_33),
.B2(n_23),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_91),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_17),
.B(n_22),
.C(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_98),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_120),
.B1(n_87),
.B2(n_98),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_97),
.B(n_82),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_49),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_115),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_52),
.B1(n_51),
.B2(n_29),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_95),
.B1(n_87),
.B2(n_70),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_0),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_57),
.B1(n_22),
.B2(n_26),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_24),
.B1(n_32),
.B2(n_27),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_27),
.B1(n_60),
.B2(n_34),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_46),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_70),
.Y(n_131)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

OR2x4_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_27),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_137),
.B(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_147),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_12),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_156),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_0),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_151),
.B(n_154),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_94),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_27),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_25),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_116),
.B(n_102),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_34),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_0),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_34),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_101),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_163),
.C(n_178),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_175),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_128),
.B(n_154),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_108),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_150),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_127),
.B1(n_133),
.B2(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_181),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_49),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_191),
.C(n_143),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_127),
.B(n_100),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_117),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_100),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_172),
.B1(n_161),
.B2(n_190),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_155),
.B1(n_133),
.B2(n_138),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_206),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_183),
.B(n_175),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_154),
.B(n_142),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_204),
.B(n_169),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_128),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_207),
.C(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_156),
.B(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_142),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_141),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_211),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_168),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_160),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_117),
.C(n_112),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_60),
.Y(n_220)
);

OAI22x1_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_174),
.B1(n_170),
.B2(n_162),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_240),
.B1(n_242),
.B2(n_192),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_187),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_207),
.C(n_218),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_238),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_232),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_168),
.B(n_174),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_244),
.B(n_8),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_180),
.B(n_177),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_237),
.B1(n_208),
.B2(n_99),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_183),
.B1(n_185),
.B2(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_205),
.B1(n_211),
.B2(n_194),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_172),
.B1(n_161),
.B2(n_176),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_114),
.B1(n_112),
.B2(n_99),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_9),
.B(n_13),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_99),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_2),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_9),
.B(n_13),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_201),
.B(n_210),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_197),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.C(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_262),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_259),
.B1(n_224),
.B2(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_202),
.B(n_209),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_256),
.B(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_220),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_7),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_8),
.B1(n_11),
.B2(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_6),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_225),
.C(n_227),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_227),
.C(n_222),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_222),
.C(n_230),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_242),
.C(n_221),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_232),
.CI(n_237),
.CON(n_281),
.SN(n_281)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_246),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_235),
.B(n_226),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_282),
.A2(n_252),
.B(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_286),
.B(n_292),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_235),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_274),
.B(n_11),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_257),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_265),
.B(n_255),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_296),
.B(n_279),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_253),
.B(n_259),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_268),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_304),
.C(n_306),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_285),
.A2(n_276),
.B1(n_281),
.B2(n_275),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_293),
.B1(n_291),
.B2(n_3),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_287),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_268),
.C(n_270),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_272),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_281),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_306),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_12),
.B(n_2),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_2),
.B(n_3),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_3),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_303),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_320),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_299),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_305),
.B(n_317),
.C(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_317),
.B(n_322),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_324),
.C(n_326),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_329),
.Y(n_330)
);


endmodule