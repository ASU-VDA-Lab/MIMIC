module real_jpeg_7236_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_43),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_43),
.B1(n_113),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_43),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_142),
.C(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_2),
.B(n_250),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_2),
.A2(n_257),
.B(n_259),
.C(n_260),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_2),
.B(n_270),
.C(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_2),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_2),
.B(n_217),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_22),
.Y(n_296)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_6),
.A2(n_47),
.B1(n_51),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_39),
.B1(n_54),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_6),
.A2(n_54),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_54),
.B1(n_72),
.B2(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_8),
.Y(n_235)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_9),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_10),
.A2(n_81),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_88),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_10),
.A2(n_88),
.B1(n_165),
.B2(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_12),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_354),
.B(n_356),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_144),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_143),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_18),
.B(n_131),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_117),
.B2(n_118),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.C(n_89),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_21),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_21),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_21),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_21),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_21),
.B(n_205),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_21),
.A2(n_136),
.B1(n_182),
.B2(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_21),
.A2(n_136),
.B1(n_253),
.B2(n_263),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_21),
.B(n_174),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_21),
.A2(n_136),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_21),
.A2(n_182),
.B(n_220),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_21),
.A2(n_132),
.B1(n_136),
.B2(n_350),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_32),
.B(n_41),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_28),
.Y(n_141)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_43),
.A2(n_69),
.B(n_72),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_45),
.A2(n_89),
.B1(n_90),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_55),
.B1(n_68),
.B2(n_80),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_46),
.A2(n_55),
.B1(n_68),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_68),
.B(n_80),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AO21x2_ASAP7_75t_SL g152 ( 
.A1(n_56),
.A2(n_68),
.B(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_57)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_68),
.Y(n_250)
);

OA22x2_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_77),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_87),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_89),
.A2(n_90),
.B1(n_138),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_136),
.C(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_111),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_100),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_91),
.A2(n_100),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_100),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_95),
.Y(n_271)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_106),
.B2(n_110),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_101),
.B(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_114),
.Y(n_272)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_130),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_132),
.Y(n_350)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_136),
.A2(n_152),
.B(n_207),
.C(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_137),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_138),
.Y(n_344)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_338),
.B(n_351),
.Y(n_145)
);

OAI211xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_243),
.B(n_332),
.C(n_337),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_225),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_148),
.A2(n_225),
.B(n_333),
.C(n_336),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_208),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_149),
.B(n_208),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_181),
.C(n_193),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_181),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_179),
.B2(n_180),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_151),
.B(n_194),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_151),
.A2(n_179),
.B1(n_232),
.B2(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_214),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_152),
.A2(n_174),
.B1(n_205),
.B2(n_229),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_152),
.A2(n_205),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_153),
.A2(n_204),
.B(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_154),
.A2(n_174),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_161),
.B1(n_167),
.B2(n_171),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_159),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_161),
.B1(n_196),
.B2(n_202),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_174),
.A2(n_229),
.B1(n_249),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_174),
.A2(n_229),
.B1(n_267),
.B2(n_268),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_174),
.A2(n_229),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_174),
.A2(n_205),
.B(n_255),
.C(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_174),
.B(n_205),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_174),
.A2(n_195),
.B1(n_229),
.B2(n_323),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_192),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_186),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_197),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_189),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_204),
.B(n_206),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_195),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_213),
.B(n_218),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_205),
.B(n_240),
.C(n_295),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AND3x1_ASAP7_75t_L g325 ( 
.A(n_207),
.B(n_302),
.C(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_224),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_212),
.B(n_219),
.C(n_224),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

FAx1_ASAP7_75t_L g340 ( 
.A(n_218),
.B(n_341),
.CI(n_345),
.CON(n_340),
.SN(n_340)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_241),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_226),
.B(n_241),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.C(n_231),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_227),
.B(n_228),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_249),
.C(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_292),
.C(n_299),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_231),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_233),
.A2(n_234),
.B1(n_240),
.B2(n_251),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_251),
.B1(n_256),
.B2(n_262),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_240),
.A2(n_251),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_256),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_314),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_304),
.B(n_313),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_290),
.B(n_303),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_264),
.B(n_289),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_263),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_276),
.B(n_288),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_273),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_300),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_327),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_317),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_324),
.C(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_340),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_346),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_348),
.Y(n_353)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_355),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);


endmodule