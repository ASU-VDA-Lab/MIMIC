module fake_netlist_1_2478_n_697 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_36), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_75), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_51), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
INVx3_ASAP7_75t_L g84 ( .A(n_10), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_53), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_54), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_34), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_60), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_37), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_7), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_7), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_74), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_38), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_76), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_43), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_47), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_64), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_50), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_26), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_56), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_31), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_58), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_63), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_35), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_20), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_125), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_125), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_85), .B(n_0), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
NOR2xp33_ASAP7_75t_R g139 ( .A(n_81), .B(n_39), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_113), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_95), .B(n_78), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_85), .B(n_1), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_126), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_121), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_92), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_110), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_87), .A2(n_33), .B(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_87), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_104), .Y(n_153) );
NOR2xp67_ASAP7_75t_L g154 ( .A(n_88), .B(n_3), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_102), .B(n_4), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_109), .B(n_5), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_82), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_92), .A2(n_5), .B1(n_6), .B2(n_9), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_111), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_96), .B(n_11), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_106), .B(n_13), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_119), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_96), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_90), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_89), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_89), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_131), .B(n_105), .Y(n_170) );
OAI21xp33_ASAP7_75t_L g171 ( .A1(n_133), .A2(n_151), .B(n_148), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_152), .B(n_93), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_131), .B(n_126), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_146), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_127), .B(n_124), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_131), .B(n_124), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_127), .B(n_91), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_144), .B(n_116), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_133), .B(n_101), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_135), .B(n_101), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_136), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_143), .B(n_123), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_137), .B(n_112), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_143), .B(n_123), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_149), .B(n_93), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_134), .B(n_94), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_141), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_135), .B(n_122), .Y(n_191) );
AO22x2_ASAP7_75t_L g192 ( .A1(n_137), .A2(n_94), .B1(n_97), .B2(n_98), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_144), .B(n_122), .Y(n_193) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_137), .B(n_120), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_129), .B(n_120), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_140), .B(n_118), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_139), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_167), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_155), .B(n_97), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_167), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_140), .B(n_118), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
BUFx6f_ASAP7_75t_SL g207 ( .A(n_148), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_167), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_132), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_162), .B(n_114), .Y(n_215) );
INVx6_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_151), .B(n_117), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_157), .B(n_98), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_157), .B(n_117), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_136), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_165), .B(n_116), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_226), .Y(n_231) );
BUFx5_ASAP7_75t_L g232 ( .A(n_185), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_219), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_219), .B(n_160), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_184), .B(n_163), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_194), .A2(n_165), .B1(n_166), .B2(n_168), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_194), .B(n_166), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_186), .B(n_153), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_226), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_192), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_215), .B(n_156), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_183), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_213), .Y(n_248) );
NOR3xp33_ASAP7_75t_SL g249 ( .A(n_198), .B(n_147), .C(n_161), .Y(n_249) );
OAI21xp33_ASAP7_75t_SL g250 ( .A1(n_206), .A2(n_159), .B(n_154), .Y(n_250) );
INVx5_ASAP7_75t_L g251 ( .A(n_185), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_209), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_203), .B(n_168), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_213), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_206), .B(n_112), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_185), .B(n_138), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_211), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_185), .A2(n_142), .B1(n_159), .B2(n_154), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_172), .B(n_138), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_190), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_185), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_227), .B(n_138), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_173), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_227), .B(n_138), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
INVx6_ASAP7_75t_L g275 ( .A(n_187), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_171), .B(n_169), .Y(n_276) );
OAI22xp5_ASAP7_75t_SL g277 ( .A1(n_174), .A2(n_99), .B1(n_103), .B2(n_114), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g278 ( .A1(n_174), .A2(n_99), .B1(n_103), .B2(n_150), .Y(n_278) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_188), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_229), .B(n_145), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_229), .B(n_145), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_208), .B(n_214), .Y(n_284) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_180), .B(n_150), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_189), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_220), .B(n_176), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_225), .B(n_169), .Y(n_288) );
INVx6_ASAP7_75t_L g289 ( .A(n_216), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_181), .B(n_158), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_191), .B(n_164), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_199), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_178), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_197), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_287), .A2(n_193), .B(n_178), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_275), .B(n_170), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_245), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_243), .A2(n_244), .B1(n_254), .B2(n_239), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_233), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_276), .A2(n_150), .B(n_193), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_237), .A2(n_222), .B1(n_205), .B2(n_177), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_246), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_275), .B(n_177), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_294), .B(n_196), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_276), .A2(n_175), .B(n_196), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_294), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_230), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_261), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_275), .B(n_175), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_150), .B(n_218), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_272), .B(n_158), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_237), .A2(n_164), .B1(n_108), .B2(n_100), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_272), .B(n_164), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_251), .B(n_115), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_246), .B(n_13), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_232), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_239), .A2(n_224), .B1(n_218), .B2(n_200), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_255), .B(n_14), .Y(n_326) );
NAND2x1_ASAP7_75t_SL g327 ( .A(n_258), .B(n_224), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_231), .B(n_14), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_251), .B(n_217), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_232), .B(n_217), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_238), .B(n_201), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_274), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_259), .A2(n_201), .B(n_200), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_232), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_247), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_241), .B(n_199), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_250), .A2(n_217), .B(n_212), .C(n_210), .Y(n_340) );
BUFx8_ASAP7_75t_L g341 ( .A(n_248), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_281), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_240), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_234), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_232), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_340), .A2(n_262), .B(n_284), .C(n_263), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_330), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_313), .B(n_236), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_313), .B(n_258), .Y(n_350) );
NOR2x1_ASAP7_75t_R g351 ( .A(n_299), .B(n_232), .Y(n_351) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_317), .A2(n_288), .B(n_273), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_309), .B(n_235), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_296), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_279), .B1(n_277), .B2(n_242), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_336), .A2(n_288), .B(n_270), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_336), .A2(n_291), .B(n_282), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_311), .B(n_263), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_303), .A2(n_291), .B(n_283), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_321), .A2(n_279), .B1(n_284), .B2(n_290), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_304), .Y(n_361) );
NOR2xp67_ASAP7_75t_SL g362 ( .A(n_330), .B(n_232), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_315), .B(n_249), .Y(n_363) );
OAI21x1_ASAP7_75t_SL g364 ( .A1(n_331), .A2(n_256), .B(n_265), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_303), .A2(n_257), .B(n_252), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_344), .A2(n_249), .B1(n_235), .B2(n_257), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_327), .A2(n_252), .B(n_264), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_327), .A2(n_264), .B(n_269), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_333), .A2(n_253), .B(n_260), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_310), .B(n_278), .C(n_285), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_335), .B(n_285), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_302), .A2(n_293), .B1(n_247), .B2(n_289), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
AOI221x1_ASAP7_75t_L g376 ( .A1(n_307), .A2(n_217), .B1(n_212), .B2(n_210), .C(n_204), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_326), .A2(n_328), .B(n_305), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_363), .A2(n_316), .B1(n_297), .B2(n_323), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_363), .A2(n_331), .B1(n_307), .B2(n_342), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_346), .A2(n_342), .B1(n_314), .B2(n_301), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_355), .A2(n_314), .B1(n_320), .B2(n_339), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_339), .B1(n_298), .B2(n_305), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_366), .A2(n_349), .B(n_353), .C(n_358), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_346), .B(n_308), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_354), .A2(n_301), .B1(n_298), .B2(n_338), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_360), .A2(n_300), .B(n_338), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_347), .A2(n_312), .B(n_295), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_372), .A2(n_312), .B(n_334), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_325), .B1(n_322), .B2(n_343), .C(n_308), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_361), .B(n_312), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_361), .B(n_343), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_371), .Y(n_393) );
OA21x2_ASAP7_75t_L g394 ( .A1(n_376), .A2(n_319), .B(n_329), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g396 ( .A1(n_354), .A2(n_337), .B1(n_324), .B2(n_341), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_368), .A2(n_341), .B1(n_308), .B2(n_306), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_351), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_374), .A2(n_341), .B(n_345), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_373), .B(n_319), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_373), .B(n_306), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_306), .B1(n_324), .B2(n_337), .C(n_271), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_350), .B(n_289), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_376), .A2(n_332), .B(n_330), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_391), .B(n_359), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_379), .B(n_377), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_392), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_391), .B(n_359), .Y(n_409) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_393), .B(n_348), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_400), .Y(n_411) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_398), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_393), .B(n_348), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_395), .B(n_377), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_377), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_392), .B(n_357), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_401), .B(n_352), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_402), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_388), .B(n_352), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_378), .B(n_352), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_389), .B(n_370), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_389), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_350), .B1(n_364), .B2(n_356), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_389), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_365), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_388), .B(n_365), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_389), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_382), .B(n_356), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_387), .B(n_364), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_389), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_383), .B(n_370), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_394), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_414), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_414), .B(n_394), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_419), .B(n_394), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_419), .B(n_384), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_436), .A2(n_397), .B1(n_386), .B2(n_404), .C(n_399), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_384), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_416), .B(n_386), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_436), .A2(n_385), .B(n_390), .C(n_403), .Y(n_450) );
BUFx8_ASAP7_75t_L g451 ( .A(n_412), .Y(n_451) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_440), .B(n_330), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_424), .B(n_405), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_421), .B(n_367), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_417), .B(n_367), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_369), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_406), .B(n_369), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_412), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_412), .B(n_289), .Y(n_461) );
INVx5_ASAP7_75t_L g462 ( .A(n_426), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_418), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_439), .B(n_421), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_406), .B(n_212), .Y(n_465) );
INVx5_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_406), .B(n_212), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_409), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_410), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_409), .B(n_210), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_410), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_210), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_420), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_425), .B(n_16), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_420), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_422), .B(n_204), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
INVx4_ASAP7_75t_L g483 ( .A(n_410), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_415), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_422), .B(n_204), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_407), .B(n_204), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_413), .Y(n_488) );
INVx5_ASAP7_75t_SL g489 ( .A(n_425), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_449), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_468), .B(n_423), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_460), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_468), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_471), .B(n_423), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_471), .B(n_423), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_441), .B(n_474), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_459), .B(n_429), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_478), .B(n_439), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
NOR2xp33_ASAP7_75t_R g503 ( .A(n_451), .B(n_439), .Y(n_503) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_483), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_474), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_459), .B(n_430), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_454), .B(n_430), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_454), .B(n_430), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_445), .B(n_429), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_477), .B(n_407), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_448), .B(n_427), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_477), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_445), .B(n_429), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_476), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_480), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_447), .B(n_438), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_447), .B(n_438), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_450), .B(n_433), .C(n_435), .D(n_432), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_448), .B(n_434), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_461), .B(n_431), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_451), .B(n_431), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_444), .B(n_438), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_452), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_446), .A2(n_435), .B(n_432), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_480), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_485), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_444), .B(n_437), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_443), .B(n_437), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_488), .B(n_433), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_453), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_459), .B(n_425), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_486), .A2(n_434), .B(n_426), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_443), .B(n_437), .Y(n_534) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_452), .A2(n_428), .A3(n_431), .B(n_425), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_481), .B(n_428), .C(n_425), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_459), .B(n_428), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_17), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
AOI33xp33_ASAP7_75t_L g540 ( .A1(n_453), .A2(n_280), .A3(n_19), .B1(n_21), .B2(n_22), .B3(n_23), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_483), .B(n_469), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_18), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_467), .B(n_25), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_483), .A2(n_332), .B1(n_330), .B2(n_362), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_467), .B(n_27), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_479), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_479), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_501), .B(n_463), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_492), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_490), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_490), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_500), .B(n_489), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_491), .B(n_463), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_531), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_509), .B(n_457), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_509), .B(n_457), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_511), .B(n_455), .C(n_470), .D(n_456), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_491), .B(n_470), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_498), .B(n_457), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_513), .B(n_457), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_500), .B(n_489), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_519), .B(n_451), .C(n_455), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_531), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_546), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_513), .B(n_457), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_497), .B(n_489), .Y(n_567) );
CKINVDCx16_ASAP7_75t_R g568 ( .A(n_503), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_496), .B(n_473), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_532), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_496), .B(n_473), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_502), .B(n_458), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_507), .B(n_489), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_540), .A2(n_475), .B(n_486), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_494), .B(n_484), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_462), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_505), .B(n_484), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_495), .B(n_458), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_514), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_504), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_512), .B(n_482), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_497), .B(n_482), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_520), .B(n_487), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_515), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_495), .B(n_475), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_527), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_541), .B(n_475), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_530), .B(n_487), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_508), .B(n_466), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_495), .B(n_475), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_510), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_530), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_523), .B(n_466), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_528), .B(n_466), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_528), .B(n_534), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_581), .A2(n_535), .B(n_504), .C(n_522), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_563), .A2(n_521), .B1(n_498), .B2(n_506), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_575), .A2(n_525), .B(n_544), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_579), .B(n_498), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_590), .A2(n_524), .B(n_536), .Y(n_605) );
AOI32xp33_ASAP7_75t_L g606 ( .A1(n_550), .A2(n_508), .A3(n_545), .B1(n_543), .B2(n_542), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_568), .A2(n_516), .B1(n_517), .B2(n_537), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_600), .B(n_529), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_595), .A2(n_499), .B1(n_516), .B2(n_517), .C(n_506), .Y(n_610) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_590), .B(n_506), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_595), .B(n_529), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_565), .B(n_462), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_554), .B(n_534), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_572), .A2(n_510), .B1(n_533), .B2(n_537), .C(n_472), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_579), .B(n_532), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_560), .B(n_532), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_572), .A2(n_540), .B(n_469), .C(n_472), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_558), .A2(n_538), .B1(n_545), .B2(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_551), .B(n_547), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_598), .B(n_547), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_552), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_549), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_565), .B(n_518), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_553), .B(n_472), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_586), .B(n_542), .C(n_538), .Y(n_627) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_560), .A2(n_594), .B1(n_593), .B2(n_577), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_588), .B(n_466), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_589), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_592), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g632 ( .A1(n_594), .A2(n_469), .A3(n_466), .B(n_462), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_587), .A2(n_466), .B1(n_462), .B2(n_332), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g635 ( .A1(n_556), .A2(n_462), .A3(n_40), .B1(n_42), .B2(n_45), .C1(n_46), .C2(n_48), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_591), .B(n_462), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_564), .B(n_28), .Y(n_637) );
NAND2x1_ASAP7_75t_SL g638 ( .A(n_613), .B(n_560), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_637), .A2(n_599), .B(n_597), .Y(n_639) );
XNOR2x2_ASAP7_75t_L g640 ( .A(n_627), .B(n_562), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_611), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_602), .A2(n_556), .B1(n_557), .B2(n_561), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_624), .B(n_557), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_620), .A2(n_567), .B1(n_570), .B2(n_559), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_610), .B(n_561), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_630), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_607), .B(n_566), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_631), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_618), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_612), .B(n_570), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_633), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_608), .A2(n_566), .A3(n_569), .B1(n_571), .B2(n_573), .C1(n_570), .C2(n_583), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_601), .A2(n_584), .B(n_582), .C(n_578), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_616), .B(n_584), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_613), .A2(n_576), .B(n_585), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_609), .B(n_580), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_606), .A2(n_580), .B1(n_574), .B2(n_362), .C(n_332), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_621), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_625), .Y(n_660) );
AOI31xp33_ASAP7_75t_L g661 ( .A1(n_644), .A2(n_619), .A3(n_603), .B(n_605), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_651), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_646), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_641), .A2(n_632), .B(n_608), .Y(n_665) );
XNOR2x1_ASAP7_75t_L g666 ( .A(n_641), .B(n_628), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_656), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_653), .A2(n_615), .B(n_629), .C(n_634), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_657), .A2(n_636), .B(n_626), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_644), .A2(n_614), .B(n_622), .C(n_604), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_652), .A2(n_635), .B(n_574), .C(n_617), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_648), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_642), .A2(n_617), .B(n_332), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_655), .A2(n_49), .B(n_52), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_662), .Y(n_675) );
AOI211x1_ASAP7_75t_SL g676 ( .A1(n_674), .A2(n_640), .B(n_645), .C(n_639), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_665), .A2(n_638), .B(n_639), .C(n_660), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_673), .A2(n_650), .B(n_649), .C(n_658), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_666), .B(n_643), .C(n_647), .Y(n_679) );
NAND2xp33_ASAP7_75t_L g680 ( .A(n_661), .B(n_654), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_663), .B(n_55), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_671), .A2(n_57), .B(n_61), .C(n_62), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_680), .B(n_667), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_676), .B(n_670), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_675), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_682), .B(n_671), .C(n_668), .Y(n_686) );
NAND2x1_ASAP7_75t_L g687 ( .A(n_679), .B(n_669), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_685), .Y(n_688) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_686), .B(n_677), .Y(n_689) );
NOR4xp75_ASAP7_75t_L g690 ( .A(n_687), .B(n_681), .C(n_678), .D(n_669), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_688), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_689), .Y(n_692) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_692), .A2(n_684), .B1(n_690), .B2(n_683), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_691), .B(n_672), .C(n_664), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_694), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_695), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_70), .B1(n_71), .B2(n_77), .Y(n_697) );
endmodule