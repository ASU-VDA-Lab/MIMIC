module fake_netlist_5_407_n_2973 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2973);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2973;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2959;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2700;
wire n_2644;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_931;
wire n_870;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_744;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2320;
wire n_2339;
wire n_1045;
wire n_1208;
wire n_2473;
wire n_2038;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2477;
wire n_761;
wire n_2277;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_2953;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_1312;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_2971;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_2722;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_2940;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_2938;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_582),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_207),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_12),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_590),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_546),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_25),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_150),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_194),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_460),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_58),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_3),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_555),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_117),
.Y(n_636)
);

BUFx8_ASAP7_75t_SL g637 ( 
.A(n_182),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_191),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_405),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_600),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_529),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_56),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_324),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_167),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_357),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_357),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_208),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_599),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_601),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_481),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_153),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_336),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_310),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_376),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_188),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_145),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_587),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_277),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_607),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_22),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_352),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_319),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_499),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_83),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_147),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_407),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_439),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_375),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_387),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_236),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_353),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_596),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_452),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_31),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_344),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_171),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_379),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_610),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_87),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_583),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_396),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_347),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_524),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_303),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_512),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_588),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_600),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_443),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_45),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_7),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_53),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_54),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_501),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_135),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_17),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_605),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_207),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_202),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_102),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_612),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_33),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_0),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_9),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_367),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_48),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_285),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_96),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_613),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_23),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_435),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_448),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_259),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_454),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_131),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_557),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_461),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_447),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_44),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_43),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_575),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_31),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_532),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_552),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_216),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_375),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_584),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_80),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_111),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_388),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_280),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_450),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_567),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_243),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_461),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_156),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_330),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_488),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_478),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_268),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_460),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_428),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_459),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_603),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_190),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_274),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_419),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_576),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_575),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_533),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_278),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_38),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_417),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_605),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_218),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_585),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_146),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_526),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_74),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_380),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_480),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_190),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_172),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_104),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_152),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_59),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_76),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_158),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_97),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_261),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_586),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_44),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_137),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_26),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_291),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_598),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_354),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_373),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_322),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_581),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_534),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_568),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_508),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_258),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_214),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_366),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_620),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_488),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_110),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_622),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_145),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_166),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_393),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_589),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_535),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_621),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_53),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_349),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_483),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_290),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_595),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_591),
.Y(n_807)
);

BUFx5_ASAP7_75t_L g808 ( 
.A(n_458),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_592),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_388),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_623),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_17),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_604),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_497),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_608),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_33),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_152),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_330),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_263),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_278),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_316),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_609),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_138),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_401),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_336),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_224),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_602),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_606),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_311),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_105),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_38),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_63),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_293),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_296),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_617),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_80),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_423),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_161),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_570),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_326),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_593),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_76),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_26),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_603),
.Y(n_844)
);

BUFx2_ASAP7_75t_SL g845 ( 
.A(n_109),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_458),
.Y(n_846)
);

BUFx10_ASAP7_75t_L g847 ( 
.A(n_623),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_171),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_15),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_16),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_463),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_594),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_215),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_569),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_528),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_449),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_385),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_11),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_112),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_258),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_325),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_412),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_216),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_509),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_54),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_622),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_173),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_64),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_263),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_371),
.Y(n_870)
);

BUFx5_ASAP7_75t_L g871 ( 
.A(n_111),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_513),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_44),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_637),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_637),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_827),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_650),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_808),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_808),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_808),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_628),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_808),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_808),
.Y(n_885)
);

CKINVDCx16_ASAP7_75t_R g886 ( 
.A(n_630),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_871),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_709),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_631),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_662),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_669),
.Y(n_891)
);

INVxp33_ASAP7_75t_SL g892 ( 
.A(n_629),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_663),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_665),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_871),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_669),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_871),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_650),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_626),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_672),
.Y(n_900)
);

INVxp33_ASAP7_75t_L g901 ( 
.A(n_705),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_871),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_871),
.Y(n_903)
);

CKINVDCx14_ASAP7_75t_R g904 ( 
.A(n_850),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_871),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_871),
.Y(n_906)
);

INVxp33_ASAP7_75t_L g907 ( 
.A(n_873),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_650),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_707),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_674),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_675),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_676),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_707),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_709),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_707),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_626),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_679),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_683),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_630),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_685),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_707),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_688),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_756),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_756),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_689),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_756),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_756),
.Y(n_927)
);

BUFx2_ASAP7_75t_SL g928 ( 
.A(n_747),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_690),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_697),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_701),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_681),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_736),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_633),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_702),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_736),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_681),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_736),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_630),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_650),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_693),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_744),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_694),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_704),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_832),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_725),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_777),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_713),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_816),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_858),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_865),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_713),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_849),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_849),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_832),
.B(n_0),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_708),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_700),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_691),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_643),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_710),
.Y(n_960)
);

CKINVDCx16_ASAP7_75t_R g961 ( 
.A(n_638),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_718),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_643),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_776),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_719),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_703),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_703),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_809),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_726),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_726),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_742),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_724),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_727),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_700),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_742),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_878),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_883),
.B(n_747),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_878),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_883),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_878),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_878),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_889),
.B(n_890),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_878),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_913),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_891),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_889),
.Y(n_986)
);

INVxp33_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_914),
.B(n_700),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_890),
.B(n_677),
.Y(n_989)
);

BUFx2_ASAP7_75t_SL g990 ( 
.A(n_876),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_893),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_908),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_908),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_893),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_940),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_894),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_940),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_896),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_898),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_963),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_932),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_898),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_894),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_898),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_927),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_957),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_957),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_974),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_900),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_974),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_927),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_937),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_900),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_909),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_910),
.B(n_695),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_915),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_910),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_911),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_921),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_911),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_923),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_912),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_942),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_924),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_886),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_902),
.A2(n_698),
.B(n_664),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_912),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_917),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_917),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_918),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_918),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_926),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_945),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_920),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_945),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_920),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_881),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_881),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_903),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_903),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_922),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1005),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1000),
.B(n_933),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1006),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1026),
.B(n_936),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1037),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1026),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1006),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1037),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1038),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1007),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_989),
.A2(n_922),
.B1(n_929),
.B2(n_925),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_L g1053 ( 
.A1(n_1018),
.A2(n_968),
.B1(n_916),
.B2(n_964),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1007),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_1015),
.B(n_919),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1038),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_976),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1008),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_977),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1039),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_976),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1039),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1014),
.B(n_938),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_L g1064 ( 
.A(n_1040),
.B(n_700),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_1040),
.B(n_729),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_984),
.B(n_925),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_983),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1008),
.Y(n_1068)
);

NAND2xp33_ASAP7_75t_L g1069 ( 
.A(n_983),
.B(n_729),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_988),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_978),
.B(n_877),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1010),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1010),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1014),
.B(n_928),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_978),
.A2(n_902),
.B(n_880),
.Y(n_1075)
);

NAND2x1p5_ASAP7_75t_L g1076 ( 
.A(n_999),
.B(n_905),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_992),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_999),
.Y(n_1078)
);

OAI22x1_ASAP7_75t_SL g1079 ( 
.A1(n_985),
.A2(n_786),
.B1(n_842),
.B2(n_744),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1016),
.B(n_953),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1011),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_1002),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_1002),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_990),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_1004),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_1018),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_980),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1016),
.B(n_954),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_982),
.A2(n_929),
.B1(n_931),
.B2(n_930),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_1004),
.A2(n_882),
.B(n_879),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1011),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_992),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_980),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_993),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_993),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_981),
.B(n_884),
.Y(n_1096)
);

AND2x6_ASAP7_75t_L g1097 ( 
.A(n_995),
.B(n_729),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_1019),
.Y(n_1098)
);

CKINVDCx11_ASAP7_75t_R g1099 ( 
.A(n_998),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_995),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_997),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_981),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_997),
.B(n_885),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1019),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_SL g1105 ( 
.A1(n_1001),
.A2(n_842),
.B1(n_844),
.B2(n_786),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_994),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1021),
.B(n_887),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1021),
.Y(n_1108)
);

INVx6_ASAP7_75t_L g1109 ( 
.A(n_1025),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1024),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1024),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_1032),
.A2(n_897),
.B(n_895),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1032),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_987),
.B(n_930),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1033),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1033),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1035),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1030),
.B(n_905),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1041),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_979),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_986),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_991),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_996),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1003),
.B(n_888),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1009),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_SL g1127 ( 
.A1(n_1012),
.A2(n_857),
.B1(n_844),
.B2(n_634),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1013),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1017),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1020),
.B(n_906),
.Y(n_1130)
);

INVxp33_ASAP7_75t_SL g1131 ( 
.A(n_1022),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_1125),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1115),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1066),
.A2(n_1028),
.B1(n_1029),
.B2(n_1027),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1109),
.B(n_990),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_1114),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1130),
.A2(n_892),
.B1(n_958),
.B2(n_939),
.Y(n_1137)
);

AO22x2_ASAP7_75t_L g1138 ( 
.A1(n_1055),
.A2(n_699),
.B1(n_723),
.B2(n_845),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1074),
.B(n_904),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1074),
.B(n_901),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1119),
.B(n_916),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1125),
.B(n_907),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1125),
.B(n_1031),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1115),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1043),
.A2(n_1036),
.B1(n_1034),
.B2(n_931),
.Y(n_1145)
);

OAI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1120),
.A2(n_961),
.B1(n_944),
.B2(n_956),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1115),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1070),
.B(n_935),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1077),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1086),
.B(n_934),
.Y(n_1150)
);

AO22x2_ASAP7_75t_L g1151 ( 
.A1(n_1120),
.A2(n_657),
.B1(n_670),
.B2(n_654),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1077),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1095),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1043),
.A2(n_935),
.B1(n_956),
.B2(n_944),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1086),
.B(n_960),
.Y(n_1155)
);

OA22x2_ASAP7_75t_L g1156 ( 
.A1(n_1053),
.A2(n_962),
.B1(n_965),
.B2(n_960),
.Y(n_1156)
);

AO22x2_ASAP7_75t_L g1157 ( 
.A1(n_1122),
.A2(n_1123),
.B1(n_1128),
.B2(n_1124),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1080),
.B(n_941),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1121),
.B(n_962),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1109),
.B(n_914),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1052),
.A2(n_965),
.B1(n_973),
.B2(n_972),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1121),
.B(n_972),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1124),
.B(n_973),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1089),
.A2(n_906),
.B1(n_874),
.B2(n_875),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1095),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1122),
.A2(n_788),
.B1(n_789),
.B2(n_768),
.Y(n_1166)
);

AND2x2_ASAP7_75t_SL g1167 ( 
.A(n_1126),
.B(n_955),
.Y(n_1167)
);

AO22x2_ASAP7_75t_L g1168 ( 
.A1(n_1123),
.A2(n_853),
.B1(n_860),
.B2(n_841),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1059),
.B(n_874),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1106),
.B(n_875),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_857),
.B1(n_966),
.B2(n_959),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1056),
.A2(n_967),
.B1(n_970),
.B2(n_969),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1105),
.A2(n_1023),
.B1(n_634),
.B2(n_642),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1045),
.Y(n_1174)
);

NOR2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1084),
.B(n_963),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1110),
.A2(n_955),
.B1(n_872),
.B2(n_862),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1045),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_1079),
.A2(n_928),
.B1(n_698),
.B2(n_730),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1115),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1049),
.A2(n_975),
.B1(n_971),
.B2(n_946),
.Y(n_1180)
);

NOR2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1084),
.B(n_888),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1111),
.A2(n_730),
.B1(n_755),
.B2(n_664),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1049),
.A2(n_947),
.B1(n_949),
.B2(n_943),
.Y(n_1183)
);

OAI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1131),
.A2(n_642),
.B1(n_661),
.B2(n_633),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1045),
.Y(n_1185)
);

AO22x2_ASAP7_75t_L g1186 ( 
.A1(n_1053),
.A2(n_794),
.B1(n_803),
.B2(n_755),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1109),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1131),
.B(n_1050),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1115),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1109),
.A2(n_843),
.B1(n_868),
.B2(n_661),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1126),
.B(n_948),
.Y(n_1191)
);

AO22x2_ASAP7_75t_L g1192 ( 
.A1(n_1127),
.A2(n_803),
.B1(n_837),
.B2(n_794),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1126),
.B(n_952),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1126),
.B(n_952),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1075),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1117),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1100),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1117),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1050),
.A2(n_950),
.B1(n_951),
.B2(n_948),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1060),
.A2(n_1062),
.B1(n_1108),
.B2(n_1100),
.Y(n_1200)
);

NAND3x1_ASAP7_75t_L g1201 ( 
.A(n_1063),
.B(n_666),
.C(n_651),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1126),
.B(n_798),
.Y(n_1202)
);

OA22x2_ASAP7_75t_L g1203 ( 
.A1(n_1080),
.A2(n_868),
.B1(n_843),
.B2(n_640),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1060),
.A2(n_837),
.B1(n_706),
.B2(n_722),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1062),
.A2(n_1082),
.B1(n_1085),
.B2(n_1083),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1047),
.A2(n_627),
.B1(n_646),
.B2(n_625),
.Y(n_1206)
);

OA22x2_ASAP7_75t_L g1207 ( 
.A1(n_1080),
.A2(n_644),
.B1(n_624),
.B2(n_635),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1117),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1129),
.B(n_638),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1082),
.A2(n_731),
.B1(n_734),
.B2(n_732),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1075),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1082),
.A2(n_737),
.B1(n_741),
.B2(n_738),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1083),
.B(n_696),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1092),
.Y(n_1214)
);

AO22x2_ASAP7_75t_L g1215 ( 
.A1(n_1047),
.A2(n_647),
.B1(n_655),
.B2(n_648),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1113),
.A2(n_779),
.B1(n_802),
.B2(n_770),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1108),
.B(n_729),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1063),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1113),
.Y(n_1219)
);

AO22x2_ASAP7_75t_L g1220 ( 
.A1(n_1088),
.A2(n_656),
.B1(n_667),
.B2(n_660),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1129),
.B(n_638),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1129),
.B(n_658),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1083),
.A2(n_748),
.B1(n_749),
.B2(n_745),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1117),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1099),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1108),
.B(n_1085),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1116),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1129),
.B(n_658),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1092),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1117),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1088),
.A2(n_673),
.B1(n_678),
.B2(n_671),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1085),
.B(n_774),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1044),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1088),
.A2(n_831),
.B1(n_812),
.B2(n_632),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1129),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1078),
.B(n_870),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1116),
.A2(n_632),
.B1(n_635),
.B2(n_624),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1093),
.A2(n_1104),
.B1(n_1118),
.B2(n_1101),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_752),
.B1(n_754),
.B2(n_750),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1118),
.B(n_658),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1094),
.B(n_855),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1094),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1042),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1101),
.B(n_774),
.Y(n_1244)
);

OAI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1107),
.A2(n_639),
.B1(n_640),
.B2(n_636),
.Y(n_1245)
);

AOI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1076),
.A2(n_639),
.B1(n_641),
.B2(n_636),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_1098),
.A2(n_680),
.B1(n_684),
.B2(n_682),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1042),
.B(n_867),
.Y(n_1248)
);

AO22x2_ASAP7_75t_L g1249 ( 
.A1(n_1098),
.A2(n_686),
.B1(n_692),
.B2(n_687),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_1076),
.B1(n_1103),
.B2(n_1071),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1104),
.A2(n_712),
.B1(n_714),
.B2(n_711),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1048),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_SL g1253 ( 
.A(n_1098),
.B(n_668),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1048),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_758),
.B1(n_759),
.B2(n_757),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1076),
.A2(n_717),
.B1(n_720),
.B2(n_716),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1096),
.A2(n_763),
.B1(n_764),
.B2(n_761),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1112),
.A2(n_766),
.B1(n_771),
.B2(n_765),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1112),
.A2(n_780),
.B1(n_782),
.B2(n_778),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1051),
.A2(n_728),
.B1(n_733),
.B2(n_721),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1087),
.B(n_784),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1051),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1057),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1057),
.B(n_774),
.Y(n_1264)
);

AO22x2_ASAP7_75t_L g1265 ( 
.A1(n_1054),
.A2(n_739),
.B1(n_740),
.B2(n_735),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1112),
.A2(n_792),
.B1(n_793),
.B2(n_787),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1112),
.A2(n_796),
.B1(n_797),
.B2(n_795),
.Y(n_1267)
);

NAND3x1_ASAP7_75t_L g1268 ( 
.A(n_1064),
.B(n_818),
.C(n_769),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1090),
.B(n_668),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1174),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1136),
.B(n_1087),
.Y(n_1271)
);

BUFx8_ASAP7_75t_SL g1272 ( 
.A(n_1135),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1174),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1132),
.B(n_798),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1177),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1132),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1185),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1185),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1214),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1141),
.B(n_1087),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1142),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1187),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1214),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1135),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1229),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1229),
.Y(n_1287)
);

AND2x6_ASAP7_75t_L g1288 ( 
.A(n_1211),
.B(n_1057),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1242),
.Y(n_1289)
);

NOR3xp33_ASAP7_75t_L g1290 ( 
.A(n_1137),
.B(n_1184),
.C(n_1146),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1242),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1134),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1233),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1150),
.B(n_840),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1235),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1193),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1263),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1211),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1154),
.B(n_804),
.C(n_801),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_R g1300 ( 
.A(n_1155),
.B(n_1148),
.Y(n_1300)
);

AND2x6_ASAP7_75t_L g1301 ( 
.A(n_1195),
.B(n_1057),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1188),
.B(n_1087),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1149),
.B(n_1087),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1227),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1252),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1254),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1194),
.B(n_1158),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1160),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1167),
.B(n_1102),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1218),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1160),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1219),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1262),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1152),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1140),
.B(n_1102),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1153),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1159),
.B(n_1102),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1143),
.B(n_840),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1165),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1263),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1202),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1197),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1133),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1139),
.B(n_1162),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1171),
.A2(n_1241),
.B1(n_1203),
.B2(n_1145),
.Y(n_1326)
);

BUFx4f_ASAP7_75t_L g1327 ( 
.A(n_1202),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1243),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1191),
.B(n_856),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1163),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_L g1331 ( 
.A(n_1226),
.B(n_1057),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1158),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1200),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1161),
.B(n_810),
.C(n_805),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1195),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1209),
.B(n_856),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1144),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1221),
.B(n_668),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1232),
.A2(n_1090),
.B(n_1073),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1238),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_1181),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1222),
.B(n_715),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1147),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1228),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1244),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_1175),
.Y(n_1346)
);

AND2x6_ASAP7_75t_L g1347 ( 
.A(n_1269),
.B(n_1061),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_L g1348 ( 
.A(n_1240),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1179),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1213),
.B(n_1102),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1248),
.B(n_715),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1157),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1205),
.B(n_1061),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1225),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1189),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1196),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1198),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1208),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1250),
.B(n_1061),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1224),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1210),
.B(n_813),
.C(n_811),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1230),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1261),
.B(n_1102),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1206),
.A2(n_1090),
.B1(n_743),
.B2(n_753),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1217),
.Y(n_1365)
);

NOR2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1236),
.B(n_641),
.Y(n_1366)
);

BUFx4f_ASAP7_75t_L g1367 ( 
.A(n_1157),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1265),
.Y(n_1368)
);

BUFx10_ASAP7_75t_L g1369 ( 
.A(n_1169),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1265),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1258),
.A2(n_1058),
.B1(n_1068),
.B2(n_1054),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1264),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1245),
.B(n_1061),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1199),
.B(n_1058),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1237),
.B(n_1061),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1207),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1259),
.B(n_1090),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1268),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1220),
.B(n_751),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1266),
.B(n_1067),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1180),
.Y(n_1381)
);

BUFx8_ASAP7_75t_SL g1382 ( 
.A(n_1173),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1183),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1206),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1267),
.B(n_1067),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1215),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1138),
.B(n_1067),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1215),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1190),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1201),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1220),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1138),
.B(n_1067),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1231),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1231),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1251),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1186),
.A2(n_762),
.B1(n_767),
.B2(n_760),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1186),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1182),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_SL g1400 ( 
.A(n_1253),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1156),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1256),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1212),
.B(n_1067),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1164),
.A2(n_1072),
.B1(n_1073),
.B2(n_1068),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1246),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1246),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1151),
.B(n_715),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1260),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1151),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1234),
.B(n_1072),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1223),
.B(n_1081),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1257),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1239),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1247),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1247),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1176),
.B(n_1081),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1255),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1178),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1204),
.B(n_1091),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1216),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1249),
.B(n_1091),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1166),
.A2(n_772),
.B1(n_781),
.B2(n_773),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1166),
.Y(n_1423)
);

NAND2xp33_ASAP7_75t_L g1424 ( 
.A(n_1168),
.B(n_1065),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1168),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1178),
.B(n_644),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1192),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1192),
.B(n_814),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1132),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1174),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_SL g1431 ( 
.A(n_1135),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1174),
.Y(n_1432)
);

XOR2xp5_ASAP7_75t_L g1433 ( 
.A(n_1225),
.B(n_815),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1174),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1174),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1136),
.B(n_817),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1174),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1174),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1174),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1174),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1174),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1136),
.B(n_819),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1132),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1174),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1174),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1167),
.B(n_774),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1142),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1173),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1149),
.B(n_1065),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1235),
.B(n_645),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1195),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1174),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1174),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1174),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1174),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1167),
.B(n_790),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1167),
.A2(n_1065),
.B1(n_1097),
.B2(n_1064),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1174),
.Y(n_1458)
);

BUFx8_ASAP7_75t_SL g1459 ( 
.A(n_1135),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1132),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1174),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1149),
.B(n_1065),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1132),
.B(n_785),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1154),
.B(n_822),
.C(n_820),
.Y(n_1464)
);

AND2x2_ASAP7_75t_SL g1465 ( 
.A(n_1167),
.B(n_790),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1174),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1142),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1458),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1333),
.B(n_790),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1429),
.B(n_790),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_L g1472 ( 
.A(n_1436),
.B(n_1069),
.C(n_800),
.Y(n_1472)
);

BUFx4_ASAP7_75t_L g1473 ( 
.A(n_1427),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1330),
.B(n_825),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1467),
.B(n_1325),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1315),
.B(n_799),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1466),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1429),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1466),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1289),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1289),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1275),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1279),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1430),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1354),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1276),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1278),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1272),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1434),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1397),
.A2(n_791),
.B1(n_823),
.B2(n_824),
.C(n_821),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1437),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1315),
.B(n_799),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1300),
.A2(n_1097),
.B1(n_1069),
.B2(n_828),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1307),
.B(n_1296),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1307),
.B(n_830),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1348),
.B(n_1465),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1439),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1317),
.B(n_799),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1317),
.B(n_799),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1432),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1441),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1444),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1397),
.A2(n_851),
.B1(n_854),
.B2(n_846),
.C(n_836),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1348),
.B(n_826),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1310),
.B(n_806),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1300),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1296),
.B(n_861),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1277),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1436),
.B(n_829),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1410),
.A2(n_1097),
.B1(n_834),
.B2(n_833),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1295),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1465),
.A2(n_807),
.B1(n_806),
.B2(n_863),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1332),
.B(n_864),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1452),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1453),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1461),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1435),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1438),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1454),
.Y(n_1519)
);

AND2x6_ASAP7_75t_L g1520 ( 
.A(n_1298),
.B(n_806),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1282),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1314),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1314),
.Y(n_1523)
);

BUFx4f_ASAP7_75t_L g1524 ( 
.A(n_1336),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1273),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1332),
.B(n_866),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1270),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1277),
.B(n_869),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1310),
.B(n_806),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1273),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1440),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1443),
.B(n_807),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1447),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1294),
.B(n_645),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1440),
.Y(n_1535)
);

BUFx10_ASAP7_75t_L g1536 ( 
.A(n_1431),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1443),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1283),
.Y(n_1538)
);

INVx8_ASAP7_75t_L g1539 ( 
.A(n_1431),
.Y(n_1539)
);

AND3x4_ASAP7_75t_L g1540 ( 
.A(n_1290),
.B(n_775),
.C(n_746),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1318),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1445),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1398),
.A2(n_807),
.B1(n_775),
.B2(n_783),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1316),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1460),
.B(n_807),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1283),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1316),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1460),
.B(n_65),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1445),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1271),
.B(n_1097),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1455),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1455),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1284),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1286),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1352),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1287),
.Y(n_1556)
);

INVx8_ASAP7_75t_L g1557 ( 
.A(n_1463),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1442),
.B(n_1412),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1280),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1344),
.B(n_65),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1291),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1376),
.B(n_66),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1304),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1318),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1320),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1295),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1311),
.B(n_66),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1410),
.A2(n_1097),
.B1(n_652),
.B2(n_653),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1295),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1442),
.B(n_649),
.Y(n_1570)
);

BUFx4_ASAP7_75t_L g1571 ( 
.A(n_1423),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1311),
.B(n_67),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1323),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1272),
.Y(n_1574)
);

AO22x2_ASAP7_75t_L g1575 ( 
.A1(n_1425),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1389),
.B(n_649),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1401),
.B(n_67),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1270),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1312),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1459),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1306),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1459),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1352),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1306),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1295),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1367),
.B(n_1097),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1271),
.B(n_652),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1298),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1367),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1356),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1292),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1322),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1356),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1370),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1293),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1337),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1305),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1313),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1408),
.B(n_653),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1324),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1324),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1281),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1281),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1349),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1338),
.B(n_1342),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1302),
.B(n_659),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1343),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1328),
.B(n_68),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1355),
.Y(n_1609)
);

AND2x6_ASAP7_75t_L g1610 ( 
.A(n_1340),
.B(n_1),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1357),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1341),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1358),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1395),
.B(n_68),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1341),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1360),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1351),
.B(n_746),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1362),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1303),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1368),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1417),
.A2(n_835),
.B1(n_838),
.B2(n_659),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1309),
.A2(n_838),
.B1(n_839),
.B2(n_835),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1335),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1297),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1297),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1319),
.B(n_1384),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1336),
.B(n_746),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1408),
.B(n_839),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1408),
.B(n_848),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1387),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1391),
.B(n_69),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1318),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1285),
.B(n_69),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1336),
.B(n_775),
.Y(n_1634)
);

NAND2x1p5_ASAP7_75t_L g1635 ( 
.A(n_1285),
.B(n_70),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1337),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1408),
.A2(n_852),
.B1(n_855),
.B2(n_848),
.Y(n_1637)
);

AO22x2_ASAP7_75t_L g1638 ( 
.A1(n_1386),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1329),
.B(n_852),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1346),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1321),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1346),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1327),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1321),
.Y(n_1644)
);

BUFx4_ASAP7_75t_L g1645 ( 
.A(n_1400),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1404),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1339),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1326),
.B(n_859),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1372),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1391),
.B(n_70),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1399),
.A2(n_867),
.B1(n_870),
.B2(n_859),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1463),
.B(n_71),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1327),
.Y(n_1653)
);

CKINVDCx8_ASAP7_75t_R g1654 ( 
.A(n_1421),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1302),
.B(n_2),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1372),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1374),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1308),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1309),
.B(n_3),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1374),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1319),
.B(n_783),
.Y(n_1661)
);

INVx8_ASAP7_75t_L g1662 ( 
.A(n_1463),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1329),
.B(n_783),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1393),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1359),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1371),
.Y(n_1666)
);

AO22x2_ASAP7_75t_L g1667 ( 
.A1(n_1384),
.A2(n_1409),
.B1(n_1415),
.B2(n_1414),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1301),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1345),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1365),
.Y(n_1670)
);

NOR2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1390),
.B(n_847),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1369),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1326),
.B(n_847),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1419),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1594),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1558),
.B(n_1420),
.Y(n_1676)
);

BUFx12f_ASAP7_75t_L g1677 ( 
.A(n_1536),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1527),
.B(n_1416),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1527),
.B(n_1413),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1602),
.B(n_1402),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1602),
.B(n_1419),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1509),
.A2(n_1406),
.B1(n_1290),
.B2(n_1366),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1539),
.B(n_1308),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1603),
.B(n_1396),
.Y(n_1684)
);

AND2x6_ASAP7_75t_L g1685 ( 
.A(n_1589),
.B(n_1390),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1603),
.B(n_1416),
.Y(n_1686)
);

INVxp33_ASAP7_75t_L g1687 ( 
.A(n_1475),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1619),
.B(n_1646),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1669),
.B(n_1446),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_SL g1690 ( 
.A1(n_1570),
.A2(n_1373),
.B(n_1375),
.C(n_1405),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1591),
.B(n_1605),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1555),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1570),
.B(n_1334),
.C(n_1361),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1494),
.B(n_1394),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1538),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1506),
.B(n_1329),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1506),
.B(n_1576),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1468),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1606),
.B(n_1383),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1496),
.A2(n_1406),
.B1(n_1448),
.B2(n_1400),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1648),
.A2(n_1394),
.B1(n_1464),
.B2(n_1299),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1494),
.B(n_1388),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1606),
.B(n_1587),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1673),
.A2(n_1448),
.B1(n_1433),
.B2(n_1415),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1587),
.B(n_1381),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1657),
.B(n_1392),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1630),
.B(n_1456),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1594),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1546),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1479),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1508),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1673),
.A2(n_1418),
.B1(n_1450),
.B2(n_1373),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1471),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1658),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1630),
.B(n_1456),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1643),
.B(n_1421),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1555),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1477),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1578),
.B(n_1446),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1563),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1508),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1565),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1576),
.B(n_1617),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1659),
.B(n_1648),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1474),
.B(n_1388),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1659),
.B(n_1364),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1621),
.A2(n_1379),
.B1(n_1426),
.B2(n_1274),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1664),
.B(n_1350),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1621),
.A2(n_1379),
.B1(n_1274),
.B2(n_1378),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1674),
.B(n_1411),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1654),
.B(n_1428),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1660),
.A2(n_1379),
.B1(n_1424),
.B2(n_1428),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1665),
.A2(n_1363),
.B(n_1451),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1665),
.B(n_1364),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1507),
.B(n_1407),
.Y(n_1735)
);

OAI22x1_ASAP7_75t_L g1736 ( 
.A1(n_1540),
.A2(n_1457),
.B1(n_1422),
.B2(n_1424),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1573),
.B(n_1422),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1666),
.B(n_1347),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1588),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1599),
.B(n_1369),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1512),
.A2(n_1589),
.B1(n_1620),
.B2(n_1554),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1522),
.B(n_1347),
.Y(n_1742)
);

AND2x2_ASAP7_75t_SL g1743 ( 
.A(n_1524),
.B(n_1512),
.Y(n_1743)
);

NOR2xp67_ASAP7_75t_L g1744 ( 
.A(n_1653),
.B(n_1403),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_L g1745 ( 
.A(n_1672),
.B(n_1347),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1507),
.B(n_1274),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1628),
.A2(n_1347),
.B1(n_1385),
.B2(n_1380),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1553),
.Y(n_1748)
);

OAI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1622),
.A2(n_1524),
.B1(n_1653),
.B2(n_1534),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1485),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1629),
.B(n_1382),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1480),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1661),
.A2(n_1347),
.B1(n_1385),
.B2(n_1377),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1592),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1643),
.B(n_1451),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1504),
.A2(n_1331),
.B1(n_1353),
.B2(n_1359),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1482),
.B(n_1365),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1643),
.B(n_1672),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1486),
.B(n_1365),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1626),
.A2(n_1331),
.B1(n_1353),
.B2(n_1449),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1655),
.A2(n_1462),
.B(n_847),
.C(n_72),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1487),
.B(n_1365),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1508),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1663),
.A2(n_1288),
.B1(n_1301),
.B2(n_1451),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1489),
.B(n_1451),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1610),
.A2(n_1288),
.B1(n_1301),
.B2(n_6),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1543),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1481),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1491),
.B(n_1288),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1511),
.B(n_1301),
.Y(n_1770)
);

NOR3x1_ASAP7_75t_L g1771 ( 
.A(n_1541),
.B(n_1632),
.C(n_1564),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_SL g1772 ( 
.A(n_1536),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1610),
.A2(n_1288),
.B1(n_1301),
.B2(n_7),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1589),
.B(n_71),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1614),
.B(n_1495),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1497),
.B(n_4),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1537),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1537),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1514),
.B(n_5),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1610),
.A2(n_9),
.B1(n_5),
.B2(n_8),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1515),
.B(n_8),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1516),
.B(n_8),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1579),
.B(n_9),
.Y(n_1784)
);

O2A1O1Ixp5_ASAP7_75t_L g1785 ( 
.A1(n_1655),
.A2(n_1499),
.B(n_1498),
.C(n_1476),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1583),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1583),
.B(n_10),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1498),
.A2(n_73),
.B(n_72),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1627),
.A2(n_74),
.B1(n_75),
.B2(n_73),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1523),
.B(n_10),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1537),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1511),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1672),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1640),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1521),
.B(n_75),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1495),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1533),
.B(n_77),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1544),
.B(n_11),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1547),
.B(n_12),
.Y(n_1799)
);

AO22x1_ASAP7_75t_L g1800 ( 
.A1(n_1652),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1639),
.Y(n_1801)
);

INVx5_ASAP7_75t_L g1802 ( 
.A(n_1668),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1637),
.B(n_1651),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1566),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1548),
.B(n_77),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1614),
.B(n_611),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1517),
.B(n_1519),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1637),
.B(n_78),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1581),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1590),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1596),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1556),
.B(n_13),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1528),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1548),
.B(n_78),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1559),
.B(n_1561),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1670),
.B(n_1525),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1528),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1651),
.B(n_79),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1513),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1634),
.A2(n_81),
.B1(n_82),
.B2(n_79),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1640),
.B(n_81),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_SL g1822 ( 
.A1(n_1499),
.A2(n_17),
.B(n_14),
.C(n_16),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1638),
.A2(n_1543),
.B1(n_1575),
.B2(n_1568),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1631),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1483),
.B(n_16),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1566),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1530),
.B(n_18),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1597),
.B(n_82),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1640),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1593),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1484),
.B(n_18),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1667),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1584),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1598),
.B(n_1595),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1608),
.B(n_618),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1566),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1490),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.C(n_21),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1645),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1513),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1839)
);

NOR2xp67_ASAP7_75t_L g1840 ( 
.A(n_1478),
.B(n_20),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1631),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1671),
.A2(n_84),
.B1(n_85),
.B2(n_83),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1526),
.B(n_84),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1500),
.B(n_1518),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1649),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1642),
.B(n_85),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1604),
.B(n_19),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1505),
.B(n_21),
.Y(n_1848)
);

INVx5_ASAP7_75t_L g1849 ( 
.A(n_1668),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1526),
.B(n_86),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1531),
.B(n_22),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1656),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1535),
.B(n_86),
.Y(n_1853)
);

INVxp67_ASAP7_75t_SL g1854 ( 
.A(n_1596),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1667),
.A2(n_1608),
.B1(n_1545),
.B2(n_1532),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1609),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1642),
.B(n_87),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1539),
.B(n_88),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1642),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1611),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1532),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1567),
.A2(n_89),
.B1(n_90),
.B2(n_88),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1539),
.B(n_89),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1613),
.Y(n_1864)
);

INVxp33_ASAP7_75t_L g1865 ( 
.A(n_1545),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1542),
.B(n_23),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1692),
.Y(n_1867)
);

INVx5_ASAP7_75t_L g1868 ( 
.A(n_1685),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1703),
.B(n_1650),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1778),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1723),
.B(n_1650),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1779),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1750),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1720),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1711),
.Y(n_1875)
);

INVx2_ASAP7_75t_SL g1876 ( 
.A(n_1695),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1693),
.A2(n_1803),
.B(n_1724),
.C(n_1682),
.Y(n_1877)
);

AND2x6_ASAP7_75t_L g1878 ( 
.A(n_1764),
.B(n_1569),
.Y(n_1878)
);

BUFx12f_ASAP7_75t_L g1879 ( 
.A(n_1677),
.Y(n_1879)
);

BUFx12f_ASAP7_75t_L g1880 ( 
.A(n_1838),
.Y(n_1880)
);

OR2x2_ASAP7_75t_SL g1881 ( 
.A(n_1676),
.B(n_1571),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1709),
.Y(n_1882)
);

AND2x4_ASAP7_75t_SL g1883 ( 
.A(n_1721),
.B(n_1478),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1697),
.B(n_1633),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1786),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1722),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1699),
.B(n_1616),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1818),
.A2(n_1575),
.B1(n_1638),
.B2(n_1652),
.Y(n_1888)
);

INVx4_ASAP7_75t_L g1889 ( 
.A(n_1778),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1807),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1856),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1748),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1678),
.B(n_1469),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1808),
.A2(n_1560),
.B1(n_1577),
.B2(n_1562),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1705),
.B(n_1577),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1687),
.B(n_1572),
.Y(n_1896)
);

O2A1O1Ixp5_ASAP7_75t_L g1897 ( 
.A1(n_1788),
.A2(n_1476),
.B(n_1492),
.C(n_1550),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1860),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1778),
.Y(n_1899)
);

NOR2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1794),
.B(n_1580),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1864),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1791),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1686),
.B(n_1562),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1829),
.Y(n_1904)
);

INVx4_ASAP7_75t_L g1905 ( 
.A(n_1791),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1698),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1833),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1691),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1739),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1713),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1859),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1725),
.B(n_1572),
.Y(n_1912)
);

AO22x1_ASAP7_75t_L g1913 ( 
.A1(n_1823),
.A2(n_1788),
.B1(n_1685),
.B2(n_1774),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_SL g1914 ( 
.A(n_1743),
.B(n_1557),
.Y(n_1914)
);

INVxp67_ASAP7_75t_SL g1915 ( 
.A(n_1679),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1791),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1718),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1752),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1717),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1729),
.A2(n_1560),
.B1(n_1503),
.B2(n_1568),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1802),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1768),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1710),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1824),
.Y(n_1924)
);

BUFx8_ASAP7_75t_L g1925 ( 
.A(n_1772),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1815),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1772),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_R g1928 ( 
.A(n_1754),
.B(n_1488),
.Y(n_1928)
);

OR2x2_ASAP7_75t_SL g1929 ( 
.A(n_1841),
.B(n_1472),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1845),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1696),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1815),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1731),
.A2(n_1510),
.B1(n_1635),
.B2(n_1633),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1736),
.A2(n_1701),
.B1(n_1767),
.B2(n_1837),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1804),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1749),
.B(n_1635),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1683),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1804),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1763),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1940)
);

BUFx5_ASAP7_75t_L g1941 ( 
.A(n_1685),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1775),
.Y(n_1942)
);

INVx5_ASAP7_75t_L g1943 ( 
.A(n_1685),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1852),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1702),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1804),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1809),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1727),
.A2(n_1662),
.B1(n_1557),
.B2(n_1472),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1810),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1793),
.Y(n_1950)
);

INVx5_ASAP7_75t_L g1951 ( 
.A(n_1802),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1830),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1675),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1708),
.Y(n_1954)
);

AO22x1_ASAP7_75t_L g1955 ( 
.A1(n_1771),
.A2(n_1582),
.B1(n_1615),
.B2(n_1612),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1844),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1802),
.B(n_1607),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1827),
.Y(n_1958)
);

NOR2xp67_ASAP7_75t_L g1959 ( 
.A(n_1802),
.B(n_1618),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1694),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1686),
.B(n_1688),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1688),
.B(n_1662),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1827),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1851),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1816),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1851),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1866),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1801),
.A2(n_1551),
.B1(n_1552),
.B2(n_1549),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1706),
.B(n_1505),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1679),
.B(n_1469),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1683),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1716),
.B(n_1569),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1728),
.B(n_1529),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1714),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1757),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1759),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_L g1977 ( 
.A(n_1707),
.B(n_1715),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1813),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1721),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1866),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1849),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1762),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1704),
.B(n_1636),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1735),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1806),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1777),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1683),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1684),
.B(n_1600),
.Y(n_1988)
);

INVx4_ASAP7_75t_L g1989 ( 
.A(n_1777),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1834),
.Y(n_1990)
);

AND3x2_ASAP7_75t_SL g1991 ( 
.A(n_1858),
.B(n_1473),
.C(n_1623),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1790),
.Y(n_1992)
);

OR2x6_ASAP7_75t_L g1993 ( 
.A(n_1744),
.B(n_1470),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1798),
.Y(n_1994)
);

AND2x6_ASAP7_75t_SL g1995 ( 
.A(n_1751),
.B(n_1574),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1712),
.A2(n_1493),
.B1(n_1601),
.B2(n_1625),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1858),
.A2(n_1493),
.B1(n_1636),
.B2(n_1470),
.Y(n_1997)
);

BUFx12f_ASAP7_75t_L g1998 ( 
.A(n_1863),
.Y(n_1998)
);

INVx5_ASAP7_75t_L g1999 ( 
.A(n_1849),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1689),
.Y(n_2000)
);

BUFx12f_ASAP7_75t_L g2001 ( 
.A(n_1863),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1781),
.A2(n_1644),
.B1(n_1520),
.B2(n_1641),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1863),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1700),
.B(n_1624),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1680),
.B(n_1492),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1689),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1746),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1681),
.Y(n_2008)
);

INVxp67_ASAP7_75t_SL g2009 ( 
.A(n_1811),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1799),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1740),
.B(n_1569),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1758),
.B(n_1585),
.Y(n_2012)
);

BUFx3_ASAP7_75t_L g2013 ( 
.A(n_1836),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_L g2014 ( 
.A(n_1737),
.B(n_1585),
.Y(n_2014)
);

INVx5_ASAP7_75t_L g2015 ( 
.A(n_1849),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1681),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_L g2017 ( 
.A(n_1766),
.B(n_1585),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1835),
.B(n_1843),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1812),
.Y(n_2019)
);

INVxp67_ASAP7_75t_SL g2020 ( 
.A(n_1854),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1836),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1765),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1812),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1797),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1730),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1680),
.B(n_1647),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1776),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1817),
.Y(n_2028)
);

AND3x1_ASAP7_75t_L g2029 ( 
.A(n_1842),
.B(n_1550),
.C(n_24),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1865),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1730),
.B(n_1728),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1849),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1792),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1826),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1780),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1882),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1960),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1933),
.B(n_1732),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2031),
.B(n_1848),
.Y(n_2039)
);

BUFx4f_ASAP7_75t_L g2040 ( 
.A(n_1960),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1874),
.Y(n_2041)
);

CKINVDCx6p67_ASAP7_75t_R g2042 ( 
.A(n_1873),
.Y(n_2042)
);

OA22x2_ASAP7_75t_L g2043 ( 
.A1(n_1888),
.A2(n_1789),
.B1(n_1862),
.B2(n_1814),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1886),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_2014),
.A2(n_1733),
.B(n_1734),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1933),
.B(n_1990),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1915),
.A2(n_1734),
.B(n_1785),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_2024),
.B(n_1805),
.Y(n_2048)
);

O2A1O1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_1877),
.A2(n_1846),
.B(n_1857),
.C(n_1821),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1892),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2025),
.B(n_1726),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_SL g2052 ( 
.A1(n_1881),
.A2(n_1820),
.B1(n_1796),
.B2(n_1819),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1897),
.A2(n_1738),
.B(n_1747),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1969),
.A2(n_1690),
.B(n_1741),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1928),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1869),
.B(n_1855),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1971),
.B(n_1832),
.Y(n_2057)
);

O2A1O1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_1884),
.A2(n_1795),
.B(n_1822),
.C(n_1761),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1936),
.A2(n_1850),
.B1(n_1773),
.B2(n_1839),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1898),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1983),
.A2(n_1741),
.B(n_1784),
.C(n_1783),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2029),
.A2(n_1828),
.B1(n_1853),
.B2(n_1800),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1925),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1903),
.B(n_1719),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1961),
.B(n_1782),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1891),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1895),
.B(n_1861),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_1960),
.Y(n_2068)
);

A2O1A1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_1920),
.A2(n_1756),
.B(n_1753),
.C(n_1840),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2008),
.B(n_1825),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1970),
.A2(n_1745),
.B(n_1738),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1970),
.A2(n_1742),
.B(n_1760),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2016),
.B(n_1831),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1907),
.Y(n_2074)
);

BUFx8_ASAP7_75t_L g2075 ( 
.A(n_1879),
.Y(n_2075)
);

OA22x2_ASAP7_75t_L g2076 ( 
.A1(n_1894),
.A2(n_1920),
.B1(n_1948),
.B2(n_1962),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1906),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1909),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1951),
.A2(n_1742),
.B(n_1769),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2027),
.B(n_1847),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1871),
.B(n_1787),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1914),
.B(n_1792),
.Y(n_2082)
);

OAI22x1_ASAP7_75t_L g2083 ( 
.A1(n_1948),
.A2(n_1894),
.B1(n_1931),
.B2(n_2019),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1899),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1914),
.B(n_1755),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_1912),
.B(n_1826),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1925),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1930),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1899),
.Y(n_2089)
);

AOI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_1951),
.A2(n_2015),
.B(n_1999),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1953),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1934),
.A2(n_1586),
.B(n_1770),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1910),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2035),
.B(n_1872),
.Y(n_2094)
);

OAI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_2022),
.A2(n_1586),
.B(n_1770),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1951),
.A2(n_1520),
.B(n_617),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_SL g2097 ( 
.A1(n_2004),
.A2(n_1520),
.B(n_26),
.C(n_24),
.Y(n_2097)
);

O2A1O1Ixp33_ASAP7_75t_SL g2098 ( 
.A1(n_1997),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_2098)
);

O2A1O1Ixp33_ASAP7_75t_L g2099 ( 
.A1(n_1992),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_2099)
);

OAI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2029),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2100)
);

O2A1O1Ixp33_ASAP7_75t_L g2101 ( 
.A1(n_1994),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_SL g2102 ( 
.A(n_1927),
.B(n_32),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1913),
.A2(n_40),
.B1(n_49),
.B2(n_32),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1984),
.B(n_90),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1944),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1974),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_2007),
.Y(n_2107)
);

A2O1A1Ixp33_ASAP7_75t_L g2108 ( 
.A1(n_2017),
.A2(n_92),
.B(n_93),
.C(n_91),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1887),
.B(n_91),
.Y(n_2109)
);

NOR3xp33_ASAP7_75t_L g2110 ( 
.A(n_2011),
.B(n_33),
.C(n_34),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_1937),
.Y(n_2111)
);

OA22x2_ASAP7_75t_L g2112 ( 
.A1(n_2003),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_1999),
.A2(n_614),
.B(n_613),
.Y(n_2113)
);

AOI22x1_ASAP7_75t_L g2114 ( 
.A1(n_2010),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1975),
.B(n_92),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1976),
.B(n_93),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1982),
.B(n_94),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1868),
.B(n_34),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1999),
.A2(n_620),
.B(n_619),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_2015),
.A2(n_1893),
.B(n_1973),
.Y(n_2120)
);

O2A1O1Ixp33_ASAP7_75t_L g2121 ( 
.A1(n_2023),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1958),
.B(n_95),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1987),
.B(n_97),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2007),
.B(n_98),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_2015),
.A2(n_99),
.B(n_98),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1868),
.B(n_99),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1931),
.B(n_100),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1963),
.B(n_100),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_SL g2129 ( 
.A(n_1868),
.B(n_37),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1964),
.B(n_101),
.Y(n_2130)
);

OR2x6_ASAP7_75t_L g2131 ( 
.A(n_1993),
.B(n_101),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1901),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_1908),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1893),
.A2(n_614),
.B(n_612),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_1890),
.B(n_102),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1973),
.A2(n_616),
.B(n_615),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1943),
.B(n_103),
.Y(n_2137)
);

INVx4_ASAP7_75t_L g2138 ( 
.A(n_1943),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_1985),
.B(n_103),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1985),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1929),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2005),
.A2(n_621),
.B(n_619),
.Y(n_2142)
);

BUFx3_ASAP7_75t_L g2143 ( 
.A(n_1911),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1943),
.B(n_104),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2028),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1966),
.B(n_105),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1942),
.B(n_106),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1967),
.B(n_106),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1917),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_1867),
.B(n_1919),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2045),
.A2(n_2026),
.B(n_2006),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_2057),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2143),
.Y(n_2153)
);

OA22x2_ASAP7_75t_L g2154 ( 
.A1(n_2062),
.A2(n_1980),
.B1(n_1954),
.B2(n_1991),
.Y(n_2154)
);

AOI211x1_ASAP7_75t_L g2155 ( 
.A1(n_2133),
.A2(n_2100),
.B(n_2145),
.C(n_2141),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_2053),
.A2(n_2000),
.B(n_1981),
.Y(n_2156)
);

AOI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2090),
.A2(n_1959),
.B(n_1957),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2132),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_2047),
.A2(n_1959),
.B(n_1957),
.Y(n_2159)
);

OAI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_2069),
.A2(n_1977),
.B(n_1996),
.Y(n_2160)
);

OAI21x1_ASAP7_75t_L g2161 ( 
.A1(n_2054),
.A2(n_1981),
.B(n_1921),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2062),
.A2(n_1954),
.B1(n_2002),
.B2(n_1885),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_2120),
.A2(n_2020),
.B(n_2009),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_2042),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2081),
.B(n_2018),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2046),
.B(n_2030),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2039),
.B(n_1926),
.Y(n_2167)
);

OAI21x1_ASAP7_75t_L g2168 ( 
.A1(n_2079),
.A2(n_1921),
.B(n_2032),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2091),
.B(n_1932),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_2036),
.Y(n_2170)
);

AND2x6_ASAP7_75t_SL g2171 ( 
.A(n_2048),
.B(n_1896),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_2072),
.A2(n_2032),
.B(n_1996),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2071),
.A2(n_1993),
.B(n_1988),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2041),
.B(n_1965),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2103),
.A2(n_1968),
.B1(n_2001),
.B2(n_1998),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_L g2176 ( 
.A1(n_2095),
.A2(n_1922),
.B(n_1918),
.Y(n_2176)
);

OA21x2_ASAP7_75t_L g2177 ( 
.A1(n_2038),
.A2(n_1947),
.B(n_1923),
.Y(n_2177)
);

OAI21x1_ASAP7_75t_L g2178 ( 
.A1(n_2061),
.A2(n_2092),
.B(n_2096),
.Y(n_2178)
);

OAI21x1_ASAP7_75t_L g2179 ( 
.A1(n_2149),
.A2(n_1952),
.B(n_1949),
.Y(n_2179)
);

OAI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2058),
.A2(n_1993),
.B(n_1924),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_2076),
.A2(n_2033),
.B(n_1956),
.Y(n_2181)
);

INVx4_ASAP7_75t_L g2182 ( 
.A(n_2138),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2044),
.B(n_1878),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_2036),
.Y(n_2184)
);

OAI21x1_ASAP7_75t_L g2185 ( 
.A1(n_2082),
.A2(n_1900),
.B(n_1941),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_2093),
.A2(n_1941),
.B(n_1878),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2050),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2060),
.B(n_1878),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_2049),
.A2(n_1940),
.B(n_1945),
.C(n_1978),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2098),
.A2(n_2051),
.B(n_2097),
.Y(n_2190)
);

AOI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2085),
.A2(n_1972),
.B(n_1940),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_2036),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2057),
.B(n_2012),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2074),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2066),
.A2(n_1941),
.B(n_1878),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2150),
.B(n_1876),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2078),
.B(n_2064),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_2084),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2103),
.A2(n_1972),
.B1(n_2012),
.B2(n_1939),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_2084),
.Y(n_2200)
);

OAI21x1_ASAP7_75t_SL g2201 ( 
.A1(n_2121),
.A2(n_1989),
.B(n_1889),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2108),
.A2(n_1875),
.B(n_1904),
.Y(n_2202)
);

INVx4_ASAP7_75t_L g2203 ( 
.A(n_2138),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_2111),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_2142),
.A2(n_1916),
.B(n_1950),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_2077),
.A2(n_1941),
.B(n_1889),
.Y(n_2206)
);

NAND2x1_ASAP7_75t_L g2207 ( 
.A(n_2131),
.B(n_1989),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2088),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2105),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2094),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2118),
.A2(n_1941),
.B(n_1883),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2065),
.B(n_2107),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2083),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2086),
.B(n_1995),
.Y(n_2214)
);

OAI21x1_ASAP7_75t_L g2215 ( 
.A1(n_2136),
.A2(n_2113),
.B(n_2119),
.Y(n_2215)
);

BUFx2_ASAP7_75t_SL g2216 ( 
.A(n_2084),
.Y(n_2216)
);

NOR2xp67_ASAP7_75t_L g2217 ( 
.A(n_2106),
.B(n_1880),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_2125),
.A2(n_1905),
.B(n_1870),
.Y(n_2218)
);

OAI22x1_ASAP7_75t_L g2219 ( 
.A1(n_2213),
.A2(n_2114),
.B1(n_2124),
.B2(n_2109),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2152),
.B(n_2131),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2210),
.B(n_2197),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2160),
.A2(n_2043),
.B1(n_2052),
.B2(n_2110),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2187),
.Y(n_2223)
);

AO31x2_ASAP7_75t_L g2224 ( 
.A1(n_2159),
.A2(n_2134),
.A3(n_2056),
.B(n_2140),
.Y(n_2224)
);

AO31x2_ASAP7_75t_L g2225 ( 
.A1(n_2173),
.A2(n_2128),
.A3(n_2130),
.B(n_2122),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2194),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2178),
.A2(n_2116),
.B(n_2115),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_2196),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_L g2229 ( 
.A1(n_2172),
.A2(n_2117),
.B(n_2146),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2177),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2214),
.B(n_1995),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2158),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2197),
.B(n_2127),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2169),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_2180),
.B(n_2070),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2160),
.A2(n_2129),
.B(n_2131),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_SL g2237 ( 
.A1(n_2154),
.A2(n_2195),
.B(n_2186),
.Y(n_2237)
);

NAND3xp33_ASAP7_75t_L g2238 ( 
.A(n_2205),
.B(n_2101),
.C(n_2099),
.Y(n_2238)
);

INVx1_ASAP7_75t_SL g2239 ( 
.A(n_2153),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2155),
.A2(n_2059),
.B1(n_2112),
.B2(n_2126),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2212),
.B(n_2169),
.Y(n_2241)
);

OAI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2215),
.A2(n_2144),
.B(n_2137),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2154),
.A2(n_2067),
.B1(n_2148),
.B2(n_2139),
.Y(n_2243)
);

CKINVDCx12_ASAP7_75t_R g2244 ( 
.A(n_2165),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2212),
.B(n_2073),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_2161),
.A2(n_2068),
.B(n_2037),
.Y(n_2246)
);

CKINVDCx11_ASAP7_75t_R g2247 ( 
.A(n_2171),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_2173),
.A2(n_2068),
.B(n_2037),
.Y(n_2248)
);

A2O1A1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2189),
.A2(n_2102),
.B(n_2147),
.C(n_2104),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_SL g2250 ( 
.A(n_2164),
.B(n_2063),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2174),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2166),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_SL g2253 ( 
.A(n_2211),
.B(n_2087),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2204),
.B(n_2080),
.Y(n_2254)
);

INVx5_ASAP7_75t_L g2255 ( 
.A(n_2182),
.Y(n_2255)
);

NOR2xp67_ASAP7_75t_L g2256 ( 
.A(n_2163),
.B(n_2135),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_2152),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2167),
.B(n_2123),
.Y(n_2258)
);

AOI31xp67_ASAP7_75t_L g2259 ( 
.A1(n_2183),
.A2(n_2123),
.A3(n_2089),
.B(n_2040),
.Y(n_2259)
);

AO31x2_ASAP7_75t_L g2260 ( 
.A1(n_2163),
.A2(n_2199),
.A3(n_2203),
.B(n_2182),
.Y(n_2260)
);

AO32x2_ASAP7_75t_L g2261 ( 
.A1(n_2199),
.A2(n_1870),
.A3(n_1905),
.B1(n_1955),
.B2(n_2089),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2167),
.B(n_2089),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2230),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2260),
.B(n_2206),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2241),
.B(n_2166),
.Y(n_2265)
);

AOI22x1_ASAP7_75t_L g2266 ( 
.A1(n_2219),
.A2(n_2190),
.B1(n_2211),
.B2(n_2205),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2252),
.B(n_2209),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2223),
.Y(n_2268)
);

INVx4_ASAP7_75t_SL g2269 ( 
.A(n_2260),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2226),
.Y(n_2270)
);

AND2x2_ASAP7_75t_SL g2271 ( 
.A(n_2253),
.B(n_2177),
.Y(n_2271)
);

AOI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2236),
.A2(n_2190),
.B(n_2180),
.Y(n_2272)
);

OAI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_2238),
.A2(n_2175),
.B1(n_2207),
.B2(n_2191),
.Y(n_2273)
);

OAI21x1_ASAP7_75t_L g2274 ( 
.A1(n_2248),
.A2(n_2156),
.B(n_2151),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2260),
.B(n_2185),
.Y(n_2275)
);

OA21x2_ASAP7_75t_L g2276 ( 
.A1(n_2227),
.A2(n_2168),
.B(n_2176),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2246),
.A2(n_2229),
.B(n_2157),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2222),
.A2(n_2247),
.B1(n_2243),
.B2(n_2240),
.Y(n_2278)
);

CKINVDCx20_ASAP7_75t_R g2279 ( 
.A(n_2244),
.Y(n_2279)
);

AO31x2_ASAP7_75t_L g2280 ( 
.A1(n_2234),
.A2(n_2188),
.A3(n_2183),
.B(n_2203),
.Y(n_2280)
);

OAI21x1_ASAP7_75t_L g2281 ( 
.A1(n_2242),
.A2(n_2188),
.B(n_2181),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2232),
.Y(n_2282)
);

OAI21x1_ASAP7_75t_L g2283 ( 
.A1(n_2235),
.A2(n_2179),
.B(n_2174),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2251),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2225),
.Y(n_2285)
);

INVx1_ASAP7_75t_SL g2286 ( 
.A(n_2239),
.Y(n_2286)
);

A2O1A1Ixp33_ASAP7_75t_L g2287 ( 
.A1(n_2249),
.A2(n_2202),
.B(n_2175),
.C(n_2162),
.Y(n_2287)
);

OAI21x1_ASAP7_75t_L g2288 ( 
.A1(n_2256),
.A2(n_2191),
.B(n_2218),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2271),
.B(n_2228),
.Y(n_2289)
);

BUFx8_ASAP7_75t_L g2290 ( 
.A(n_2266),
.Y(n_2290)
);

BUFx12f_ASAP7_75t_L g2291 ( 
.A(n_2271),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2272),
.A2(n_2231),
.B(n_2256),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2271),
.B(n_2269),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2263),
.Y(n_2294)
);

NOR2xp67_ASAP7_75t_L g2295 ( 
.A(n_2285),
.B(n_2237),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2270),
.Y(n_2296)
);

BUFx12f_ASAP7_75t_SL g2297 ( 
.A(n_2279),
.Y(n_2297)
);

OR2x6_ASAP7_75t_L g2298 ( 
.A(n_2288),
.B(n_2259),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2291),
.A2(n_2266),
.B1(n_2278),
.B2(n_2273),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2296),
.Y(n_2300)
);

OA222x2_ASAP7_75t_L g2301 ( 
.A1(n_2298),
.A2(n_2269),
.B1(n_2263),
.B2(n_2285),
.C1(n_2261),
.C2(n_2257),
.Y(n_2301)
);

AO22x1_ASAP7_75t_L g2302 ( 
.A1(n_2290),
.A2(n_2075),
.B1(n_2255),
.B2(n_2286),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2294),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2293),
.B(n_2269),
.Y(n_2304)
);

BUFx12f_ASAP7_75t_L g2305 ( 
.A(n_2290),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2297),
.B(n_2250),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_2305),
.Y(n_2307)
);

AO21x2_ASAP7_75t_L g2308 ( 
.A1(n_2301),
.A2(n_2295),
.B(n_2292),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2300),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2304),
.B(n_2293),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2303),
.Y(n_2311)
);

AOI22xp33_ASAP7_75t_L g2312 ( 
.A1(n_2299),
.A2(n_2291),
.B1(n_2290),
.B2(n_2289),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2304),
.B(n_2298),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2303),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_2306),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2302),
.B(n_2289),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2310),
.B(n_2305),
.Y(n_2317)
);

INVx5_ASAP7_75t_L g2318 ( 
.A(n_2307),
.Y(n_2318)
);

BUFx2_ASAP7_75t_L g2319 ( 
.A(n_2307),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2310),
.B(n_2302),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2314),
.Y(n_2321)
);

AND2x2_ASAP7_75t_SL g2322 ( 
.A(n_2312),
.B(n_2297),
.Y(n_2322)
);

INVx1_ASAP7_75t_SL g2323 ( 
.A(n_2307),
.Y(n_2323)
);

AND2x4_ASAP7_75t_SL g2324 ( 
.A(n_2316),
.B(n_2298),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2316),
.B(n_2300),
.Y(n_2325)
);

BUFx12f_ASAP7_75t_L g2326 ( 
.A(n_2313),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2314),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2319),
.B(n_2315),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2317),
.B(n_2315),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2317),
.B(n_2313),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2321),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2319),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2320),
.B(n_2313),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2318),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2326),
.Y(n_2335)
);

INVx2_ASAP7_75t_SL g2336 ( 
.A(n_2318),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2332),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2336),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2333),
.B(n_2320),
.Y(n_2339)
);

NAND2x1_ASAP7_75t_SL g2340 ( 
.A(n_2329),
.B(n_2325),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2339),
.B(n_2333),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2339),
.B(n_2329),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2337),
.B(n_2328),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_2340),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2341),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2342),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2343),
.B(n_2332),
.Y(n_2347)
);

INVx1_ASAP7_75t_SL g2348 ( 
.A(n_2344),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2341),
.B(n_2323),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2341),
.B(n_2330),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2350),
.B(n_2318),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2347),
.B(n_2338),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2345),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2348),
.B(n_2318),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2346),
.B(n_2330),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2348),
.B(n_2338),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2349),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2347),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2350),
.B(n_2335),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2347),
.Y(n_2360)
);

NOR2x1_ASAP7_75t_L g2361 ( 
.A(n_2356),
.B(n_2360),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_2352),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2355),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2360),
.Y(n_2364)
);

OR2x2_ASAP7_75t_L g2365 ( 
.A(n_2358),
.B(n_2335),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2359),
.B(n_2318),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2353),
.B(n_2318),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2357),
.B(n_2322),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2354),
.B(n_2351),
.Y(n_2369)
);

HB1xp67_ASAP7_75t_L g2370 ( 
.A(n_2352),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2356),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2356),
.B(n_2336),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2355),
.B(n_2322),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2361),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2373),
.B(n_2322),
.Y(n_2375)
);

INVx1_ASAP7_75t_SL g2376 ( 
.A(n_2362),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2370),
.B(n_2331),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2361),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2364),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2372),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2368),
.B(n_2326),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2371),
.B(n_2334),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2365),
.B(n_2334),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2363),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2367),
.Y(n_2385)
);

OAI21xp33_ASAP7_75t_L g2386 ( 
.A1(n_2366),
.A2(n_2331),
.B(n_2327),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2369),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2361),
.Y(n_2388)
);

A2O1A1Ixp33_ASAP7_75t_L g2389 ( 
.A1(n_2374),
.A2(n_2327),
.B(n_2321),
.C(n_2324),
.Y(n_2389)
);

OAI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_2376),
.A2(n_2325),
.B1(n_2326),
.B2(n_2311),
.C(n_2309),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2381),
.B(n_2380),
.Y(n_2391)
);

NOR3xp33_ASAP7_75t_L g2392 ( 
.A(n_2387),
.B(n_2075),
.C(n_2055),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2375),
.B(n_2308),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2383),
.B(n_2308),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2378),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2384),
.A2(n_2324),
.B1(n_2308),
.B2(n_2309),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2382),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2379),
.B(n_2324),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2388),
.B(n_2308),
.Y(n_2399)
);

INVx1_ASAP7_75t_SL g2400 ( 
.A(n_2377),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2386),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2386),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2399),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2394),
.Y(n_2404)
);

OAI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2392),
.A2(n_2385),
.B(n_2311),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_2393),
.B(n_2311),
.Y(n_2406)
);

NOR4xp25_ASAP7_75t_L g2407 ( 
.A(n_2389),
.B(n_2287),
.C(n_2294),
.D(n_45),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2396),
.B(n_2217),
.Y(n_2408)
);

OAI21xp33_ASAP7_75t_L g2409 ( 
.A1(n_2391),
.A2(n_2298),
.B(n_2254),
.Y(n_2409)
);

OAI32xp33_ASAP7_75t_L g2410 ( 
.A1(n_2401),
.A2(n_2237),
.A3(n_2296),
.B1(n_2021),
.B2(n_2013),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2398),
.Y(n_2411)
);

AOI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2397),
.A2(n_2295),
.B1(n_2170),
.B2(n_2192),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2400),
.B(n_2265),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2402),
.B(n_2275),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_SL g2415 ( 
.A(n_2395),
.B(n_2184),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2390),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2398),
.B(n_2275),
.Y(n_2417)
);

AND2x2_ASAP7_75t_SL g2418 ( 
.A(n_2398),
.B(n_2184),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2393),
.B(n_2267),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2399),
.Y(n_2420)
);

AOI21xp33_ASAP7_75t_SL g2421 ( 
.A1(n_2401),
.A2(n_45),
.B(n_43),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2398),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2398),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2399),
.Y(n_2424)
);

INVxp67_ASAP7_75t_L g2425 ( 
.A(n_2411),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2422),
.B(n_2184),
.Y(n_2426)
);

NAND3xp33_ASAP7_75t_L g2427 ( 
.A(n_2421),
.B(n_2192),
.C(n_42),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2406),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2421),
.B(n_46),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2423),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2413),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2418),
.B(n_2269),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2407),
.B(n_46),
.Y(n_2433)
);

AOI321xp33_ASAP7_75t_SL g2434 ( 
.A1(n_2405),
.A2(n_48),
.A3(n_50),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_2434)
);

O2A1O1Ixp33_ASAP7_75t_L g2435 ( 
.A1(n_2415),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2414),
.Y(n_2436)
);

OAI33xp33_ASAP7_75t_L g2437 ( 
.A1(n_2416),
.A2(n_51),
.A3(n_53),
.B1(n_47),
.B2(n_50),
.B3(n_52),
.Y(n_2437)
);

XNOR2xp5_ASAP7_75t_L g2438 ( 
.A(n_2408),
.B(n_50),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2404),
.B(n_51),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2419),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2417),
.B(n_2275),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2403),
.Y(n_2442)
);

AOI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2409),
.A2(n_2192),
.B1(n_2264),
.B2(n_2255),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2420),
.B(n_51),
.Y(n_2444)
);

INVx1_ASAP7_75t_SL g2445 ( 
.A(n_2424),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2412),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2410),
.B(n_2280),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2422),
.B(n_2280),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2407),
.B(n_2233),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2408),
.A2(n_52),
.B(n_54),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2421),
.B(n_52),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2411),
.Y(n_2452)
);

AOI32xp33_ASAP7_75t_L g2453 ( 
.A1(n_2416),
.A2(n_2264),
.A3(n_2220),
.B1(n_2288),
.B2(n_2162),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2422),
.B(n_2280),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_SL g2455 ( 
.A1(n_2405),
.A2(n_2245),
.B1(n_2284),
.B2(n_2258),
.C(n_2268),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2423),
.B(n_55),
.Y(n_2456)
);

AOI221xp5_ASAP7_75t_L g2457 ( 
.A1(n_2407),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.C(n_58),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2411),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2411),
.Y(n_2459)
);

OAI211xp5_ASAP7_75t_L g2460 ( 
.A1(n_2405),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_2460)
);

AND4x1_ASAP7_75t_L g2461 ( 
.A(n_2411),
.B(n_59),
.C(n_57),
.D(n_58),
.Y(n_2461)
);

AOI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2452),
.A2(n_2264),
.B1(n_2255),
.B2(n_2220),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2461),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2429),
.A2(n_59),
.B(n_60),
.Y(n_2464)
);

OAI21xp33_ASAP7_75t_L g2465 ( 
.A1(n_2458),
.A2(n_2264),
.B(n_2202),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2459),
.A2(n_1986),
.B1(n_1979),
.B2(n_2034),
.Y(n_2466)
);

OAI221xp5_ASAP7_75t_SL g2467 ( 
.A1(n_2457),
.A2(n_2284),
.B1(n_62),
.B2(n_60),
.C(n_61),
.Y(n_2467)
);

OAI222xp33_ASAP7_75t_L g2468 ( 
.A1(n_2445),
.A2(n_2268),
.B1(n_2282),
.B2(n_2270),
.C1(n_62),
.C2(n_64),
.Y(n_2468)
);

OAI222xp33_ASAP7_75t_L g2469 ( 
.A1(n_2425),
.A2(n_2433),
.B1(n_2430),
.B2(n_2442),
.C1(n_2449),
.C2(n_2439),
.Y(n_2469)
);

OAI211xp5_ASAP7_75t_SL g2470 ( 
.A1(n_2436),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_2470)
);

AOI222xp33_ASAP7_75t_L g2471 ( 
.A1(n_2427),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.C1(n_108),
.C2(n_107),
.Y(n_2471)
);

AOI211xp5_ASAP7_75t_SL g2472 ( 
.A1(n_2456),
.A2(n_63),
.B(n_108),
.C(n_107),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2443),
.A2(n_2431),
.B1(n_2438),
.B2(n_2446),
.Y(n_2473)
);

O2A1O1Ixp33_ASAP7_75t_L g2474 ( 
.A1(n_2451),
.A2(n_2460),
.B(n_2435),
.C(n_2444),
.Y(n_2474)
);

AOI22xp33_ASAP7_75t_L g2475 ( 
.A1(n_2437),
.A2(n_1986),
.B1(n_1979),
.B2(n_2034),
.Y(n_2475)
);

INVx2_ASAP7_75t_SL g2476 ( 
.A(n_2461),
.Y(n_2476)
);

AOI321xp33_ASAP7_75t_L g2477 ( 
.A1(n_2450),
.A2(n_2440),
.A3(n_2428),
.B1(n_2426),
.B2(n_2454),
.C(n_2448),
.Y(n_2477)
);

AOI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2426),
.A2(n_2432),
.B1(n_2447),
.B2(n_2453),
.C(n_2441),
.Y(n_2478)
);

OAI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2455),
.A2(n_1986),
.B1(n_1979),
.B2(n_2282),
.Y(n_2479)
);

AOI221xp5_ASAP7_75t_L g2480 ( 
.A1(n_2434),
.A2(n_112),
.B1(n_109),
.B2(n_110),
.C(n_113),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2425),
.A2(n_2200),
.B1(n_2198),
.B2(n_1902),
.Y(n_2481)
);

AOI322xp5_ASAP7_75t_L g2482 ( 
.A1(n_2452),
.A2(n_2261),
.A3(n_2200),
.B1(n_2262),
.B2(n_2221),
.C1(n_2257),
.C2(n_1902),
.Y(n_2482)
);

OAI21xp33_ASAP7_75t_L g2483 ( 
.A1(n_2452),
.A2(n_1902),
.B(n_1899),
.Y(n_2483)
);

AOI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2452),
.A2(n_2034),
.B1(n_1938),
.B2(n_1946),
.Y(n_2484)
);

AOI21xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2427),
.A2(n_113),
.B(n_114),
.Y(n_2485)
);

OAI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2457),
.A2(n_2040),
.B1(n_116),
.B2(n_114),
.C(n_115),
.Y(n_2486)
);

OAI221xp5_ASAP7_75t_L g2487 ( 
.A1(n_2457),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_2487)
);

O2A1O1Ixp33_ASAP7_75t_L g2488 ( 
.A1(n_2433),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2461),
.Y(n_2489)
);

OAI22x1_ASAP7_75t_L g2490 ( 
.A1(n_2461),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2461),
.Y(n_2491)
);

AOI221xp5_ASAP7_75t_SL g2492 ( 
.A1(n_2425),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_2492)
);

OAI211xp5_ASAP7_75t_SL g2493 ( 
.A1(n_2425),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_2493)
);

OAI222xp33_ASAP7_75t_L g2494 ( 
.A1(n_2445),
.A2(n_150),
.B1(n_133),
.B2(n_159),
.C1(n_141),
.C2(n_125),
.Y(n_2494)
);

AOI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2429),
.A2(n_125),
.B(n_126),
.Y(n_2495)
);

OAI222xp33_ASAP7_75t_L g2496 ( 
.A1(n_2445),
.A2(n_153),
.B1(n_134),
.B2(n_161),
.C1(n_142),
.C2(n_126),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2461),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2461),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2461),
.Y(n_2499)
);

NOR3xp33_ASAP7_75t_L g2500 ( 
.A(n_2469),
.B(n_129),
.C(n_128),
.Y(n_2500)
);

NOR4xp25_ASAP7_75t_SL g2501 ( 
.A(n_2463),
.B(n_129),
.C(n_127),
.D(n_128),
.Y(n_2501)
);

OAI222xp33_ASAP7_75t_L g2502 ( 
.A1(n_2476),
.A2(n_131),
.B1(n_133),
.B2(n_127),
.C1(n_130),
.C2(n_132),
.Y(n_2502)
);

OAI221xp5_ASAP7_75t_SL g2503 ( 
.A1(n_2480),
.A2(n_134),
.B1(n_130),
.B2(n_132),
.C(n_135),
.Y(n_2503)
);

AOI211xp5_ASAP7_75t_L g2504 ( 
.A1(n_2467),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2489),
.B(n_136),
.Y(n_2505)
);

AOI221xp5_ASAP7_75t_L g2506 ( 
.A1(n_2485),
.A2(n_2473),
.B1(n_2486),
.B2(n_2497),
.C(n_2491),
.Y(n_2506)
);

AOI222xp33_ASAP7_75t_L g2507 ( 
.A1(n_2498),
.A2(n_141),
.B1(n_143),
.B2(n_139),
.C1(n_140),
.C2(n_142),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2464),
.A2(n_151),
.B(n_139),
.Y(n_2508)
);

NAND4xp25_ASAP7_75t_SL g2509 ( 
.A(n_2471),
.B(n_144),
.C(n_140),
.D(n_143),
.Y(n_2509)
);

AOI21xp33_ASAP7_75t_L g2510 ( 
.A1(n_2488),
.A2(n_144),
.B(n_146),
.Y(n_2510)
);

AOI211xp5_ASAP7_75t_L g2511 ( 
.A1(n_2487),
.A2(n_2470),
.B(n_2499),
.C(n_2474),
.Y(n_2511)
);

OAI211xp5_ASAP7_75t_L g2512 ( 
.A1(n_2478),
.A2(n_2477),
.B(n_2495),
.C(n_2492),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_SL g2513 ( 
.A(n_2493),
.B(n_147),
.C(n_148),
.Y(n_2513)
);

AOI221xp5_ASAP7_75t_L g2514 ( 
.A1(n_2468),
.A2(n_151),
.B1(n_155),
.B2(n_149),
.C(n_154),
.Y(n_2514)
);

OAI211xp5_ASAP7_75t_L g2515 ( 
.A1(n_2472),
.A2(n_154),
.B(n_148),
.C(n_149),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2490),
.Y(n_2516)
);

AOI211xp5_ASAP7_75t_L g2517 ( 
.A1(n_2483),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2475),
.B(n_157),
.C(n_158),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2462),
.A2(n_1938),
.B1(n_1946),
.B2(n_1935),
.Y(n_2519)
);

HB1xp67_ASAP7_75t_L g2520 ( 
.A(n_2494),
.Y(n_2520)
);

OAI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2481),
.A2(n_177),
.B1(n_185),
.B2(n_168),
.C(n_159),
.Y(n_2521)
);

OAI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2484),
.A2(n_1938),
.B1(n_1946),
.B2(n_1935),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2466),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2496),
.A2(n_169),
.B(n_160),
.Y(n_2524)
);

NAND2x1_ASAP7_75t_L g2525 ( 
.A(n_2479),
.B(n_2201),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2465),
.A2(n_1935),
.B1(n_2198),
.B2(n_2277),
.Y(n_2526)
);

AOI221xp5_ASAP7_75t_L g2527 ( 
.A1(n_2482),
.A2(n_163),
.B1(n_165),
.B2(n_162),
.C(n_164),
.Y(n_2527)
);

NAND4xp25_ASAP7_75t_L g2528 ( 
.A(n_2480),
.B(n_169),
.C(n_178),
.D(n_160),
.Y(n_2528)
);

AOI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_2485),
.A2(n_164),
.B1(n_166),
.B2(n_163),
.C(n_165),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2476),
.B(n_162),
.Y(n_2530)
);

OAI21xp5_ASAP7_75t_SL g2531 ( 
.A1(n_2469),
.A2(n_167),
.B(n_168),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2469),
.A2(n_170),
.B(n_172),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2490),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2490),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2476),
.B(n_170),
.Y(n_2535)
);

NAND3xp33_ASAP7_75t_SL g2536 ( 
.A(n_2471),
.B(n_173),
.C(n_174),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2476),
.A2(n_174),
.B(n_175),
.Y(n_2537)
);

XNOR2x1_ASAP7_75t_L g2538 ( 
.A(n_2490),
.B(n_175),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2490),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_SL g2540 ( 
.A(n_2471),
.B(n_176),
.C(n_177),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2476),
.B(n_176),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2476),
.A2(n_2198),
.B1(n_2216),
.B2(n_2281),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2476),
.B(n_178),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2476),
.B(n_179),
.Y(n_2544)
);

AOI322xp5_ASAP7_75t_L g2545 ( 
.A1(n_2480),
.A2(n_2261),
.A3(n_184),
.B1(n_181),
.B2(n_183),
.C1(n_179),
.C2(n_180),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2476),
.B(n_180),
.Y(n_2546)
);

AOI221xp5_ASAP7_75t_L g2547 ( 
.A1(n_2485),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2476),
.B(n_2280),
.Y(n_2548)
);

OAI21xp33_ASAP7_75t_SL g2549 ( 
.A1(n_2476),
.A2(n_2277),
.B(n_2281),
.Y(n_2549)
);

AOI221xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2480),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_2550)
);

OAI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2480),
.A2(n_2283),
.B(n_2193),
.Y(n_2551)
);

OAI211xp5_ASAP7_75t_L g2552 ( 
.A1(n_2471),
.A2(n_189),
.B(n_186),
.C(n_187),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_SL g2553 ( 
.A1(n_2490),
.A2(n_189),
.B(n_191),
.Y(n_2553)
);

AOI221x1_ASAP7_75t_SL g2554 ( 
.A1(n_2473),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_2554)
);

OAI211xp5_ASAP7_75t_SL g2555 ( 
.A1(n_2478),
.A2(n_195),
.B(n_192),
.C(n_193),
.Y(n_2555)
);

OAI221xp5_ASAP7_75t_L g2556 ( 
.A1(n_2476),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_2556)
);

AOI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2485),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_2557)
);

AOI21xp33_ASAP7_75t_SL g2558 ( 
.A1(n_2490),
.A2(n_200),
.B(n_201),
.Y(n_2558)
);

AOI211xp5_ASAP7_75t_L g2559 ( 
.A1(n_2467),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_2559)
);

NAND4xp25_ASAP7_75t_L g2560 ( 
.A(n_2480),
.B(n_205),
.C(n_203),
.D(n_204),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2476),
.A2(n_203),
.B(n_204),
.Y(n_2561)
);

AOI211xp5_ASAP7_75t_L g2562 ( 
.A1(n_2467),
.A2(n_208),
.B(n_205),
.C(n_206),
.Y(n_2562)
);

AOI221xp5_ASAP7_75t_L g2563 ( 
.A1(n_2485),
.A2(n_210),
.B1(n_206),
.B2(n_209),
.C(n_211),
.Y(n_2563)
);

OAI221xp5_ASAP7_75t_SL g2564 ( 
.A1(n_2531),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_2564)
);

AOI31xp33_ASAP7_75t_L g2565 ( 
.A1(n_2538),
.A2(n_214),
.A3(n_212),
.B(n_213),
.Y(n_2565)
);

OAI221xp5_ASAP7_75t_SL g2566 ( 
.A1(n_2532),
.A2(n_217),
.B1(n_213),
.B2(n_215),
.C(n_218),
.Y(n_2566)
);

AOI222xp33_ASAP7_75t_L g2567 ( 
.A1(n_2518),
.A2(n_220),
.B1(n_222),
.B2(n_217),
.C1(n_219),
.C2(n_221),
.Y(n_2567)
);

NAND4xp75_ASAP7_75t_L g2568 ( 
.A(n_2506),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2568)
);

AOI211xp5_ASAP7_75t_L g2569 ( 
.A1(n_2503),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2554),
.B(n_223),
.Y(n_2570)
);

OAI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2514),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.C(n_228),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2516),
.A2(n_2276),
.B1(n_2208),
.B2(n_227),
.Y(n_2572)
);

AOI21xp33_ASAP7_75t_L g2573 ( 
.A1(n_2505),
.A2(n_225),
.B(n_226),
.Y(n_2573)
);

OAI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2550),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_2574)
);

OAI211xp5_ASAP7_75t_L g2575 ( 
.A1(n_2553),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2508),
.A2(n_232),
.B(n_233),
.Y(n_2576)
);

NOR4xp25_ASAP7_75t_SL g2577 ( 
.A(n_2558),
.B(n_234),
.C(n_232),
.D(n_233),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2528),
.B(n_234),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2530),
.A2(n_235),
.B(n_236),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2535),
.Y(n_2580)
);

AOI22xp5_ASAP7_75t_L g2581 ( 
.A1(n_2500),
.A2(n_2276),
.B1(n_2283),
.B2(n_2274),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2541),
.Y(n_2582)
);

A2O1A1Ixp33_ASAP7_75t_L g2583 ( 
.A1(n_2537),
.A2(n_238),
.B(n_235),
.C(n_237),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2544),
.B(n_237),
.Y(n_2584)
);

AOI221xp5_ASAP7_75t_L g2585 ( 
.A1(n_2510),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2529),
.B(n_239),
.Y(n_2586)
);

OAI32xp33_ASAP7_75t_L g2587 ( 
.A1(n_2543),
.A2(n_242),
.A3(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_2587)
);

OAI221xp5_ASAP7_75t_SL g2588 ( 
.A1(n_2545),
.A2(n_245),
.B1(n_242),
.B2(n_244),
.C(n_246),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2524),
.A2(n_244),
.B(n_245),
.Y(n_2589)
);

AOI211xp5_ASAP7_75t_L g2590 ( 
.A1(n_2515),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_2590)
);

NOR3xp33_ASAP7_75t_L g2591 ( 
.A(n_2512),
.B(n_247),
.C(n_248),
.Y(n_2591)
);

NOR3xp33_ASAP7_75t_L g2592 ( 
.A(n_2511),
.B(n_249),
.C(n_250),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2533),
.B(n_2280),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2546),
.A2(n_249),
.B(n_250),
.Y(n_2594)
);

AOI221xp5_ASAP7_75t_L g2595 ( 
.A1(n_2555),
.A2(n_2509),
.B1(n_2560),
.B2(n_2527),
.C(n_2539),
.Y(n_2595)
);

NAND3xp33_ASAP7_75t_SL g2596 ( 
.A(n_2501),
.B(n_251),
.C(n_252),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2534),
.B(n_251),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_SL g2598 ( 
.A(n_2502),
.B(n_252),
.Y(n_2598)
);

AOI21xp33_ASAP7_75t_L g2599 ( 
.A1(n_2552),
.A2(n_253),
.B(n_254),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2561),
.B(n_253),
.Y(n_2600)
);

NOR3xp33_ASAP7_75t_L g2601 ( 
.A(n_2536),
.B(n_2540),
.C(n_2547),
.Y(n_2601)
);

OAI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2504),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_2602)
);

NOR4xp25_ASAP7_75t_L g2603 ( 
.A(n_2523),
.B(n_257),
.C(n_255),
.D(n_256),
.Y(n_2603)
);

AOI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2520),
.A2(n_2276),
.B1(n_2274),
.B2(n_261),
.Y(n_2604)
);

OAI221xp5_ASAP7_75t_SL g2605 ( 
.A1(n_2559),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.C(n_264),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2513),
.Y(n_2606)
);

AOI211xp5_ASAP7_75t_L g2607 ( 
.A1(n_2521),
.A2(n_2557),
.B(n_2563),
.C(n_2562),
.Y(n_2607)
);

OAI21xp33_ASAP7_75t_SL g2608 ( 
.A1(n_2526),
.A2(n_260),
.B(n_262),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2548),
.A2(n_2276),
.B1(n_266),
.B2(n_264),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2525),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2551),
.B(n_2519),
.Y(n_2611)
);

AOI211xp5_ASAP7_75t_L g2612 ( 
.A1(n_2556),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2612)
);

AOI221xp5_ASAP7_75t_L g2613 ( 
.A1(n_2522),
.A2(n_268),
.B1(n_265),
.B2(n_267),
.C(n_269),
.Y(n_2613)
);

AOI211xp5_ASAP7_75t_SL g2614 ( 
.A1(n_2517),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2549),
.B(n_270),
.Y(n_2615)
);

NOR3xp33_ASAP7_75t_L g2616 ( 
.A(n_2507),
.B(n_271),
.C(n_272),
.Y(n_2616)
);

NOR3xp33_ASAP7_75t_L g2617 ( 
.A(n_2507),
.B(n_272),
.C(n_273),
.Y(n_2617)
);

AOI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2542),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2618)
);

AOI322xp5_ASAP7_75t_L g2619 ( 
.A1(n_2516),
.A2(n_281),
.A3(n_280),
.B1(n_277),
.B2(n_275),
.C1(n_276),
.C2(n_279),
.Y(n_2619)
);

AOI211xp5_ASAP7_75t_L g2620 ( 
.A1(n_2503),
.A2(n_281),
.B(n_276),
.C(n_279),
.Y(n_2620)
);

AOI221x1_ASAP7_75t_L g2621 ( 
.A1(n_2500),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2621)
);

OAI211xp5_ASAP7_75t_SL g2622 ( 
.A1(n_2506),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_SL g2623 ( 
.A1(n_2531),
.A2(n_286),
.B(n_287),
.Y(n_2623)
);

AOI221x1_ASAP7_75t_L g2624 ( 
.A1(n_2500),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.C(n_289),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_SL g2625 ( 
.A1(n_2520),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2553),
.A2(n_291),
.B(n_292),
.Y(n_2626)
);

AOI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2500),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2528),
.B(n_294),
.Y(n_2628)
);

OAI211xp5_ASAP7_75t_L g2629 ( 
.A1(n_2531),
.A2(n_297),
.B(n_295),
.C(n_296),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2558),
.B(n_295),
.Y(n_2630)
);

AOI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2500),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_2631)
);

AO21x2_ASAP7_75t_L g2632 ( 
.A1(n_2530),
.A2(n_298),
.B(n_299),
.Y(n_2632)
);

AOI221xp5_ASAP7_75t_L g2633 ( 
.A1(n_2558),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.C(n_303),
.Y(n_2633)
);

OAI321xp33_ASAP7_75t_L g2634 ( 
.A1(n_2555),
.A2(n_302),
.A3(n_305),
.B1(n_300),
.B2(n_301),
.C(n_304),
.Y(n_2634)
);

OAI22xp33_ASAP7_75t_SL g2635 ( 
.A1(n_2530),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_2635)
);

OAI221xp5_ASAP7_75t_L g2636 ( 
.A1(n_2554),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.C(n_309),
.Y(n_2636)
);

AOI22xp33_ASAP7_75t_SL g2637 ( 
.A1(n_2520),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_2637)
);

AOI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2558),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.C(n_313),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2535),
.Y(n_2639)
);

NAND4xp25_ASAP7_75t_SL g2640 ( 
.A(n_2550),
.B(n_314),
.C(n_312),
.D(n_313),
.Y(n_2640)
);

NAND3xp33_ASAP7_75t_L g2641 ( 
.A(n_2591),
.B(n_314),
.C(n_315),
.Y(n_2641)
);

OAI21xp33_ASAP7_75t_L g2642 ( 
.A1(n_2598),
.A2(n_315),
.B(n_316),
.Y(n_2642)
);

NAND3xp33_ASAP7_75t_L g2643 ( 
.A(n_2592),
.B(n_2585),
.C(n_2633),
.Y(n_2643)
);

NAND3xp33_ASAP7_75t_L g2644 ( 
.A(n_2638),
.B(n_317),
.C(n_318),
.Y(n_2644)
);

O2A1O1Ixp5_ASAP7_75t_L g2645 ( 
.A1(n_2630),
.A2(n_319),
.B(n_317),
.C(n_318),
.Y(n_2645)
);

NOR4xp25_ASAP7_75t_L g2646 ( 
.A(n_2596),
.B(n_322),
.C(n_320),
.D(n_321),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_2565),
.B(n_320),
.Y(n_2647)
);

NOR3xp33_ASAP7_75t_L g2648 ( 
.A(n_2606),
.B(n_321),
.C(n_323),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2597),
.B(n_323),
.Y(n_2649)
);

OAI211xp5_ASAP7_75t_L g2650 ( 
.A1(n_2627),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_2650)
);

NAND3xp33_ASAP7_75t_SL g2651 ( 
.A(n_2577),
.B(n_327),
.C(n_328),
.Y(n_2651)
);

XNOR2xp5_ASAP7_75t_L g2652 ( 
.A(n_2568),
.B(n_327),
.Y(n_2652)
);

NOR2x1_ASAP7_75t_L g2653 ( 
.A(n_2632),
.B(n_328),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2634),
.B(n_329),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2564),
.B(n_329),
.Y(n_2655)
);

NAND3xp33_ASAP7_75t_L g2656 ( 
.A(n_2590),
.B(n_331),
.C(n_332),
.Y(n_2656)
);

NAND3xp33_ASAP7_75t_SL g2657 ( 
.A(n_2626),
.B(n_331),
.C(n_332),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2570),
.Y(n_2658)
);

NAND4xp25_ASAP7_75t_L g2659 ( 
.A(n_2628),
.B(n_335),
.C(n_333),
.D(n_334),
.Y(n_2659)
);

NOR3xp33_ASAP7_75t_L g2660 ( 
.A(n_2584),
.B(n_333),
.C(n_334),
.Y(n_2660)
);

OAI32xp33_ASAP7_75t_L g2661 ( 
.A1(n_2616),
.A2(n_2617),
.A3(n_2608),
.B1(n_2578),
.B2(n_2600),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2603),
.B(n_335),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2631),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_2663)
);

AOI31xp33_ASAP7_75t_L g2664 ( 
.A1(n_2569),
.A2(n_339),
.A3(n_337),
.B(n_338),
.Y(n_2664)
);

NAND4xp75_ASAP7_75t_L g2665 ( 
.A(n_2621),
.B(n_342),
.C(n_340),
.D(n_341),
.Y(n_2665)
);

OAI21xp5_ASAP7_75t_SL g2666 ( 
.A1(n_2623),
.A2(n_340),
.B(n_341),
.Y(n_2666)
);

NOR2x1_ASAP7_75t_L g2667 ( 
.A(n_2632),
.B(n_342),
.Y(n_2667)
);

NAND3x1_ASAP7_75t_L g2668 ( 
.A(n_2601),
.B(n_2589),
.C(n_2580),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2636),
.B(n_343),
.Y(n_2669)
);

OAI221xp5_ASAP7_75t_L g2670 ( 
.A1(n_2618),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_2670)
);

NAND3xp33_ASAP7_75t_L g2671 ( 
.A(n_2567),
.B(n_345),
.C(n_346),
.Y(n_2671)
);

AOI221xp5_ASAP7_75t_L g2672 ( 
.A1(n_2599),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.C(n_350),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2575),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2576),
.A2(n_348),
.B(n_350),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2586),
.A2(n_351),
.B(n_352),
.Y(n_2675)
);

O2A1O1Ixp33_ASAP7_75t_L g2676 ( 
.A1(n_2583),
.A2(n_354),
.B(n_351),
.C(n_353),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2615),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2629),
.Y(n_2678)
);

NAND4xp25_ASAP7_75t_L g2679 ( 
.A(n_2595),
.B(n_358),
.C(n_355),
.D(n_356),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2574),
.B(n_355),
.Y(n_2680)
);

NAND4xp75_ASAP7_75t_L g2681 ( 
.A(n_2624),
.B(n_359),
.C(n_356),
.D(n_358),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2614),
.B(n_2225),
.Y(n_2682)
);

AOI22xp5_ASAP7_75t_L g2683 ( 
.A1(n_2640),
.A2(n_2622),
.B1(n_2639),
.B2(n_2593),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2635),
.Y(n_2684)
);

NOR3x1_ASAP7_75t_L g2685 ( 
.A(n_2602),
.B(n_2571),
.C(n_2611),
.Y(n_2685)
);

OR3x1_ASAP7_75t_L g2686 ( 
.A(n_2587),
.B(n_359),
.C(n_360),
.Y(n_2686)
);

AOI211xp5_ASAP7_75t_L g2687 ( 
.A1(n_2588),
.A2(n_2605),
.B(n_2566),
.C(n_2594),
.Y(n_2687)
);

INVx2_ASAP7_75t_SL g2688 ( 
.A(n_2610),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2620),
.Y(n_2689)
);

NAND3xp33_ASAP7_75t_SL g2690 ( 
.A(n_2612),
.B(n_360),
.C(n_361),
.Y(n_2690)
);

NOR4xp25_ASAP7_75t_L g2691 ( 
.A(n_2582),
.B(n_363),
.C(n_361),
.D(n_362),
.Y(n_2691)
);

OAI221xp5_ASAP7_75t_L g2692 ( 
.A1(n_2609),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.C(n_365),
.Y(n_2692)
);

AOI211xp5_ASAP7_75t_L g2693 ( 
.A1(n_2613),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_2693)
);

NOR2x1_ASAP7_75t_L g2694 ( 
.A(n_2579),
.B(n_367),
.Y(n_2694)
);

NOR3xp33_ASAP7_75t_L g2695 ( 
.A(n_2573),
.B(n_368),
.C(n_369),
.Y(n_2695)
);

OAI21xp33_ASAP7_75t_L g2696 ( 
.A1(n_2604),
.A2(n_2607),
.B(n_2625),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2637),
.A2(n_2572),
.B(n_2581),
.Y(n_2697)
);

NOR2x1_ASAP7_75t_L g2698 ( 
.A(n_2619),
.B(n_368),
.Y(n_2698)
);

NAND4xp25_ASAP7_75t_L g2699 ( 
.A(n_2595),
.B(n_371),
.C(n_369),
.D(n_370),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_SL g2700 ( 
.A(n_2577),
.B(n_370),
.C(n_372),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2597),
.B(n_372),
.Y(n_2701)
);

NOR3x1_ASAP7_75t_L g2702 ( 
.A(n_2568),
.B(n_373),
.C(n_374),
.Y(n_2702)
);

NAND5xp2_ASAP7_75t_L g2703 ( 
.A(n_2595),
.B(n_377),
.C(n_374),
.D(n_376),
.E(n_378),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2597),
.B(n_377),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_SL g2705 ( 
.A(n_2568),
.B(n_378),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2634),
.B(n_379),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2630),
.A2(n_380),
.B(n_381),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2634),
.B(n_381),
.Y(n_2708)
);

NAND3xp33_ASAP7_75t_L g2709 ( 
.A(n_2591),
.B(n_382),
.C(n_383),
.Y(n_2709)
);

AND4x1_ASAP7_75t_L g2710 ( 
.A(n_2646),
.B(n_384),
.C(n_382),
.D(n_383),
.Y(n_2710)
);

OAI211xp5_ASAP7_75t_SL g2711 ( 
.A1(n_2642),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_2711)
);

OAI211xp5_ASAP7_75t_SL g2712 ( 
.A1(n_2696),
.A2(n_389),
.B(n_386),
.C(n_387),
.Y(n_2712)
);

NOR3xp33_ASAP7_75t_L g2713 ( 
.A(n_2688),
.B(n_389),
.C(n_390),
.Y(n_2713)
);

NAND4xp25_ASAP7_75t_SL g2714 ( 
.A(n_2672),
.B(n_392),
.C(n_390),
.D(n_391),
.Y(n_2714)
);

NAND4xp25_ASAP7_75t_L g2715 ( 
.A(n_2687),
.B(n_393),
.C(n_391),
.D(n_392),
.Y(n_2715)
);

AOI222xp33_ASAP7_75t_L g2716 ( 
.A1(n_2651),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.C1(n_397),
.C2(n_398),
.Y(n_2716)
);

OAI211xp5_ASAP7_75t_SL g2717 ( 
.A1(n_2683),
.A2(n_397),
.B(n_394),
.C(n_395),
.Y(n_2717)
);

NAND3xp33_ASAP7_75t_SL g2718 ( 
.A(n_2705),
.B(n_398),
.C(n_399),
.Y(n_2718)
);

AOI221xp5_ASAP7_75t_L g2719 ( 
.A1(n_2664),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.C(n_402),
.Y(n_2719)
);

XNOR2x1_ASAP7_75t_L g2720 ( 
.A(n_2653),
.B(n_400),
.Y(n_2720)
);

OAI221xp5_ASAP7_75t_L g2721 ( 
.A1(n_2666),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.C(n_405),
.Y(n_2721)
);

AOI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2655),
.A2(n_406),
.B1(n_403),
.B2(n_404),
.Y(n_2722)
);

OAI211xp5_ASAP7_75t_SL g2723 ( 
.A1(n_2698),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2723)
);

NOR4xp25_ASAP7_75t_L g2724 ( 
.A(n_2668),
.B(n_410),
.C(n_408),
.D(n_409),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2703),
.B(n_2659),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2667),
.B(n_409),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2700),
.B(n_410),
.Y(n_2727)
);

NOR3xp33_ASAP7_75t_L g2728 ( 
.A(n_2673),
.B(n_411),
.C(n_412),
.Y(n_2728)
);

NOR4xp25_ASAP7_75t_L g2729 ( 
.A(n_2690),
.B(n_414),
.C(n_411),
.D(n_413),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2647),
.B(n_2225),
.Y(n_2730)
);

NAND4xp25_ASAP7_75t_L g2731 ( 
.A(n_2685),
.B(n_415),
.C(n_413),
.D(n_414),
.Y(n_2731)
);

NOR3xp33_ASAP7_75t_L g2732 ( 
.A(n_2684),
.B(n_415),
.C(n_416),
.Y(n_2732)
);

AND4x1_ASAP7_75t_L g2733 ( 
.A(n_2702),
.B(n_418),
.C(n_416),
.D(n_417),
.Y(n_2733)
);

AOI221x1_ASAP7_75t_L g2734 ( 
.A1(n_2677),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.C(n_421),
.Y(n_2734)
);

NOR3xp33_ASAP7_75t_SL g2735 ( 
.A(n_2657),
.B(n_420),
.C(n_421),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2694),
.B(n_422),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2669),
.B(n_2691),
.Y(n_2737)
);

INVx1_ASAP7_75t_SL g2738 ( 
.A(n_2686),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2665),
.Y(n_2739)
);

NAND3xp33_ASAP7_75t_SL g2740 ( 
.A(n_2695),
.B(n_422),
.C(n_423),
.Y(n_2740)
);

INVxp33_ASAP7_75t_L g2741 ( 
.A(n_2679),
.Y(n_2741)
);

OAI221xp5_ASAP7_75t_L g2742 ( 
.A1(n_2692),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.C(n_427),
.Y(n_2742)
);

NOR3xp33_ASAP7_75t_L g2743 ( 
.A(n_2678),
.B(n_424),
.C(n_425),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2648),
.B(n_426),
.Y(n_2744)
);

NOR2x1_ASAP7_75t_SL g2745 ( 
.A(n_2681),
.B(n_427),
.Y(n_2745)
);

NAND3xp33_ASAP7_75t_L g2746 ( 
.A(n_2660),
.B(n_428),
.C(n_429),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2676),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_2747)
);

INVxp67_ASAP7_75t_L g2748 ( 
.A(n_2680),
.Y(n_2748)
);

AND4x1_ASAP7_75t_L g2749 ( 
.A(n_2645),
.B(n_432),
.C(n_430),
.D(n_431),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2659),
.B(n_432),
.Y(n_2750)
);

NAND3xp33_ASAP7_75t_SL g2751 ( 
.A(n_2693),
.B(n_433),
.C(n_434),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2652),
.B(n_2224),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2649),
.Y(n_2753)
);

NOR3xp33_ASAP7_75t_L g2754 ( 
.A(n_2689),
.B(n_433),
.C(n_434),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_SL g2755 ( 
.A(n_2641),
.B(n_435),
.Y(n_2755)
);

NAND4xp25_ASAP7_75t_L g2756 ( 
.A(n_2709),
.B(n_438),
.C(n_436),
.D(n_437),
.Y(n_2756)
);

NAND2x1_ASAP7_75t_SL g2757 ( 
.A(n_2658),
.B(n_436),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2701),
.Y(n_2758)
);

NOR2x1_ASAP7_75t_L g2759 ( 
.A(n_2699),
.B(n_437),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2704),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2682),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2674),
.B(n_438),
.Y(n_2762)
);

NAND4xp25_ASAP7_75t_L g2763 ( 
.A(n_2656),
.B(n_2643),
.C(n_2671),
.D(n_2644),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2707),
.B(n_439),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2757),
.Y(n_2765)
);

NOR2x1_ASAP7_75t_L g2766 ( 
.A(n_2720),
.B(n_2662),
.Y(n_2766)
);

NOR2x1_ASAP7_75t_L g2767 ( 
.A(n_2726),
.B(n_2650),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2725),
.A2(n_2708),
.B1(n_2706),
.B2(n_2654),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2727),
.Y(n_2769)
);

INVx1_ASAP7_75t_SL g2770 ( 
.A(n_2736),
.Y(n_2770)
);

NOR2x1_ASAP7_75t_L g2771 ( 
.A(n_2731),
.B(n_2663),
.Y(n_2771)
);

OAI21xp33_ASAP7_75t_L g2772 ( 
.A1(n_2741),
.A2(n_2675),
.B(n_2661),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2745),
.B(n_2697),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2739),
.B(n_2670),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2710),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2750),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2724),
.B(n_440),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_SL g2778 ( 
.A1(n_2729),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_2778)
);

NOR2x1_ASAP7_75t_L g2779 ( 
.A(n_2736),
.B(n_444),
.Y(n_2779)
);

AO22x2_ASAP7_75t_L g2780 ( 
.A1(n_2738),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2733),
.Y(n_2781)
);

NOR2x1_ASAP7_75t_L g2782 ( 
.A(n_2718),
.B(n_445),
.Y(n_2782)
);

AOI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2714),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2764),
.Y(n_2784)
);

AO22x1_ASAP7_75t_L g2785 ( 
.A1(n_2732),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2717),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2749),
.Y(n_2787)
);

AOI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2723),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2716),
.B(n_455),
.Y(n_2789)
);

NOR2xp33_ASAP7_75t_L g2790 ( 
.A(n_2756),
.B(n_456),
.Y(n_2790)
);

NOR2x1_ASAP7_75t_L g2791 ( 
.A(n_2715),
.B(n_456),
.Y(n_2791)
);

NOR2x1_ASAP7_75t_L g2792 ( 
.A(n_2746),
.B(n_457),
.Y(n_2792)
);

AND3x4_ASAP7_75t_L g2793 ( 
.A(n_2735),
.B(n_457),
.C(n_459),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2713),
.B(n_462),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2712),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2728),
.B(n_2743),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2759),
.Y(n_2797)
);

NOR2x1_ASAP7_75t_L g2798 ( 
.A(n_2763),
.B(n_464),
.Y(n_2798)
);

AO22x2_ASAP7_75t_L g2799 ( 
.A1(n_2761),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_2799)
);

INVx3_ASAP7_75t_L g2800 ( 
.A(n_2764),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2722),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2711),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_2802)
);

BUFx3_ASAP7_75t_L g2803 ( 
.A(n_2737),
.Y(n_2803)
);

NOR2x1_ASAP7_75t_L g2804 ( 
.A(n_2740),
.B(n_468),
.Y(n_2804)
);

NAND3xp33_ASAP7_75t_L g2805 ( 
.A(n_2719),
.B(n_469),
.C(n_470),
.Y(n_2805)
);

NOR2x1_ASAP7_75t_L g2806 ( 
.A(n_2751),
.B(n_471),
.Y(n_2806)
);

NOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2762),
.B(n_471),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2734),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2754),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2744),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2730),
.Y(n_2811)
);

AO22x2_ASAP7_75t_L g2812 ( 
.A1(n_2753),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_2812)
);

HB1xp67_ASAP7_75t_L g2813 ( 
.A(n_2721),
.Y(n_2813)
);

NOR3xp33_ASAP7_75t_L g2814 ( 
.A(n_2772),
.B(n_2748),
.C(n_2758),
.Y(n_2814)
);

NOR4xp25_ASAP7_75t_L g2815 ( 
.A(n_2770),
.B(n_2755),
.C(n_2760),
.D(n_2747),
.Y(n_2815)
);

NOR3xp33_ASAP7_75t_L g2816 ( 
.A(n_2800),
.B(n_2742),
.C(n_2752),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2777),
.B(n_472),
.Y(n_2817)
);

NOR2x1_ASAP7_75t_L g2818 ( 
.A(n_2779),
.B(n_473),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2785),
.B(n_474),
.Y(n_2819)
);

NAND5xp2_ASAP7_75t_L g2820 ( 
.A(n_2768),
.B(n_475),
.C(n_476),
.D(n_477),
.E(n_478),
.Y(n_2820)
);

NOR3xp33_ASAP7_75t_L g2821 ( 
.A(n_2765),
.B(n_475),
.C(n_476),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2783),
.B(n_477),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2778),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2791),
.B(n_2224),
.Y(n_2824)
);

NAND4xp25_ASAP7_75t_L g2825 ( 
.A(n_2790),
.B(n_481),
.C(n_479),
.D(n_480),
.Y(n_2825)
);

NAND3x1_ASAP7_75t_L g2826 ( 
.A(n_2798),
.B(n_479),
.C(n_482),
.Y(n_2826)
);

NAND3xp33_ASAP7_75t_SL g2827 ( 
.A(n_2808),
.B(n_482),
.C(n_483),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2793),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_2828)
);

NAND3xp33_ASAP7_75t_L g2829 ( 
.A(n_2807),
.B(n_484),
.C(n_485),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2780),
.Y(n_2830)
);

NAND3xp33_ASAP7_75t_L g2831 ( 
.A(n_2775),
.B(n_486),
.C(n_487),
.Y(n_2831)
);

NAND3xp33_ASAP7_75t_L g2832 ( 
.A(n_2787),
.B(n_487),
.C(n_489),
.Y(n_2832)
);

NOR4xp25_ASAP7_75t_L g2833 ( 
.A(n_2781),
.B(n_491),
.C(n_489),
.D(n_490),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2794),
.B(n_490),
.Y(n_2834)
);

NOR3x2_ASAP7_75t_L g2835 ( 
.A(n_2799),
.B(n_491),
.C(n_492),
.Y(n_2835)
);

NOR2x1_ASAP7_75t_L g2836 ( 
.A(n_2766),
.B(n_492),
.Y(n_2836)
);

NOR3xp33_ASAP7_75t_L g2837 ( 
.A(n_2797),
.B(n_2773),
.C(n_2769),
.Y(n_2837)
);

NOR3xp33_ASAP7_75t_SL g2838 ( 
.A(n_2789),
.B(n_493),
.C(n_494),
.Y(n_2838)
);

NAND3xp33_ASAP7_75t_L g2839 ( 
.A(n_2803),
.B(n_493),
.C(n_494),
.Y(n_2839)
);

NAND4xp75_ASAP7_75t_L g2840 ( 
.A(n_2767),
.B(n_495),
.C(n_496),
.D(n_497),
.Y(n_2840)
);

NAND4xp25_ASAP7_75t_SL g2841 ( 
.A(n_2802),
.B(n_495),
.C(n_496),
.D(n_498),
.Y(n_2841)
);

NOR2x1_ASAP7_75t_L g2842 ( 
.A(n_2784),
.B(n_498),
.Y(n_2842)
);

AND3x2_ASAP7_75t_L g2843 ( 
.A(n_2809),
.B(n_499),
.C(n_500),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2788),
.B(n_500),
.Y(n_2844)
);

INVx1_ASAP7_75t_SL g2845 ( 
.A(n_2835),
.Y(n_2845)
);

NOR3xp33_ASAP7_75t_L g2846 ( 
.A(n_2837),
.B(n_2823),
.C(n_2814),
.Y(n_2846)
);

NAND4xp25_ASAP7_75t_SL g2847 ( 
.A(n_2828),
.B(n_2786),
.C(n_2795),
.D(n_2805),
.Y(n_2847)
);

NAND4xp25_ASAP7_75t_L g2848 ( 
.A(n_2816),
.B(n_2771),
.C(n_2806),
.D(n_2782),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2843),
.Y(n_2849)
);

NAND3x1_ASAP7_75t_L g2850 ( 
.A(n_2818),
.B(n_2804),
.C(n_2792),
.Y(n_2850)
);

AOI221xp5_ASAP7_75t_L g2851 ( 
.A1(n_2815),
.A2(n_2774),
.B1(n_2801),
.B2(n_2813),
.C(n_2811),
.Y(n_2851)
);

HB1xp67_ASAP7_75t_L g2852 ( 
.A(n_2842),
.Y(n_2852)
);

AO22x1_ASAP7_75t_L g2853 ( 
.A1(n_2836),
.A2(n_2810),
.B1(n_2796),
.B2(n_2799),
.Y(n_2853)
);

OAI211xp5_ASAP7_75t_L g2854 ( 
.A1(n_2817),
.A2(n_2776),
.B(n_2780),
.C(n_2812),
.Y(n_2854)
);

AOI211xp5_ASAP7_75t_L g2855 ( 
.A1(n_2827),
.A2(n_2812),
.B(n_502),
.C(n_503),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2838),
.B(n_2224),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2819),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2833),
.B(n_501),
.Y(n_2858)
);

NAND3xp33_ASAP7_75t_SL g2859 ( 
.A(n_2830),
.B(n_502),
.C(n_503),
.Y(n_2859)
);

NAND4xp75_ASAP7_75t_L g2860 ( 
.A(n_2834),
.B(n_504),
.C(n_505),
.D(n_506),
.Y(n_2860)
);

NAND4xp75_ASAP7_75t_L g2861 ( 
.A(n_2822),
.B(n_504),
.C(n_505),
.D(n_506),
.Y(n_2861)
);

OR2x2_ASAP7_75t_L g2862 ( 
.A(n_2820),
.B(n_507),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2829),
.Y(n_2863)
);

NOR2xp67_ASAP7_75t_SL g2864 ( 
.A(n_2825),
.B(n_507),
.Y(n_2864)
);

AND2x4_ASAP7_75t_L g2865 ( 
.A(n_2844),
.B(n_508),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2841),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2826),
.Y(n_2867)
);

AOI22xp33_ASAP7_75t_L g2868 ( 
.A1(n_2824),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_2868)
);

INVxp67_ASAP7_75t_L g2869 ( 
.A(n_2839),
.Y(n_2869)
);

NAND3xp33_ASAP7_75t_L g2870 ( 
.A(n_2821),
.B(n_513),
.C(n_514),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2831),
.B(n_514),
.Y(n_2871)
);

AND3x4_ASAP7_75t_L g2872 ( 
.A(n_2840),
.B(n_515),
.C(n_516),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2832),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2835),
.Y(n_2874)
);

NAND3xp33_ASAP7_75t_SL g2875 ( 
.A(n_2837),
.B(n_515),
.C(n_516),
.Y(n_2875)
);

OAI211xp5_ASAP7_75t_SL g2876 ( 
.A1(n_2823),
.A2(n_517),
.B(n_518),
.C(n_519),
.Y(n_2876)
);

AOI22x1_ASAP7_75t_L g2877 ( 
.A1(n_2830),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_2877)
);

AND4x1_ASAP7_75t_L g2878 ( 
.A(n_2815),
.B(n_520),
.C(n_521),
.D(n_522),
.Y(n_2878)
);

OR2x6_ASAP7_75t_L g2879 ( 
.A(n_2830),
.B(n_520),
.Y(n_2879)
);

NAND5xp2_ASAP7_75t_L g2880 ( 
.A(n_2814),
.B(n_521),
.C(n_522),
.D(n_523),
.E(n_524),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2835),
.Y(n_2881)
);

O2A1O1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2830),
.A2(n_523),
.B(n_525),
.C(n_526),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2862),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2879),
.Y(n_2884)
);

AND3x4_ASAP7_75t_L g2885 ( 
.A(n_2846),
.B(n_525),
.C(n_527),
.Y(n_2885)
);

AND4x1_ASAP7_75t_L g2886 ( 
.A(n_2851),
.B(n_527),
.C(n_529),
.D(n_530),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2871),
.B(n_530),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2872),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2879),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2878),
.B(n_531),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2854),
.B(n_531),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2866),
.B(n_532),
.Y(n_2892)
);

NOR3xp33_ASAP7_75t_L g2893 ( 
.A(n_2848),
.B(n_533),
.C(n_534),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2845),
.B(n_535),
.Y(n_2894)
);

NAND3x1_ASAP7_75t_SL g2895 ( 
.A(n_2850),
.B(n_536),
.C(n_537),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2865),
.B(n_536),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2855),
.B(n_2865),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2870),
.Y(n_2898)
);

OAI21xp33_ASAP7_75t_L g2899 ( 
.A1(n_2847),
.A2(n_537),
.B(n_538),
.Y(n_2899)
);

AND3x4_ASAP7_75t_L g2900 ( 
.A(n_2849),
.B(n_538),
.C(n_539),
.Y(n_2900)
);

NOR4xp25_ASAP7_75t_L g2901 ( 
.A(n_2874),
.B(n_2881),
.C(n_2867),
.D(n_2869),
.Y(n_2901)
);

NOR2x2_ASAP7_75t_L g2902 ( 
.A(n_2861),
.B(n_539),
.Y(n_2902)
);

NOR2x1_ASAP7_75t_L g2903 ( 
.A(n_2859),
.B(n_540),
.Y(n_2903)
);

INVxp67_ASAP7_75t_L g2904 ( 
.A(n_2864),
.Y(n_2904)
);

XNOR2x1_ASAP7_75t_SL g2905 ( 
.A(n_2857),
.B(n_540),
.Y(n_2905)
);

NAND4xp75_ASAP7_75t_L g2906 ( 
.A(n_2863),
.B(n_541),
.C(n_542),
.D(n_543),
.Y(n_2906)
);

NOR3xp33_ASAP7_75t_L g2907 ( 
.A(n_2853),
.B(n_541),
.C(n_542),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2891),
.A2(n_2875),
.B1(n_2858),
.B2(n_2876),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2905),
.Y(n_2909)
);

CKINVDCx20_ASAP7_75t_R g2910 ( 
.A(n_2884),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2907),
.A2(n_2873),
.B1(n_2868),
.B2(n_2852),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2896),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2890),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2887),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2906),
.Y(n_2915)
);

OR2x2_ASAP7_75t_L g2916 ( 
.A(n_2892),
.B(n_2880),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2900),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2901),
.B(n_2889),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2885),
.Y(n_2919)
);

OR3x2_ASAP7_75t_L g2920 ( 
.A(n_2895),
.B(n_2882),
.C(n_2860),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_2903),
.A2(n_2856),
.B1(n_2877),
.B2(n_545),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2886),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2893),
.B(n_543),
.Y(n_2923)
);

INVxp67_ASAP7_75t_L g2924 ( 
.A(n_2894),
.Y(n_2924)
);

INVx2_ASAP7_75t_SL g2925 ( 
.A(n_2888),
.Y(n_2925)
);

HB1xp67_ASAP7_75t_L g2926 ( 
.A(n_2897),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2899),
.Y(n_2927)
);

NAND3xp33_ASAP7_75t_L g2928 ( 
.A(n_2918),
.B(n_2904),
.C(n_2883),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2920),
.Y(n_2929)
);

OR3x2_ASAP7_75t_L g2930 ( 
.A(n_2927),
.B(n_2898),
.C(n_2902),
.Y(n_2930)
);

XNOR2x1_ASAP7_75t_L g2931 ( 
.A(n_2916),
.B(n_2926),
.Y(n_2931)
);

XNOR2x1_ASAP7_75t_L g2932 ( 
.A(n_2922),
.B(n_544),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2917),
.Y(n_2933)
);

AND3x4_ASAP7_75t_L g2934 ( 
.A(n_2919),
.B(n_544),
.C(n_545),
.Y(n_2934)
);

OAI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2910),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2923),
.Y(n_2936)
);

XOR2xp5_ASAP7_75t_L g2937 ( 
.A(n_2908),
.B(n_547),
.Y(n_2937)
);

OAI22x1_ASAP7_75t_L g2938 ( 
.A1(n_2911),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_2938)
);

OAI221xp5_ASAP7_75t_L g2939 ( 
.A1(n_2921),
.A2(n_2925),
.B1(n_2909),
.B2(n_2915),
.C(n_2924),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2912),
.Y(n_2940)
);

OAI22x1_ASAP7_75t_L g2941 ( 
.A1(n_2928),
.A2(n_2940),
.B1(n_2914),
.B2(n_2929),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2930),
.A2(n_2913),
.B1(n_550),
.B2(n_551),
.Y(n_2942)
);

OR5x1_ASAP7_75t_L g2943 ( 
.A(n_2931),
.B(n_549),
.C(n_551),
.D(n_552),
.E(n_553),
.Y(n_2943)
);

OAI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2939),
.A2(n_553),
.B(n_554),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2932),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2937),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2933),
.A2(n_554),
.B(n_555),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_SL g2948 ( 
.A1(n_2943),
.A2(n_2936),
.B1(n_2934),
.B2(n_2938),
.Y(n_2948)
);

O2A1O1Ixp33_ASAP7_75t_L g2949 ( 
.A1(n_2945),
.A2(n_2935),
.B(n_557),
.C(n_558),
.Y(n_2949)
);

OAI22xp5_ASAP7_75t_L g2950 ( 
.A1(n_2944),
.A2(n_556),
.B1(n_558),
.B2(n_559),
.Y(n_2950)
);

XNOR2xp5_ASAP7_75t_L g2951 ( 
.A(n_2941),
.B(n_556),
.Y(n_2951)
);

NOR2x1_ASAP7_75t_L g2952 ( 
.A(n_2946),
.B(n_559),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2942),
.B(n_560),
.Y(n_2953)
);

HB1xp67_ASAP7_75t_L g2954 ( 
.A(n_2947),
.Y(n_2954)
);

AO22x1_ASAP7_75t_L g2955 ( 
.A1(n_2952),
.A2(n_560),
.B1(n_561),
.B2(n_562),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2948),
.A2(n_561),
.B(n_562),
.Y(n_2956)
);

A2O1A1Ixp33_ASAP7_75t_L g2957 ( 
.A1(n_2949),
.A2(n_563),
.B(n_564),
.C(n_565),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2953),
.A2(n_563),
.B(n_564),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2956),
.A2(n_2951),
.B1(n_2950),
.B2(n_2954),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2955),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2958),
.A2(n_565),
.B1(n_566),
.B2(n_567),
.Y(n_2961)
);

XNOR2xp5_ASAP7_75t_L g2962 ( 
.A(n_2959),
.B(n_2957),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2960),
.Y(n_2963)
);

OR2x2_ASAP7_75t_L g2964 ( 
.A(n_2961),
.B(n_566),
.Y(n_2964)
);

AOI222xp33_ASAP7_75t_L g2965 ( 
.A1(n_2963),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.C1(n_571),
.C2(n_572),
.Y(n_2965)
);

NAND3xp33_ASAP7_75t_L g2966 ( 
.A(n_2962),
.B(n_571),
.C(n_572),
.Y(n_2966)
);

AOI221xp5_ASAP7_75t_L g2967 ( 
.A1(n_2966),
.A2(n_2964),
.B1(n_574),
.B2(n_576),
.C(n_577),
.Y(n_2967)
);

NOR3x1_ASAP7_75t_L g2968 ( 
.A(n_2967),
.B(n_2965),
.C(n_574),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2968),
.Y(n_2969)
);

OA21x2_ASAP7_75t_L g2970 ( 
.A1(n_2969),
.A2(n_573),
.B(n_577),
.Y(n_2970)
);

OAI221xp5_ASAP7_75t_R g2971 ( 
.A1(n_2970),
.A2(n_573),
.B1(n_578),
.B2(n_579),
.C(n_580),
.Y(n_2971)
);

AOI21xp33_ASAP7_75t_L g2972 ( 
.A1(n_2971),
.A2(n_578),
.B(n_579),
.Y(n_2972)
);

AOI211xp5_ASAP7_75t_L g2973 ( 
.A1(n_2972),
.A2(n_580),
.B(n_581),
.C(n_582),
.Y(n_2973)
);


endmodule