module real_jpeg_15943_n_2 (n_1, n_0, n_2);

input n_1;
input n_0;

output n_2;

wire n_4;
wire n_3;

AND2x6_ASAP7_75t_L g4 ( 
.A(n_0),
.B(n_1),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g2 ( 
.A(n_3),
.Y(n_2)
);

BUFx12_ASAP7_75t_L g3 ( 
.A(n_4),
.Y(n_3)
);


endmodule