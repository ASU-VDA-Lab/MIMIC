module fake_ibex_2037_n_19 (n_4, n_2, n_5, n_6, n_0, n_3, n_1, n_19);

input n_4;
input n_2;
input n_5;
input n_6;
input n_0;
input n_3;
input n_1;

output n_19;

wire n_7;
wire n_17;
wire n_18;
wire n_11;
wire n_13;
wire n_8;
wire n_14;
wire n_9;
wire n_12;
wire n_15;
wire n_10;
wire n_16;

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_6),
.Y(n_8)
);

OAI22xp33_ASAP7_75t_L g9 ( 
.A1(n_2),
.A2(n_4),
.B1(n_0),
.B2(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR4xp25_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

AOI221xp5_ASAP7_75t_L g15 ( 
.A1(n_14),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

OAI22x1_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_8),
.B1(n_11),
.B2(n_0),
.Y(n_18)
);

AOI31xp67_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_16),
.A3(n_17),
.B(n_5),
.Y(n_19)
);


endmodule