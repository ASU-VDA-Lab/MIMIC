module fake_jpeg_13961_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_11),
.B(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_45),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_50),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_32),
.B1(n_43),
.B2(n_38),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_61),
.B1(n_40),
.B2(n_15),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_32),
.B1(n_43),
.B2(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_33),
.B1(n_44),
.B2(n_42),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_5),
.B(n_6),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_33),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_80),
.B1(n_62),
.B2(n_63),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_87),
.A3(n_83),
.B1(n_81),
.B2(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_68),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_84),
.C(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_89),
.B1(n_86),
.B2(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_74),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_85),
.A3(n_10),
.B1(n_14),
.B2(n_16),
.C1(n_18),
.C2(n_7),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_23),
.B(n_26),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_27),
.Y(n_96)
);


endmodule