module fake_jpeg_20148_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_25),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_26),
.B1(n_34),
.B2(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_48),
.B1(n_52),
.B2(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_26),
.B1(n_16),
.B2(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_41),
.B1(n_36),
.B2(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_41),
.B1(n_30),
.B2(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_73),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_80),
.Y(n_100)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_33),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_29),
.B1(n_23),
.B2(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_42),
.B1(n_37),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_82),
.B1(n_49),
.B2(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_42),
.B1(n_37),
.B2(n_20),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_38),
.B(n_37),
.C(n_21),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_58),
.B(n_68),
.C(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_59),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_21),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_38),
.C(n_47),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_87),
.B1(n_49),
.B2(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_101),
.B1(n_70),
.B2(n_74),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_73),
.B1(n_88),
.B2(n_66),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_114),
.B(n_67),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_59),
.C(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_19),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_120),
.B1(n_137),
.B2(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_121),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_100),
.B1(n_92),
.B2(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_80),
.C(n_9),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_112),
.Y(n_143)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_78),
.B1(n_72),
.B2(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_136),
.B1(n_138),
.B2(n_108),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_131),
.B(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_111),
.B(n_109),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_72),
.B1(n_71),
.B2(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_83),
.B1(n_76),
.B2(n_85),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_82),
.B1(n_66),
.B2(n_73),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_11),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_99),
.B(n_113),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_146),
.B(n_152),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_113),
.B(n_93),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_108),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_148),
.B(n_150),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_91),
.B1(n_94),
.B2(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_149),
.A2(n_168),
.B1(n_169),
.B2(n_115),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_93),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_103),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_128),
.B(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_104),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_160),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_94),
.B(n_97),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_111),
.B(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_164),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_104),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_162),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_111),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_66),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_95),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_18),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_7),
.B1(n_15),
.B2(n_12),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_129),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_121),
.B1(n_131),
.B2(n_130),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_132),
.C(n_117),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_182),
.C(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_118),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_118),
.C(n_123),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_115),
.C(n_18),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_162),
.B1(n_155),
.B2(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_155),
.Y(n_199)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

XNOR2x2_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_145),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_183),
.B(n_147),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_144),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_211),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_171),
.B1(n_183),
.B2(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_157),
.B1(n_163),
.B2(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_191),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_193),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_160),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_181),
.C(n_180),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_219),
.B1(n_224),
.B2(n_209),
.Y(n_236)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_230),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_171),
.B1(n_190),
.B2(n_192),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_173),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_166),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_168),
.B1(n_188),
.B2(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_227),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_180),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_210),
.B1(n_205),
.B2(n_208),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_210),
.B1(n_216),
.B2(n_222),
.Y(n_234)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_214),
.C(n_200),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_238),
.C(n_239),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_236),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_214),
.C(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_213),
.C(n_212),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_194),
.B1(n_166),
.B2(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_247),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_219),
.C(n_223),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_216),
.B1(n_228),
.B2(n_226),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_232),
.B1(n_231),
.B2(n_239),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_9),
.B1(n_8),
.B2(n_3),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_1),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_230),
.B1(n_2),
.B2(n_3),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_1),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_12),
.B(n_11),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_9),
.B(n_8),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_1),
.C(n_2),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_246),
.B1(n_248),
.B2(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.C(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_244),
.C(n_247),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_250),
.B(n_260),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_271),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_262),
.C(n_4),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

OAI31xp33_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_272),
.A3(n_5),
.B(n_6),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_5),
.Y(n_276)
);


endmodule