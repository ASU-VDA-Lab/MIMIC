module real_jpeg_16833_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_1),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_90),
.Y(n_171)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_5),
.A2(n_9),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_5),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_5),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_5),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_5),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_5),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_5),
.B(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_7),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_7),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_7),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_7),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_8),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_8),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_8),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_8),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_8),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_8),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_9),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_9),
.B(n_74),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g124 ( 
.A(n_12),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_12),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_14),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_14),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_14),
.B(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_17),
.Y(n_136)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_223),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_183),
.B(n_220),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_25),
.B(n_184),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_112),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_68),
.C(n_94),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_27),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_44),
.C(n_57),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_29),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_30),
.B(n_38),
.C(n_43),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_44),
.B(n_57),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_45),
.B(n_51),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_48),
.Y(n_271)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.C(n_64),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_58),
.B(n_61),
.Y(n_231)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_61),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_61),
.B(n_309),
.C(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_63),
.Y(n_265)
);

XOR2x1_ASAP7_75t_SL g230 ( 
.A(n_64),
.B(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_68),
.B(n_94),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_79),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_77),
.C(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.C(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_80),
.A2(n_89),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_84),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_85),
.B(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_89),
.B(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_101),
.C(n_110),
.Y(n_153)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_105),
.A2(n_110),
.B1(n_234),
.B2(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_110),
.B(n_234),
.C(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_151),
.B1(n_181),
.B2(n_182),
.Y(n_112)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_138),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.C(n_137),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_115),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_121),
.C(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_128),
.A2(n_129),
.B1(n_137),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_129),
.A2(n_193),
.B(n_200),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_138)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_142),
.A2(n_143),
.B1(n_213),
.B2(n_214),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_207),
.C(n_213),
.Y(n_206)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_168),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_160),
.Y(n_167)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_166),
.Y(n_278)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_217),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_217),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.C(n_206),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_192),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_190),
.B(n_259),
.C(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_207),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_SL g293 ( 
.A(n_208),
.B(n_211),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_208),
.A2(n_303),
.B1(n_304),
.B2(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_250),
.B(n_361),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_248),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_226),
.B(n_248),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_245),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_227),
.B(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_229),
.B(n_246),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.C(n_243),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_230),
.B(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_233),
.B(n_244),
.Y(n_346)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_356),
.B(n_360),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_342),
.B(n_355),
.Y(n_253)
);

OAI21x1_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_299),
.B(n_341),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_284),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_256),
.B(n_284),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.C(n_275),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_257),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_268),
.B(n_272),
.Y(n_310)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

AO22x1_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_279),
.B1(n_282),
.B2(n_283),
.Y(n_275)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_279),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_282),
.Y(n_291)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_286),
.B(n_287),
.C(n_290),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_334),
.B(n_340),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_318),
.B(n_333),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_308),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_328),
.B(n_332),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_338),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_354),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_347),
.B2(n_348),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_349),
.C(n_353),
.Y(n_357)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_358),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);


endmodule