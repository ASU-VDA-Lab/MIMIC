module fake_jpeg_14863_n_87 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_87);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx11_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_10),
.Y(n_60)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_40),
.B1(n_43),
.B2(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_42),
.B1(n_37),
.B2(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_32),
.B1(n_14),
.B2(n_17),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_4),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_22),
.B(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_11),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.C(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_70),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_65),
.Y(n_78)
);

BUFx24_ASAP7_75t_SL g77 ( 
.A(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_63),
.C(n_72),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_81),
.A2(n_69),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_56),
.B1(n_26),
.B2(n_29),
.Y(n_87)
);


endmodule