module real_jpeg_32670_n_15 (n_8, n_0, n_2, n_132, n_125, n_10, n_9, n_129, n_12, n_124, n_130, n_134, n_6, n_128, n_133, n_11, n_14, n_131, n_7, n_127, n_3, n_5, n_4, n_1, n_126, n_13, n_15);

input n_8;
input n_0;
input n_2;
input n_132;
input n_125;
input n_10;
input n_9;
input n_129;
input n_12;
input n_124;
input n_130;
input n_134;
input n_6;
input n_128;
input n_133;
input n_11;
input n_14;
input n_131;
input n_7;
input n_127;
input n_3;
input n_5;
input n_4;
input n_1;
input n_126;
input n_13;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI221xp5_ASAP7_75t_L g76 ( 
.A1(n_0),
.A2(n_14),
.B1(n_77),
.B2(n_83),
.C(n_85),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_45),
.A3(n_47),
.B1(n_53),
.B2(n_117),
.C1(n_119),
.C2(n_134),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_79),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_17),
.B1(n_18),
.B2(n_24),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_77),
.C(n_83),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_25),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_34),
.B(n_122),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI31xp67_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_68),
.A3(n_106),
.B(n_112),
.Y(n_35)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_52),
.C(n_61),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_37),
.A2(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_45),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_39),
.B(n_61),
.C(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_125),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

OA21x2_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_97),
.C(n_98),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_89),
.B(n_96),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_130),
.Y(n_83)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_124),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_126),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_127),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_128),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_129),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_131),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_132),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_133),
.Y(n_109)
);


endmodule