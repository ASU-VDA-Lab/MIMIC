module fake_aes_321_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_4), .A2(n_0), .B(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_7), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_16), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_11), .B(n_1), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_12), .B(n_2), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
BUFx12f_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_15), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_13), .B1(n_16), .B2(n_14), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_20), .B(n_17), .Y(n_26) );
AO21x2_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_19), .B(n_20), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_16), .B1(n_18), .B2(n_21), .C(n_22), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_23), .B(n_14), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_27), .B(n_25), .Y(n_31) );
INVx3_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_29), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_33), .B(n_31), .Y(n_34) );
AOI211xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_28), .B(n_16), .C(n_31), .Y(n_35) );
AOI22xp33_ASAP7_75t_SL g36 ( .A1(n_32), .A2(n_18), .B1(n_21), .B2(n_25), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
NOR2x2_ASAP7_75t_L g38 ( .A(n_35), .B(n_5), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_36), .Y(n_39) );
XNOR2xp5_ASAP7_75t_L g40 ( .A(n_39), .B(n_6), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_37), .Y(n_41) );
AOI322xp5_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_8), .A3(n_9), .B1(n_10), .B2(n_37), .C1(n_38), .C2(n_40), .Y(n_42) );
endmodule