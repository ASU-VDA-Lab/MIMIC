module fake_jpeg_7831_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_1),
.B(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_23),
.B1(n_27),
.B2(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_54),
.B1(n_21),
.B2(n_15),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_23),
.B1(n_27),
.B2(n_22),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_51),
.B(n_59),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_23),
.B1(n_31),
.B2(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_21),
.B1(n_41),
.B2(n_29),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_25),
.B1(n_16),
.B2(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_31),
.B1(n_15),
.B2(n_19),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_64),
.Y(n_66)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_76),
.B1(n_48),
.B2(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_79),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_1),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_36),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_72),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_55),
.B1(n_61),
.B2(n_43),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_99),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_43),
.C(n_63),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_107),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_55),
.B1(n_52),
.B2(n_61),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_65),
.B1(n_86),
.B2(n_71),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_36),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_80),
.B1(n_77),
.B2(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_67),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_95),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_35),
.C(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_83),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_84),
.B1(n_83),
.B2(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_117),
.B1(n_127),
.B2(n_2),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_104),
.B1(n_98),
.B2(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_84),
.B1(n_83),
.B2(n_70),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_101),
.B(n_33),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_88),
.B(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_65),
.B1(n_71),
.B2(n_61),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_107),
.B1(n_94),
.B2(n_106),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_65),
.B1(n_55),
.B2(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_66),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_29),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_109),
.B(n_95),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_136),
.B(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_88),
.C(n_81),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_152),
.C(n_117),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_146),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_145),
.CI(n_116),
.CON(n_174),
.SN(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_154),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_30),
.B(n_33),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_30),
.B(n_3),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_127),
.B(n_116),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_98),
.C(n_89),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_3),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_124),
.B1(n_112),
.B2(n_129),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_158),
.B(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_135),
.C(n_134),
.Y(n_181)
);

BUFx12f_ASAP7_75t_SL g164 ( 
.A(n_145),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_167),
.B(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_118),
.CON(n_167),
.SN(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_175),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_174),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_169),
.B1(n_168),
.B2(n_176),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_184),
.B1(n_187),
.B2(n_148),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_192),
.C(n_171),
.Y(n_196)
);

HAxp5_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_137),
.CON(n_206),
.SN(n_206)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_150),
.B1(n_153),
.B2(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_144),
.B1(n_143),
.B2(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_194),
.B(n_122),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_140),
.C(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_164),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_179),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_198),
.C(n_204),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_170),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_201),
.B(n_180),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_175),
.C(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_159),
.B1(n_173),
.B2(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_179),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_160),
.B1(n_159),
.B2(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_174),
.C(n_121),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_194),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_205),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_182),
.C(n_178),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_122),
.C(n_130),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_177),
.B1(n_187),
.B2(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_214),
.B1(n_198),
.B2(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_197),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_217),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_180),
.B(n_189),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_216),
.C(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_178),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_227),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_213),
.Y(n_236)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_235),
.B(n_236),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_230),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_216),
.C(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_231),
.C(n_233),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_224),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_232),
.A2(n_220),
.B1(n_226),
.B2(n_130),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_5),
.C(n_6),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_233),
.B(n_7),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_8),
.B(n_9),
.Y(n_248)
);

AOI321xp33_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_245),
.A3(n_244),
.B1(n_12),
.B2(n_13),
.C(n_11),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_249),
.A2(n_247),
.B(n_12),
.C(n_13),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_9),
.Y(n_251)
);


endmodule