module fake_jpeg_31782_n_366 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_64),
.Y(n_73)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_0),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_31),
.C(n_38),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_8),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_85),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_74),
.A2(n_76),
.B1(n_96),
.B2(n_37),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_95),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_84),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_93),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_16),
.B1(n_17),
.B2(n_40),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_106),
.B1(n_108),
.B2(n_20),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_44),
.B(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_112),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_53),
.A2(n_16),
.B1(n_17),
.B2(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_40),
.B1(n_17),
.B2(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_34),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_46),
.B(n_19),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_66),
.B1(n_63),
.B2(n_46),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_121),
.B1(n_125),
.B2(n_110),
.Y(n_163)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_68),
.B1(n_51),
.B2(n_50),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_32),
.B(n_28),
.C(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_68),
.B1(n_51),
.B2(n_50),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_153),
.B1(n_79),
.B2(n_102),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_47),
.B1(n_23),
.B2(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_28),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_132),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_79),
.B1(n_86),
.B2(n_89),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_81),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_19),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_84),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_135),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_79),
.B1(n_87),
.B2(n_83),
.Y(n_167)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_141),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_49),
.B1(n_56),
.B2(n_26),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_140),
.A2(n_81),
.B1(n_2),
.B2(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_11),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_11),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_94),
.B(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_147),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_49),
.C(n_47),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_151),
.C(n_75),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_37),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_89),
.A2(n_37),
.B1(n_30),
.B2(n_49),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_110),
.A2(n_30),
.B1(n_39),
.B2(n_3),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_83),
.B1(n_113),
.B2(n_94),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_174),
.B1(n_187),
.B2(n_190),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_167),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_178),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_39),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_166),
.B(n_155),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_149),
.B1(n_129),
.B2(n_122),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_91),
.B(n_98),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_140),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_113),
.B1(n_71),
.B2(n_102),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_189),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_183),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_101),
.C(n_107),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_188),
.C(n_193),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_118),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_185),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_119),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_75),
.B1(n_71),
.B2(n_107),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_101),
.C(n_98),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_127),
.B(n_13),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_13),
.C(n_12),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_124),
.B1(n_131),
.B2(n_150),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_197),
.B1(n_225),
.B2(n_190),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_126),
.B(n_154),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_210),
.B(n_159),
.Y(n_238)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_116),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_148),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_217),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_214),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_120),
.B1(n_139),
.B2(n_138),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_169),
.B(n_178),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_147),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_10),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_182),
.B(n_129),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_173),
.B(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_140),
.C(n_144),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_224),
.C(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_153),
.C(n_135),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_163),
.A2(n_119),
.B1(n_12),
.B2(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_1),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_161),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_12),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_178),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_246),
.C(n_221),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_239),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_233),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_166),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_245),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_166),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_240),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_220),
.B(n_210),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_159),
.B1(n_170),
.B2(n_171),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_193),
.C(n_175),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_173),
.B1(n_164),
.B2(n_175),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_249),
.B1(n_254),
.B2(n_211),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_253),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_176),
.B1(n_156),
.B2(n_161),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_209),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_252),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_276),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_272),
.C(n_277),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_261),
.B(n_267),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_247),
.B1(n_254),
.B2(n_237),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_214),
.B(n_195),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_271),
.B(n_236),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_241),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_274),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_213),
.B(n_208),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_223),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_242),
.B(n_207),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.Y(n_287)
);

FAx1_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_224),
.CI(n_226),
.CON(n_274),
.SN(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_279),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_208),
.C(n_200),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_242),
.B(n_201),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_200),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_290),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_239),
.B1(n_231),
.B2(n_236),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_285),
.B1(n_291),
.B2(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_202),
.B1(n_225),
.B2(n_232),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_290),
.B1(n_169),
.B2(n_176),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_202),
.B1(n_255),
.B2(n_233),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_256),
.A2(n_262),
.B1(n_261),
.B2(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_199),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_294),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_260),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_217),
.B1(n_219),
.B2(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_235),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_201),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_169),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_235),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_270),
.B(n_222),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_304),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_259),
.C(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_303),
.C(n_289),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_274),
.C(n_279),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_278),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_271),
.B(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_308),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_286),
.B1(n_288),
.B2(n_282),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_284),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_316),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_294),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_299),
.B1(n_281),
.B2(n_298),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_178),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_303),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_328),
.B1(n_313),
.B2(n_300),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_324),
.A2(n_304),
.B1(n_4),
.B2(n_5),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_310),
.A2(n_289),
.B1(n_156),
.B2(n_177),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_177),
.C(n_156),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_316),
.C(n_301),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_335),
.C(n_329),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_335),
.Y(n_347)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_333),
.Y(n_342)
);

XOR2x2_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_305),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g348 ( 
.A(n_334),
.B(n_6),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_309),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_317),
.C(n_327),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_2),
.B(n_5),
.Y(n_338)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_318),
.B(n_283),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_6),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_341),
.B(n_345),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_324),
.C(n_2),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_330),
.C(n_339),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_342),
.A2(n_332),
.B(n_338),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_353),
.B(n_355),
.Y(n_360)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_347),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_357),
.B(n_358),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_345),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_360),
.A2(n_350),
.B(n_359),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_361),
.A2(n_351),
.B(n_354),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_363),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_362),
.B1(n_331),
.B2(n_347),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_365),
.Y(n_366)
);


endmodule