module fake_ariane_575_n_451 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_451);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_451;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_410;
wire n_379;
wire n_445;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;

BUFx3_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_115),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_17),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_21),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_38),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_44),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_39),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_16),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_49),
.B(n_19),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_50),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_87),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_52),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_34),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_121),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_18),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_113),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_59),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_11),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_61),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_45),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_20),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_69),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_62),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_103),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_64),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_30),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_40),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_12),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_0),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_132),
.B(n_136),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_0),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

CKINVDCx6p67_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_169),
.A2(n_200),
.B1(n_137),
.B2(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_138),
.B(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_174),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

AO21x2_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_133),
.B(n_207),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_209),
.B(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_181),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_172),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_183),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_184),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_147),
.B1(n_165),
.B2(n_142),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_204),
.B1(n_185),
.B2(n_201),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_187),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_192),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_134),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_238),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_148),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_224),
.B1(n_236),
.B2(n_225),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_208),
.B1(n_237),
.B2(n_236),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_223),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_212),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_193),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_258),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

NOR2x1p5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_164),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

NAND2x1_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_197),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_241),
.B(n_199),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_146),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_149),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_153),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_249),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_157),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_263),
.B(n_158),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_146),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_257),
.A2(n_140),
.B(n_156),
.C(n_150),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_265),
.B(n_160),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_255),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_257),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_262),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_288),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_259),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_288),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_260),
.B(n_255),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_260),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_255),
.Y(n_326)
);

BUFx8_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_246),
.B(n_244),
.C(n_253),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_161),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_170),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_276),
.B(n_180),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_245),
.B(n_247),
.C(n_190),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_278),
.B(n_182),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_293),
.A2(n_146),
.B1(n_179),
.B2(n_194),
.Y(n_341)
);

OR2x6_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_242),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_189),
.B1(n_186),
.B2(n_202),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_188),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_4),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_334),
.A2(n_299),
.B1(n_293),
.B2(n_310),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_327),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_299),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_350),
.A2(n_332),
.B1(n_319),
.B2(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_290),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_300),
.B(n_298),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_317),
.A2(n_308),
.B1(n_286),
.B2(n_280),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_297),
.B(n_314),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_335),
.A2(n_297),
.B(n_194),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_194),
.B(n_179),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_331),
.A2(n_194),
.B(n_179),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_314),
.B1(n_7),
.B2(n_5),
.Y(n_365)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_349),
.A2(n_194),
.B(n_179),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_146),
.B(n_14),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_323),
.A2(n_8),
.B(n_15),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_250),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_337),
.A2(n_250),
.B1(n_25),
.B2(n_26),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_316),
.A2(n_29),
.B(n_32),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_33),
.B(n_35),
.Y(n_376)
);

NAND2x1p5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_345),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_366),
.A2(n_326),
.B(n_348),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_355),
.B(n_324),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_342),
.Y(n_381)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_344),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

OAI221xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_343),
.B1(n_322),
.B2(n_320),
.C(n_328),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_328),
.B1(n_345),
.B2(n_348),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_348),
.C(n_37),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_354),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

AO21x2_ASAP7_75t_L g390 ( 
.A1(n_363),
.A2(n_362),
.B(n_361),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_352),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_353),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_369),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_358),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_373),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_373),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_377),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_370),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_403),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_387),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_403),
.Y(n_408)
);

AO31x2_ASAP7_75t_L g409 ( 
.A1(n_396),
.A2(n_388),
.A3(n_390),
.B(n_376),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_375),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_404),
.A2(n_384),
.B1(n_391),
.B2(n_392),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_368),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_394),
.B(n_367),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_360),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_397),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_398),
.Y(n_419)
);

NAND2x1p5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_402),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_402),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_63),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_129),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_417),
.Y(n_428)
);

NOR3xp33_ASAP7_75t_SL g429 ( 
.A(n_421),
.B(n_415),
.C(n_413),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_409),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_422),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_427),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_410),
.Y(n_433)
);

NOR4xp25_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_421),
.C(n_428),
.D(n_425),
.Y(n_434)
);

NAND2x1_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_423),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_433),
.B(n_418),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_432),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

NAND4xp25_ASAP7_75t_SL g440 ( 
.A(n_438),
.B(n_430),
.C(n_424),
.D(n_436),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_426),
.B1(n_409),
.B2(n_79),
.Y(n_441)
);

OAI221xp5_ASAP7_75t_L g442 ( 
.A1(n_440),
.A2(n_409),
.B1(n_73),
.B2(n_80),
.C(n_81),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_72),
.Y(n_443)
);

NOR5xp2_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_84),
.C(n_86),
.D(n_88),
.E(n_89),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_443),
.B(n_91),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_444),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_447),
.Y(n_448)
);

AOI222xp33_ASAP7_75t_SL g449 ( 
.A1(n_448),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.C1(n_101),
.C2(n_104),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_118),
.B1(n_120),
.B2(n_123),
.Y(n_451)
);


endmodule