module fake_jpeg_12262_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_41),
.Y(n_76)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_58),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_28),
.B(n_34),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_27),
.B(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_13),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_2),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_62),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_63),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_15),
.A2(n_5),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_5),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_25),
.B1(n_29),
.B2(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_45),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_22),
.B1(n_20),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_74),
.B1(n_91),
.B2(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_89),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_14),
.B1(n_21),
.B2(n_27),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_5),
.B1(n_27),
.B2(n_44),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_96),
.C(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_37),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_60),
.B1(n_47),
.B2(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_46),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_39),
.B(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_82),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_107),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_67),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_119),
.B(n_112),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_118),
.B(n_120),
.C(n_121),
.D(n_69),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_81),
.C(n_69),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_73),
.B(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_87),
.B1(n_68),
.B2(n_94),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_130),
.B1(n_133),
.B2(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_94),
.B1(n_80),
.B2(n_70),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_80),
.B1(n_93),
.B2(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_145),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_108),
.B1(n_106),
.B2(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_141),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_134),
.B(n_133),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_118),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_136),
.B(n_128),
.C(n_141),
.D(n_121),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_103),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_119),
.C(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_142),
.C(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_141),
.B1(n_125),
.B2(n_135),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_150),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_144),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_149),
.B(n_138),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_129),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_148),
.C(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_109),
.B1(n_155),
.B2(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_142),
.B1(n_157),
.B2(n_102),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_162),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_164),
.B1(n_163),
.B2(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_102),
.B(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_117),
.C(n_169),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_168),
.C(n_171),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_174),
.Y(n_177)
);


endmodule