module fake_jpeg_11766_n_42 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_42);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_42;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_1),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_15),
.C(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B(n_2),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_30),
.B(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_15),
.B1(n_14),
.B2(n_16),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_12),
.B1(n_11),
.B2(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_3),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_3),
.B(n_4),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.C(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_5),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_34),
.B(n_7),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_6),
.C(n_8),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_9),
.B(n_10),
.C(n_31),
.Y(n_42)
);


endmodule