module real_jpeg_4105_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_27),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_76),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_1),
.A2(n_76),
.B1(n_149),
.B2(n_325),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_1),
.A2(n_76),
.B1(n_347),
.B2(n_350),
.Y(n_346)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_26),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_31),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_26),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_3),
.A2(n_26),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_3),
.A2(n_313),
.B(n_315),
.C(n_319),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_3),
.B(n_337),
.C(n_339),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_3),
.B(n_120),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_3),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_3),
.B(n_134),
.Y(n_376)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_5),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_5),
.Y(n_364)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_5),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_47),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_47),
.B1(n_173),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_47),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_7),
.Y(n_158)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_10),
.Y(n_430)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_11),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_167),
.B1(n_168),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_13),
.A2(n_167),
.B1(n_241),
.B2(n_245),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_13),
.A2(n_167),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_13),
.A2(n_167),
.B1(n_427),
.B2(n_431),
.Y(n_426)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_456),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_61),
.B1(n_65),
.B2(n_451),
.C(n_454),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_22),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_22),
.B(n_61),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_23),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_24),
.B(n_218),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_50),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g315 ( 
.A1(n_26),
.A2(n_316),
.B(n_318),
.Y(n_315)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_28),
.Y(n_160)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_31),
.B(n_44),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_35),
.Y(n_162)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_37),
.Y(n_156)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_43),
.B(n_74),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_43),
.A2(n_63),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_50),
.B(n_75),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_53),
.Y(n_432)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_55),
.Y(n_164)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_61),
.A2(n_267),
.B1(n_273),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_61),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_61),
.A2(n_273),
.B(n_279),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_62),
.A2(n_217),
.B(n_426),
.Y(n_447)
);

A2O1A1O1Ixp25_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_405),
.B(n_440),
.C(n_443),
.D(n_450),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_397),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_255),
.C(n_302),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_228),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_200),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_70),
.B(n_200),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_152),
.C(n_184),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_71),
.B(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_72),
.B(n_79),
.C(n_122),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_73),
.B(n_217),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_121),
.B1(n_122),
.B2(n_151),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_114),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_81),
.A2(n_120),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_81),
.B(n_221),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_107),
.Y(n_81)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_82),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_97),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_87),
.Y(n_317)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_90),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_90),
.Y(n_289)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_97),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_101),
.Y(n_246)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_101),
.Y(n_327)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_106),
.Y(n_314)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_108),
.B(n_120),
.Y(n_186)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_113),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_114),
.B(n_265),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_115),
.B(n_188),
.Y(n_187)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_120),
.A2(n_188),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_121),
.A2(n_122),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_121),
.B(n_412),
.C(n_415),
.Y(n_438)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_122),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_122),
.B(n_436),
.C(n_437),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_143),
.B(n_144),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_123),
.A2(n_207),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_145),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_124),
.B(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_124),
.B(n_324),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_135),
.B1(n_137),
.B2(n_141),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_133),
.Y(n_244)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_134),
.B(n_324),
.Y(n_341)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_138),
.Y(n_350)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_142),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_142),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_143),
.A2(n_240),
.B(n_247),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_143),
.B(n_144),
.Y(n_294)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_148),
.Y(n_335)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_152),
.A2(n_153),
.B1(n_184),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_165),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_154),
.B(n_165),
.Y(n_214)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.A3(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_175),
.B(n_177),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_199),
.B(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_178),
.A2(n_193),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_178),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_182),
.Y(n_199)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_185),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_186),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_186),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_188),
.B(n_223),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_188),
.A2(n_287),
.B(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_191),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_192),
.B(n_362),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_199),
.B(n_345),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_200),
.B(n_229),
.Y(n_401)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.CI(n_213),
.CON(n_200),
.SN(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_205),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_206),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_207),
.B(n_323),
.Y(n_352)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.C(n_219),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_228),
.A2(n_400),
.B(n_401),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_232),
.C(n_248),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_248),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_234),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_238),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_247),
.B(n_341),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_251),
.A2(n_253),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_251),
.B(n_447),
.C(n_448),
.Y(n_453)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_298),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_256),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_275),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_257),
.B(n_275),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.C(n_274),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_266),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_272),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_267),
.A2(n_273),
.B1(n_312),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_297),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_285),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_278),
.B(n_284),
.C(n_297),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_293),
.B(n_296),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_293),
.Y(n_296)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_296),
.A2(n_409),
.B1(n_410),
.B2(n_417),
.Y(n_408)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_296),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_299),
.B(n_301),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_328),
.B(n_396),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_304),
.B(n_307),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.C(n_320),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_308),
.B(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_311),
.A2(n_320),
.B1(n_321),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_390),
.B(n_395),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_380),
.B(n_389),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_356),
.B(n_379),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_342),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_332),
.B(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_340),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_334),
.B1(n_340),
.B2(n_359),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_354),
.C(n_382),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_365),
.B(n_378),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_360),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_374),
.B(n_377),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_373),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_376),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_394),
.Y(n_395)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_399),
.B(n_402),
.C(n_403),
.D(n_404),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_420),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_419),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_419),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_418),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_417),
.C(n_418),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_411),
.A2(n_412),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_423),
.C(n_438),
.Y(n_449)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_439),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_439),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_438),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_433),
.B1(n_434),
.B2(n_437),
.Y(n_424)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_425),
.Y(n_437)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_449),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_449),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_453),
.Y(n_455)
);


endmodule