module real_jpeg_23916_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_49),
.B1(n_53),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_33),
.B1(n_49),
.B2(n_53),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_23),
.C(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_6),
.B(n_37),
.C(n_39),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_49),
.C(n_62),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_6),
.B(n_101),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_111),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_109),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_88),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_14),
.B(n_88),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_67),
.C(n_77),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_16),
.B1(n_67),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_46),
.B2(n_66),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_17),
.A2(n_18),
.B1(n_123),
.B2(n_130),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_17),
.A2(n_18),
.B1(n_78),
.B2(n_79),
.Y(n_199)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_34),
.B2(n_45),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_45),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_19),
.A2(n_20),
.B1(n_68),
.B2(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_19),
.A2(n_20),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_34),
.Y(n_86)
);

AOI211xp5_ASAP7_75t_L g120 ( 
.A1(n_20),
.A2(n_58),
.B(n_87),
.C(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_22),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_27),
.B1(n_37),
.B2(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_23),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_34),
.A2(n_45),
.B1(n_58),
.B2(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_34),
.B(n_124),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_34),
.A2(n_45),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_34),
.A2(n_58),
.B(n_121),
.C(n_185),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_36),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_36)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_39),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_39),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_98),
.B(n_104),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_45),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_45),
.B(n_119),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_86),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_47),
.A2(n_58),
.B1(n_119),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_52),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_49),
.B(n_174),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_80),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_58),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_58),
.A2(n_119),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_58),
.A2(n_119),
.B1(n_161),
.B2(n_162),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_58),
.A2(n_119),
.B1(n_149),
.B2(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_64),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_82),
.Y(n_125)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_77),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_87),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_86),
.A2(n_107),
.B(n_123),
.Y(n_202)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_204),
.B(n_209),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_142),
.B(n_195),
.C(n_203),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_132),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_132),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_122),
.B2(n_131),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_120),
.C(n_131),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_146),
.C(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_125),
.C(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_125),
.B1(n_139),
.B2(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_125),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_124),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_124),
.A2(n_125),
.B1(n_150),
.B2(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_125),
.B(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_137),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_134),
.A2(n_135),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_194),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_156),
.B(n_193),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_145),
.B(n_153),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_187),
.B(n_192),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_181),
.B(n_186),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_170),
.B(n_180),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_164),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_208),
.Y(n_209)
);


endmodule