module fake_ariane_3246_n_1605 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1605);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1605;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_5),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_21),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_35),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_26),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_43),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_27),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_35),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_22),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_38),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_42),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_30),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_85),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_40),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_90),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_29),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_45),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_89),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_57),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_20),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_44),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_57),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_44),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_31),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_32),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_28),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_61),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_58),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_36),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_114),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_39),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_28),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_105),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_100),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_59),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_46),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_60),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_56),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_39),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_102),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_108),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_58),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_50),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_54),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_80),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_72),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_49),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_81),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_99),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_43),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_118),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_87),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_71),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_5),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_145),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_67),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_11),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_133),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_16),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_75),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_141),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_110),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_65),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_78),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_131),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_129),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_88),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_36),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_12),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_111),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_1),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_206),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_184),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_168),
.B(n_193),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_221),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_155),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_147),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_157),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_151),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_212),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_151),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_219),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_157),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_231),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_156),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_266),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_214),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_166),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_268),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_269),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_172),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_172),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_214),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_170),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_260),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_168),
.B(n_1),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_148),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_260),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_149),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_186),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_170),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_194),
.B(n_3),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_177),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_194),
.B(n_3),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_150),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_202),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_179),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_202),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_207),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_207),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_154),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_173),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_222),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_162),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_158),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_200),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_179),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_256),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_213),
.B(n_4),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_181),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_213),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_8),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_220),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_222),
.B(n_10),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_274),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_280),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_163),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_158),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_181),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_216),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_208),
.B(n_11),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_188),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_290),
.B(n_160),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_295),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_299),
.A2(n_236),
.B(n_217),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_314),
.B(n_167),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_299),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_160),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_337),
.B(n_163),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_291),
.B(n_208),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_291),
.B(n_217),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_321),
.B(n_236),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_352),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_287),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_350),
.A2(n_230),
.B1(n_285),
.B2(n_284),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

NOR2x1_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_164),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_252),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_331),
.B(n_160),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_325),
.A2(n_229),
.B1(n_281),
.B2(n_278),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_303),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_333),
.A2(n_254),
.B(n_252),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_164),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_164),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_355),
.B(n_254),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_335),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_355),
.B(n_258),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_288),
.A2(n_246),
.B1(n_175),
.B2(n_180),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_425),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_354),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_354),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_320),
.B1(n_289),
.B2(n_329),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_380),
.A2(n_346),
.B1(n_349),
.B2(n_327),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

CKINVDCx11_ASAP7_75t_R g441 ( 
.A(n_401),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_337),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_317),
.B1(n_351),
.B2(n_358),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_324),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_376),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_357),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_377),
.B(n_330),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_395),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_409),
.B(n_351),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

NAND2x1p5_ASAP7_75t_L g458 ( 
.A(n_369),
.B(n_357),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_376),
.B(n_336),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_362),
.B(n_327),
.C(n_359),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_374),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_379),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_364),
.B(n_258),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_317),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_366),
.B(n_306),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_364),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_395),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_380),
.A2(n_306),
.B1(n_358),
.B2(n_316),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_367),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_367),
.B(n_339),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_409),
.A2(n_293),
.B1(n_311),
.B2(n_310),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_368),
.B(n_340),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_372),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_372),
.B(n_292),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_369),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_369),
.A2(n_360),
.B1(n_356),
.B2(n_292),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_410),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_375),
.B(n_222),
.C(n_261),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_398),
.B(n_322),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_383),
.B(n_294),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_383),
.B(n_294),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_361),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_384),
.B(n_386),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_386),
.B(n_296),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_390),
.B(n_296),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_410),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_391),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_428),
.A2(n_332),
.B1(n_347),
.B2(n_302),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_391),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_361),
.B(n_302),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_393),
.B(n_152),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_312),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_396),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_389),
.A2(n_332),
.B1(n_347),
.B2(n_312),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_401),
.B(n_169),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_402),
.B(n_313),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_405),
.B(n_313),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_411),
.B(n_328),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_369),
.A2(n_360),
.B1(n_356),
.B2(n_344),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_416),
.Y(n_530)
);

INVxp67_ASAP7_75t_R g531 ( 
.A(n_400),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_407),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_412),
.A2(n_262),
.B(n_261),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_416),
.B(n_264),
.C(n_262),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_361),
.B(n_328),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_417),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_417),
.B(n_270),
.C(n_264),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_369),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_370),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_408),
.A2(n_344),
.B1(n_210),
.B2(n_209),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_414),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_414),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_400),
.B(n_188),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_408),
.B(n_235),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_370),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_378),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_424),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_408),
.B(n_169),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_424),
.B(n_298),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_408),
.B(n_169),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_363),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_407),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_408),
.B(n_169),
.Y(n_559)
);

AO21x2_ASAP7_75t_L g560 ( 
.A1(n_412),
.A2(n_273),
.B(n_270),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_423),
.Y(n_561)
);

AND3x2_ASAP7_75t_L g562 ( 
.A(n_370),
.B(n_192),
.C(n_189),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_423),
.B(n_277),
.C(n_273),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_406),
.B(n_195),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_426),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_406),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_426),
.B(n_204),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_414),
.A2(n_195),
.B1(n_209),
.B2(n_210),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_414),
.A2(n_232),
.B1(n_224),
.B2(n_259),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_414),
.B(n_235),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_378),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_433),
.B(n_412),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_422),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_422),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_300),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_444),
.A2(n_286),
.B1(n_277),
.B2(n_422),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_532),
.B(n_414),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_432),
.B(n_171),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_561),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_431),
.B(n_182),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_432),
.B(n_171),
.Y(n_582)
);

AOI221xp5_ASAP7_75t_L g583 ( 
.A1(n_506),
.A2(n_229),
.B1(n_232),
.B2(n_224),
.C(n_197),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_498),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_561),
.B(n_565),
.Y(n_586)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_470),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_523),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_517),
.Y(n_591)
);

O2A1O1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_497),
.A2(n_189),
.B(n_243),
.C(n_248),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_432),
.B(n_404),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_456),
.A2(n_242),
.B1(n_243),
.B2(n_238),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_497),
.A2(n_278),
.B(n_248),
.C(n_242),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_436),
.A2(n_247),
.B(n_192),
.C(n_238),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_432),
.B(n_185),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_565),
.B(n_404),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_523),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_482),
.B(n_422),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_448),
.B(n_545),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_447),
.B(n_187),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_485),
.B(n_422),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_436),
.A2(n_422),
.B1(n_307),
.B2(n_304),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_422),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_247),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_460),
.B(n_247),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_510),
.B(n_197),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_487),
.A2(n_281),
.B(n_404),
.C(n_394),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_448),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_448),
.B(n_536),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_472),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_448),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_456),
.A2(n_343),
.B1(n_353),
.B2(n_345),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_473),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_442),
.B(n_196),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_522),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_536),
.B(n_198),
.Y(n_623)
);

OAI221xp5_ASAP7_75t_L g624 ( 
.A1(n_439),
.A2(n_225),
.B1(n_240),
.B2(n_251),
.C(n_199),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_443),
.A2(n_183),
.B1(n_161),
.B2(n_282),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_496),
.B(n_501),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_467),
.B(n_475),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_201),
.Y(n_628)
);

BUFx8_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_522),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_502),
.B(n_203),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_521),
.B(n_218),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_468),
.Y(n_634)
);

INVx8_ASAP7_75t_L g635 ( 
.A(n_467),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_545),
.B(n_404),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_445),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_527),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_475),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_553),
.B(n_165),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_524),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_538),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_525),
.B(n_234),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_554),
.B(n_165),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_526),
.A2(n_404),
.B(n_403),
.C(n_394),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_L g647 ( 
.A1(n_499),
.A2(n_275),
.B(n_263),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_453),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_503),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_489),
.B(n_528),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_462),
.A2(n_276),
.B1(n_265),
.B2(n_272),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_566),
.B(n_204),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_545),
.B(n_274),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_538),
.Y(n_654)
);

AND2x6_ASAP7_75t_SL g655 ( 
.A(n_441),
.B(n_204),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_467),
.A2(n_226),
.B1(n_249),
.B2(n_223),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_559),
.B(n_223),
.Y(n_657)
);

BUFx8_ASAP7_75t_L g658 ( 
.A(n_550),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_494),
.B(n_223),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_564),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_458),
.B(n_274),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_223),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_467),
.A2(n_226),
.B1(n_249),
.B2(n_239),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_481),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_484),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_484),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_486),
.B(n_174),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_446),
.A2(n_403),
.B(n_394),
.C(n_381),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_453),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_547),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_555),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_462),
.B(n_12),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_L g674 ( 
.A(n_477),
.B(n_176),
.C(n_178),
.Y(n_674)
);

NAND2x1p5_ASAP7_75t_L g675 ( 
.A(n_463),
.B(n_165),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_490),
.B(n_190),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_445),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_463),
.B(n_13),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_458),
.B(n_274),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_490),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_SL g681 ( 
.A(n_477),
.B(n_191),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_540),
.B(n_378),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_531),
.B(n_226),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_540),
.B(n_378),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_547),
.B(n_13),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_449),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_540),
.B(n_378),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_249),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_491),
.B(n_239),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_505),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_507),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_507),
.B(n_205),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_540),
.B(n_378),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_450),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_509),
.B(n_211),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_518),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_564),
.B(n_239),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_491),
.B(n_479),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_488),
.B(n_440),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_518),
.A2(n_403),
.B(n_381),
.C(n_373),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_450),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_483),
.B(n_283),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_562),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_529),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_529),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_530),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_459),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_488),
.B(n_378),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_467),
.A2(n_563),
.B1(n_564),
.B2(n_544),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_537),
.B(n_215),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_467),
.B(n_537),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_541),
.B(n_542),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_541),
.B(n_15),
.Y(n_715)
);

BUFx8_ASAP7_75t_L g716 ( 
.A(n_467),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_542),
.Y(n_717)
);

NAND2x1_ASAP7_75t_L g718 ( 
.A(n_519),
.B(n_363),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_549),
.A2(n_283),
.B(n_371),
.C(n_373),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_552),
.B(n_267),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_548),
.B(n_283),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_543),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_552),
.B(n_257),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_611),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_576),
.Y(n_725)
);

INVx11_ASAP7_75t_L g726 ( 
.A(n_629),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_602),
.B(n_548),
.Y(n_727)
);

AOI21x1_ASAP7_75t_L g728 ( 
.A1(n_661),
.A2(n_457),
.B(n_464),
.Y(n_728)
);

AOI33xp33_ASAP7_75t_L g729 ( 
.A1(n_671),
.A2(n_515),
.A3(n_548),
.B1(n_455),
.B2(n_457),
.B3(n_454),
.Y(n_729)
);

AND2x2_ASAP7_75t_SL g730 ( 
.A(n_627),
.B(n_569),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_572),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_634),
.B(n_543),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_670),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_629),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_710),
.A2(n_465),
.B(n_459),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_636),
.B(n_564),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_613),
.B(n_488),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_710),
.A2(n_480),
.B(n_504),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_687),
.A2(n_461),
.B1(n_535),
.B2(n_539),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_596),
.A2(n_511),
.B(n_454),
.C(n_455),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_581),
.B(n_626),
.Y(n_741)
);

AOI21x1_ASAP7_75t_L g742 ( 
.A1(n_661),
.A2(n_464),
.B(n_469),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_613),
.B(n_519),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_613),
.B(n_519),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_629),
.Y(n_745)
);

AOI33xp33_ASAP7_75t_L g746 ( 
.A1(n_594),
.A2(n_568),
.A3(n_474),
.B1(n_492),
.B2(n_471),
.B3(n_500),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_700),
.B(n_564),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_683),
.A2(n_480),
.B(n_478),
.Y(n_748)
);

AO21x1_ASAP7_75t_L g749 ( 
.A1(n_573),
.A2(n_570),
.B(n_434),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_715),
.A2(n_535),
.B(n_539),
.C(n_563),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_603),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_581),
.B(n_520),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_587),
.B(n_452),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_520),
.Y(n_754)
);

INVx11_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_683),
.A2(n_480),
.B(n_474),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_686),
.A2(n_492),
.B(n_500),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_714),
.A2(n_452),
.B1(n_534),
.B2(n_504),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_452),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_677),
.Y(n_761)
);

NAND2x1_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_534),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_613),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_686),
.A2(n_508),
.B(n_434),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_689),
.A2(n_469),
.B(n_430),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_689),
.A2(n_451),
.B(n_430),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_597),
.B(n_435),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_715),
.A2(n_493),
.B(n_451),
.C(n_435),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_624),
.B(n_493),
.C(n_438),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_616),
.B(n_440),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_677),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_649),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_695),
.A2(n_440),
.B(n_533),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_665),
.A2(n_615),
.B(n_619),
.C(n_617),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_557),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_640),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_620),
.B(n_557),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

BUFx2_ASAP7_75t_SL g779 ( 
.A(n_639),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_628),
.A2(n_440),
.B1(n_560),
.B2(n_533),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_591),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_716),
.B(n_600),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_618),
.A2(n_227),
.B1(n_237),
.B2(n_241),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_614),
.B(n_605),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_663),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_701),
.A2(n_440),
.B(n_560),
.Y(n_786)
);

AND2x2_ASAP7_75t_SL g787 ( 
.A(n_713),
.B(n_551),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_652),
.B(n_560),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_721),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_666),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_722),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_578),
.A2(n_546),
.B(n_512),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_638),
.B(n_546),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_606),
.A2(n_546),
.B(n_512),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_667),
.A2(n_571),
.B1(n_551),
.B2(n_546),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_658),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_635),
.B(n_571),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_716),
.B(n_571),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_701),
.A2(n_571),
.B(n_551),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_652),
.B(n_571),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_647),
.A2(n_271),
.B(n_245),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_716),
.B(n_551),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_677),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_637),
.A2(n_551),
.B(n_546),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_685),
.A2(n_512),
.B1(n_437),
.B2(n_244),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_610),
.B(n_512),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_610),
.B(n_512),
.Y(n_808)
);

BUFx12f_ASAP7_75t_SL g809 ( 
.A(n_645),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_15),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_637),
.A2(n_437),
.B(n_373),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_598),
.A2(n_437),
.B(n_381),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_692),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_677),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_693),
.A2(n_437),
.B1(n_250),
.B2(n_279),
.Y(n_815)
);

OAI21xp33_ASAP7_75t_L g816 ( 
.A1(n_673),
.A2(n_253),
.B(n_255),
.Y(n_816)
);

OAI321xp33_ASAP7_75t_L g817 ( 
.A1(n_583),
.A2(n_371),
.A3(n_385),
.B1(n_388),
.B2(n_392),
.C(n_397),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_584),
.B(n_585),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_588),
.B(n_17),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_623),
.B(n_632),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_621),
.Y(n_822)
);

BUFx2_ASAP7_75t_SL g823 ( 
.A(n_721),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_698),
.A2(n_392),
.B(n_388),
.C(n_385),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_18),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_644),
.B(n_18),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_593),
.A2(n_397),
.B(n_392),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_684),
.B(n_19),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_622),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_593),
.A2(n_397),
.B(n_392),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_706),
.A2(n_397),
.B1(n_392),
.B2(n_388),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_658),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_24),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_641),
.B(n_25),
.Y(n_834)
);

AOI21xp33_ASAP7_75t_L g835 ( 
.A1(n_659),
.A2(n_25),
.B(n_26),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_604),
.B(n_635),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_691),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_641),
.B(n_31),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_679),
.A2(n_388),
.B(n_385),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_579),
.A2(n_388),
.B(n_385),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_641),
.B(n_707),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_582),
.A2(n_33),
.B(n_34),
.C(n_41),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_609),
.A2(n_385),
.B(n_46),
.C(n_47),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_635),
.B(n_385),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_699),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_601),
.A2(n_86),
.B(n_143),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_574),
.A2(n_83),
.B(n_140),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_688),
.A2(n_79),
.B(n_137),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_659),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_708),
.B(n_717),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_575),
.B(n_48),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_91),
.B(n_135),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_589),
.B(n_51),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_674),
.B(n_51),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_590),
.B(n_52),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_696),
.A2(n_92),
.B(n_127),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_673),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_678),
.A2(n_711),
.B1(n_709),
.B2(n_599),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_R g859 ( 
.A(n_655),
.B(n_101),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_709),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_696),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_705),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_703),
.B(n_56),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_678),
.A2(n_60),
.B(n_62),
.C(n_74),
.Y(n_864)
);

CKINVDCx6p67_ASAP7_75t_R g865 ( 
.A(n_645),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_607),
.B(n_62),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_669),
.A2(n_106),
.B(n_122),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_703),
.A2(n_123),
.B(n_126),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_646),
.A2(n_146),
.B(n_675),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_718),
.A2(n_668),
.B(n_720),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_699),
.B(n_721),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_657),
.B(n_662),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_630),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_699),
.B(n_645),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_657),
.B(n_662),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_625),
.B(n_660),
.Y(n_876)
);

AOI21x1_ASAP7_75t_L g877 ( 
.A1(n_653),
.A2(n_642),
.B(n_672),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_704),
.B(n_723),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_651),
.B(n_694),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_630),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_681),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_L g882 ( 
.A(n_592),
.B(n_595),
.C(n_712),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_675),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_676),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_631),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_872),
.A2(n_697),
.B(n_612),
.C(n_719),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_741),
.A2(n_653),
.B(n_702),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_726),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_875),
.A2(n_577),
.B(n_656),
.C(n_664),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_821),
.B(n_747),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_789),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_854),
.A2(n_643),
.B(n_672),
.C(n_631),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_884),
.B(n_650),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_724),
.Y(n_894)
);

OR2x6_ASAP7_75t_SL g895 ( 
.A(n_862),
.B(n_755),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_835),
.A2(n_642),
.B(n_654),
.C(n_682),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_SL g897 ( 
.A(n_779),
.B(n_654),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_809),
.B(n_797),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_747),
.B(n_878),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_772),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_787),
.B(n_754),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_751),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_850),
.A2(n_774),
.B1(n_841),
.B2(n_760),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_784),
.A2(n_750),
.B(n_879),
.C(n_774),
.Y(n_904)
);

O2A1O1Ixp5_ASAP7_75t_L g905 ( 
.A1(n_867),
.A2(n_869),
.B(n_851),
.C(n_749),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_784),
.A2(n_732),
.B1(n_725),
.B2(n_791),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_819),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_753),
.B(n_760),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_L g909 ( 
.A1(n_851),
.A2(n_863),
.B(n_767),
.C(n_843),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_832),
.B(n_734),
.Y(n_910)
);

O2A1O1Ixp5_ASAP7_75t_SL g911 ( 
.A1(n_863),
.A2(n_737),
.B(n_866),
.C(n_788),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_733),
.B(n_731),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_857),
.A2(n_864),
.B(n_833),
.C(n_828),
.Y(n_913)
);

OA22x2_ASAP7_75t_L g914 ( 
.A1(n_783),
.A2(n_837),
.B1(n_736),
.B2(n_849),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_857),
.B(n_864),
.C(n_739),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_756),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_753),
.B(n_729),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_752),
.A2(n_870),
.B(n_801),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_874),
.A2(n_876),
.B1(n_730),
.B2(n_871),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_750),
.A2(n_820),
.B(n_825),
.C(n_826),
.Y(n_920)
);

XNOR2xp5_ASAP7_75t_L g921 ( 
.A(n_745),
.B(n_874),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_799),
.B(n_803),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_731),
.B(n_876),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_773),
.A2(n_766),
.B(n_765),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_776),
.B(n_785),
.Y(n_925)
);

BUFx2_ASAP7_75t_SL g926 ( 
.A(n_871),
.Y(n_926)
);

AO32x1_ASAP7_75t_L g927 ( 
.A1(n_858),
.A2(n_831),
.A3(n_759),
.B1(n_861),
.B2(n_883),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_764),
.A2(n_758),
.B(n_800),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_881),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_739),
.A2(n_730),
.B1(n_882),
.B2(n_790),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_786),
.A2(n_742),
.B(n_877),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_881),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_789),
.B(n_845),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_882),
.B(n_816),
.C(n_842),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_796),
.A2(n_813),
.B1(n_787),
.B2(n_860),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_860),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_853),
.A2(n_855),
.B(n_810),
.C(n_838),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_818),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_860),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_798),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_818),
.Y(n_942)
);

NAND2x1_ASAP7_75t_SL g943 ( 
.A(n_763),
.B(n_780),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_823),
.B(n_775),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_768),
.A2(n_757),
.B(n_748),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_860),
.A2(n_777),
.B1(n_834),
.B2(n_763),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_778),
.A2(n_885),
.B1(n_880),
.B2(n_873),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_799),
.B(n_803),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_738),
.A2(n_735),
.B(n_737),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_740),
.A2(n_802),
.B(n_824),
.C(n_770),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_819),
.B(n_746),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_761),
.B(n_814),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_761),
.B(n_814),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_819),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_761),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_781),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_769),
.A2(n_847),
.B(n_817),
.C(n_839),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_859),
.B(n_819),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_771),
.B(n_814),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_822),
.A2(n_829),
.B1(n_769),
.B2(n_807),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_771),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_836),
.A2(n_770),
.B(n_805),
.Y(n_963)
);

AOI33xp33_ASAP7_75t_L g964 ( 
.A1(n_859),
.A2(n_743),
.A3(n_744),
.B1(n_830),
.B2(n_827),
.B3(n_728),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_743),
.A2(n_744),
.B1(n_808),
.B2(n_771),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_804),
.B(n_814),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_804),
.Y(n_967)
);

BUFx6f_ASAP7_75t_SL g968 ( 
.A(n_804),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_844),
.B(n_804),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_782),
.B(n_815),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_782),
.A2(n_795),
.B1(n_844),
.B2(n_806),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_762),
.B(n_793),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_846),
.B(n_868),
.C(n_856),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_844),
.B(n_793),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_844),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_844),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_794),
.A2(n_792),
.B(n_811),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_812),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_848),
.B(n_852),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_741),
.A2(n_875),
.B1(n_872),
.B2(n_727),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_872),
.B(n_431),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_751),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_799),
.B(n_803),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_751),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_741),
.B(n_602),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_732),
.B(n_366),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_741),
.B(n_602),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_741),
.A2(n_586),
.B(n_580),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_741),
.A2(n_586),
.B(n_580),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_741),
.B(n_602),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_SL g992 ( 
.A1(n_783),
.A2(n_477),
.B1(n_491),
.B2(n_453),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_872),
.A2(n_875),
.B(n_602),
.C(n_431),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_860),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_741),
.B(n_602),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_860),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_872),
.A2(n_602),
.B1(n_477),
.B2(n_491),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_872),
.B(n_431),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_741),
.B(n_602),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_741),
.A2(n_875),
.B1(n_872),
.B2(n_727),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_761),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_823),
.B(n_797),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_872),
.A2(n_875),
.B(n_602),
.C(n_431),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_797),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_872),
.A2(n_875),
.B(n_602),
.C(n_431),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_809),
.B(n_453),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_726),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_761),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_787),
.B(n_727),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_867),
.A2(n_869),
.B(n_851),
.C(n_749),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_741),
.A2(n_586),
.B(n_580),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_741),
.A2(n_875),
.B1(n_872),
.B2(n_727),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_431),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_786),
.A2(n_773),
.B(n_766),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_982),
.B(n_998),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_900),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_894),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_1007),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_SL g1021 ( 
.A1(n_913),
.A2(n_938),
.B(n_930),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_890),
.A2(n_915),
.B1(n_1014),
.B2(n_982),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_981),
.A2(n_1013),
.B(n_1000),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_993),
.A2(n_1005),
.B(n_1003),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_898),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_1014),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_986),
.A2(n_991),
.B(n_988),
.C(n_995),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_999),
.B(n_890),
.Y(n_1029)
);

AO32x2_ASAP7_75t_L g1030 ( 
.A1(n_935),
.A2(n_946),
.A3(n_903),
.B1(n_915),
.B2(n_965),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_987),
.B(n_997),
.Y(n_1031)
);

BUFx4f_ASAP7_75t_L g1032 ( 
.A(n_1002),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_SL g1033 ( 
.A1(n_930),
.A2(n_917),
.B(n_950),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_980),
.A2(n_904),
.B(n_941),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_980),
.A2(n_924),
.B(n_928),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_945),
.A2(n_977),
.B(n_963),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_902),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_894),
.Y(n_1038)
);

CKINVDCx6p67_ASAP7_75t_R g1039 ( 
.A(n_929),
.Y(n_1039)
);

CKINVDCx11_ASAP7_75t_R g1040 ( 
.A(n_895),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_898),
.Y(n_1041)
);

AOI211x1_ASAP7_75t_L g1042 ( 
.A1(n_939),
.A2(n_942),
.B(n_925),
.C(n_983),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_893),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_992),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1002),
.B(n_888),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_889),
.A2(n_1009),
.B(n_970),
.C(n_934),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_911),
.A2(n_905),
.B(n_1010),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_909),
.A2(n_887),
.B(n_905),
.Y(n_1048)
);

NOR2xp67_ASAP7_75t_SL g1049 ( 
.A(n_888),
.B(n_932),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_909),
.A2(n_886),
.B(n_1009),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_1004),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_919),
.A2(n_923),
.B1(n_914),
.B2(n_908),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_901),
.A2(n_960),
.B(n_952),
.C(n_953),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1006),
.B(n_906),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_891),
.B(n_933),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_901),
.A2(n_892),
.B(n_927),
.Y(n_1056)
);

AO21x2_ASAP7_75t_L g1057 ( 
.A1(n_973),
.A2(n_951),
.B(n_971),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_952),
.A2(n_960),
.B(n_953),
.C(n_974),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_927),
.A2(n_944),
.B(n_966),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_927),
.A2(n_978),
.B(n_976),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_961),
.A2(n_896),
.B(n_973),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_914),
.B(n_933),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_962),
.Y(n_1063)
);

AO32x2_ASAP7_75t_L g1064 ( 
.A1(n_907),
.A2(n_954),
.A3(n_943),
.B1(n_919),
.B2(n_964),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1002),
.B(n_959),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_912),
.B(n_969),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_972),
.A2(n_975),
.B(n_916),
.C(n_985),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_968),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_891),
.A2(n_897),
.B1(n_910),
.B2(n_948),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_936),
.B(n_907),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_937),
.A2(n_996),
.B(n_994),
.C(n_940),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_978),
.A2(n_1012),
.B(n_956),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_SL g1073 ( 
.A1(n_926),
.A2(n_948),
.B1(n_969),
.B2(n_922),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_956),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_922),
.A2(n_984),
.B(n_967),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_921),
.B(n_957),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_937),
.B(n_940),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_947),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_956),
.A2(n_1012),
.B(n_1008),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_955),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1001),
.A2(n_618),
.B1(n_483),
.B2(n_554),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_1001),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1012),
.B(n_1001),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1008),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1008),
.B(n_982),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_993),
.A2(n_1005),
.B(n_1003),
.C(n_602),
.Y(n_1086)
);

NOR4xp25_ASAP7_75t_L g1087 ( 
.A(n_993),
.B(n_1003),
.C(n_1005),
.D(n_904),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_1006),
.B(n_809),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_993),
.A2(n_875),
.B(n_872),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_986),
.A2(n_991),
.B1(n_995),
.B2(n_988),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_904),
.A2(n_920),
.B(n_986),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_982),
.B(n_998),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_890),
.A2(n_915),
.B1(n_602),
.B2(n_982),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_997),
.B(n_453),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_986),
.A2(n_991),
.B(n_988),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_926),
.B(n_823),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_SL g1103 ( 
.A1(n_980),
.A2(n_979),
.B(n_835),
.C(n_863),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_982),
.B(n_998),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1002),
.B(n_871),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_982),
.B(n_998),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_902),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_924),
.A2(n_1015),
.B(n_1010),
.Y(n_1111)
);

AO22x2_ASAP7_75t_L g1112 ( 
.A1(n_915),
.A2(n_899),
.B1(n_1000),
.B2(n_981),
.Y(n_1112)
);

INVx6_ASAP7_75t_L g1113 ( 
.A(n_888),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_900),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_962),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_987),
.B(n_732),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_904),
.A2(n_920),
.B(n_986),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_888),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_894),
.B(n_576),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_894),
.B(n_576),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_902),
.Y(n_1123)
);

NOR4xp25_ASAP7_75t_L g1124 ( 
.A(n_993),
.B(n_1003),
.C(n_1005),
.D(n_904),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_931),
.A2(n_1015),
.B(n_949),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_902),
.Y(n_1126)
);

NOR4xp25_ASAP7_75t_L g1127 ( 
.A(n_993),
.B(n_1003),
.C(n_1005),
.D(n_904),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_1007),
.Y(n_1128)
);

INVx8_ASAP7_75t_L g1129 ( 
.A(n_1002),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_904),
.A2(n_920),
.B(n_986),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_894),
.B(n_576),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_902),
.Y(n_1132)
);

NAND3x1_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_906),
.C(n_923),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_980),
.A2(n_924),
.B(n_918),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_895),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_914),
.A2(n_618),
.B1(n_483),
.B2(n_554),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_958),
.A2(n_749),
.A3(n_918),
.B(n_920),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_902),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_904),
.A2(n_920),
.B(n_986),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_986),
.A2(n_991),
.B1(n_995),
.B2(n_988),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_989),
.A2(n_1011),
.B(n_990),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1040),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_1081),
.B2(n_1062),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1052),
.A2(n_1099),
.B1(n_1022),
.B2(n_1021),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1099),
.A2(n_1022),
.B1(n_1054),
.B2(n_1100),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1044),
.A2(n_1016),
.B1(n_1096),
.B2(n_1104),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1109),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1123),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1133),
.A2(n_1108),
.B1(n_1027),
.B2(n_1029),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_1112),
.A2(n_1033),
.B1(n_1130),
.B2(n_1118),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1126),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1135),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1023),
.A2(n_1090),
.B(n_1020),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1065),
.A2(n_1043),
.B1(n_1031),
.B2(n_1141),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1132),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1113),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1139),
.Y(n_1158)
);

CKINVDCx6p67_ASAP7_75t_R g1159 ( 
.A(n_1119),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1116),
.A2(n_1112),
.B1(n_1118),
.B2(n_1094),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1086),
.A2(n_1028),
.B1(n_1093),
.B2(n_1141),
.Y(n_1161)
);

CKINVDCx11_ASAP7_75t_R g1162 ( 
.A(n_1019),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1094),
.A2(n_1130),
.B1(n_1140),
.B2(n_1121),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1113),
.Y(n_1164)
);

BUFx2_ASAP7_75t_SL g1165 ( 
.A(n_1119),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1038),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1025),
.Y(n_1167)
);

INVx6_ASAP7_75t_L g1168 ( 
.A(n_1068),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1140),
.A2(n_1120),
.B1(n_1131),
.B2(n_1078),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1075),
.Y(n_1170)
);

CKINVDCx11_ASAP7_75t_R g1171 ( 
.A(n_1019),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1083),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1069),
.A2(n_1055),
.B1(n_1018),
.B2(n_1095),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1093),
.A2(n_1076),
.B1(n_1024),
.B2(n_1089),
.Y(n_1174)
);

INVx6_ASAP7_75t_L g1175 ( 
.A(n_1068),
.Y(n_1175)
);

INVx6_ASAP7_75t_L g1176 ( 
.A(n_1128),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1088),
.A2(n_1061),
.B1(n_1065),
.B2(n_1069),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1087),
.B(n_1124),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1114),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1042),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1061),
.A2(n_1032),
.B1(n_1057),
.B2(n_1085),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1041),
.A2(n_1087),
.B1(n_1127),
.B2(n_1124),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1084),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1057),
.A2(n_1073),
.B1(n_1066),
.B2(n_1105),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1048),
.A2(n_1050),
.B(n_1045),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1039),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1105),
.A2(n_1102),
.B1(n_1059),
.B2(n_1050),
.Y(n_1187)
);

INVx6_ASAP7_75t_L g1188 ( 
.A(n_1128),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1034),
.A2(n_1070),
.B1(n_1115),
.B2(n_1063),
.Y(n_1189)
);

CKINVDCx11_ASAP7_75t_R g1190 ( 
.A(n_1051),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1082),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1080),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1056),
.A2(n_1060),
.B1(n_1127),
.B2(n_1074),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1077),
.Y(n_1194)
);

INVx8_ASAP7_75t_L g1195 ( 
.A(n_1049),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1064),
.B(n_1030),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1101),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1047),
.A2(n_1091),
.B1(n_1137),
.B2(n_1122),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_1117),
.B1(n_1110),
.B2(n_1142),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1046),
.A2(n_1064),
.B(n_1030),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1071),
.B(n_1079),
.Y(n_1201)
);

BUFx12f_ASAP7_75t_L g1202 ( 
.A(n_1053),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1072),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1067),
.Y(n_1204)
);

INVx8_ASAP7_75t_L g1205 ( 
.A(n_1058),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1030),
.Y(n_1206)
);

INVx11_ASAP7_75t_L g1207 ( 
.A(n_1103),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1111),
.A2(n_1036),
.B1(n_1026),
.B2(n_1125),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1138),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1035),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1134),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1097),
.A2(n_1098),
.B1(n_1106),
.B2(n_1107),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1052),
.A2(n_914),
.B1(n_618),
.B2(n_298),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1113),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1052),
.A2(n_914),
.B1(n_618),
.B2(n_298),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1099),
.A2(n_602),
.B1(n_997),
.B2(n_1022),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1037),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1017),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1052),
.A2(n_914),
.B1(n_618),
.B2(n_298),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1112),
.B(n_1022),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1037),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1052),
.A2(n_914),
.B1(n_618),
.B2(n_298),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1037),
.Y(n_1226)
);

INVx8_ASAP7_75t_L g1227 ( 
.A(n_1129),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1017),
.Y(n_1228)
);

INVx6_ASAP7_75t_L g1229 ( 
.A(n_1119),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1040),
.Y(n_1230)
);

CKINVDCx6p67_ASAP7_75t_R g1231 ( 
.A(n_1119),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1099),
.A2(n_1022),
.B1(n_997),
.B2(n_1016),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1017),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1075),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1040),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1136),
.A2(n_1052),
.B1(n_618),
.B2(n_914),
.Y(n_1238)
);

BUFx4f_ASAP7_75t_SL g1239 ( 
.A(n_1039),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1052),
.A2(n_914),
.B1(n_618),
.B2(n_298),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1040),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1204),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1190),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1196),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1150),
.B(n_1155),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1196),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_R g1247 ( 
.A(n_1239),
.B(n_1190),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1193),
.A2(n_1200),
.B(n_1154),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1199),
.A2(n_1198),
.B(n_1208),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1216),
.A2(n_1146),
.B1(n_1145),
.B2(n_1163),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1209),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1220),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1209),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1206),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1178),
.B(n_1172),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1170),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1210),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1213),
.A2(n_1240),
.B1(n_1219),
.B2(n_1215),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1170),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1161),
.B(n_1151),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1152),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1167),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1156),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_R g1265 ( 
.A(n_1143),
.B(n_1153),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1158),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1217),
.B(n_1222),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1236),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1226),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1166),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1201),
.A2(n_1180),
.B(n_1185),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1232),
.A2(n_1233),
.B1(n_1221),
.B2(n_1235),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1160),
.B(n_1173),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1174),
.B(n_1169),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1236),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1211),
.A2(n_1187),
.B(n_1181),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1147),
.B(n_1194),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1223),
.A2(n_1238),
.B1(n_1225),
.B2(n_1224),
.Y(n_1278)
);

OR2x6_ASAP7_75t_L g1279 ( 
.A(n_1204),
.B(n_1173),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1184),
.A2(n_1183),
.B(n_1177),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1191),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1179),
.B(n_1228),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1203),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1203),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1189),
.A2(n_1212),
.B(n_1144),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1218),
.Y(n_1286)
);

CKINVDCx14_ASAP7_75t_R g1287 ( 
.A(n_1143),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1202),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1207),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1207),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1202),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1182),
.B(n_1205),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1197),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1197),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1159),
.A2(n_1231),
.B(n_1229),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1262),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1262),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1261),
.A2(n_1194),
.B(n_1234),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1286),
.B(n_1176),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1255),
.B(n_1192),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1255),
.B(n_1176),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1279),
.B(n_1195),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1244),
.B(n_1176),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_1270),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1272),
.A2(n_1195),
.B1(n_1153),
.B2(n_1237),
.C(n_1230),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1243),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1244),
.B(n_1188),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1272),
.A2(n_1195),
.B(n_1157),
.C(n_1164),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1246),
.B(n_1214),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1261),
.A2(n_1214),
.B(n_1164),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1290),
.B(n_1162),
.C(n_1171),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1264),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1295),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1271),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1290),
.A2(n_1165),
.B(n_1241),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1243),
.A2(n_1241),
.B1(n_1237),
.B2(n_1230),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1282),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1250),
.A2(n_1186),
.B1(n_1168),
.B2(n_1175),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1281),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1252),
.B(n_1186),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1281),
.Y(n_1321)
);

NOR3xp33_ASAP7_75t_SL g1322 ( 
.A(n_1265),
.B(n_1162),
.C(n_1171),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1271),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1250),
.A2(n_1167),
.B(n_1227),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1245),
.A2(n_1285),
.B(n_1292),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1257),
.B(n_1254),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1266),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1243),
.B(n_1287),
.Y(n_1328)
);

AO32x2_ASAP7_75t_L g1329 ( 
.A1(n_1256),
.A2(n_1260),
.A3(n_1268),
.B1(n_1242),
.B2(n_1271),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1283),
.B(n_1259),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1285),
.A2(n_1292),
.B(n_1274),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1278),
.A2(n_1274),
.B1(n_1258),
.B2(n_1277),
.C(n_1283),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1267),
.B(n_1266),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1247),
.Y(n_1335)
);

CKINVDCx6p67_ASAP7_75t_R g1336 ( 
.A(n_1288),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1296),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1319),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1297),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1332),
.A2(n_1273),
.B1(n_1248),
.B2(n_1279),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1333),
.B(n_1248),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1329),
.B(n_1248),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1321),
.B(n_1269),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1318),
.B(n_1282),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1329),
.B(n_1275),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1312),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1329),
.B(n_1275),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1329),
.B(n_1275),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1327),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1304),
.B(n_1269),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1325),
.A2(n_1273),
.B1(n_1293),
.B2(n_1294),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1334),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1326),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1329),
.B(n_1249),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1326),
.Y(n_1355)
);

OAI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1331),
.A2(n_1289),
.B(n_1294),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1317),
.B(n_1330),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1314),
.B(n_1284),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1305),
.A2(n_1279),
.B1(n_1253),
.B2(n_1251),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1317),
.B(n_1249),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1323),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1315),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1300),
.B(n_1289),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1300),
.B(n_1254),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1309),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1337),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1342),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1337),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1337),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1338),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1341),
.B(n_1303),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_SL g1373 ( 
.A(n_1342),
.B(n_1302),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1345),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1341),
.B(n_1307),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1356),
.B(n_1336),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1342),
.B(n_1313),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1356),
.B(n_1336),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1339),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1345),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1339),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1363),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1338),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1345),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1353),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1340),
.A2(n_1298),
.B1(n_1279),
.B2(n_1324),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1347),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1363),
.B(n_1313),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1347),
.B(n_1301),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1353),
.B(n_1320),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1363),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1344),
.B(n_1320),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1340),
.A2(n_1293),
.B1(n_1276),
.B2(n_1280),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1351),
.A2(n_1308),
.B(n_1315),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1351),
.A2(n_1293),
.B1(n_1302),
.B2(n_1310),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1354),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1354),
.A2(n_1288),
.B1(n_1291),
.B2(n_1306),
.C(n_1311),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1347),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1348),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1390),
.B(n_1355),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1371),
.B(n_1352),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1396),
.B(n_1366),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1371),
.B(n_1367),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1367),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1369),
.B(n_1346),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1387),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1396),
.B(n_1372),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1369),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1390),
.B(n_1374),
.Y(n_1409)
);

AND2x2_ASAP7_75t_SL g1410 ( 
.A(n_1391),
.B(n_1354),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1396),
.B(n_1366),
.Y(n_1411)
);

OAI33xp33_ASAP7_75t_L g1412 ( 
.A1(n_1388),
.A2(n_1362),
.A3(n_1359),
.B1(n_1350),
.B2(n_1343),
.B3(n_1383),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1396),
.B(n_1348),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1370),
.B(n_1349),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1370),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1396),
.B(n_1372),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1379),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1392),
.B(n_1335),
.Y(n_1418)
);

INVx8_ASAP7_75t_L g1419 ( 
.A(n_1383),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1390),
.B(n_1365),
.Y(n_1420)
);

NOR2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1387),
.B(n_1306),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1382),
.B(n_1315),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1396),
.B(n_1364),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1391),
.B(n_1348),
.Y(n_1424)
);

OAI33xp33_ASAP7_75t_L g1425 ( 
.A1(n_1388),
.A2(n_1359),
.A3(n_1362),
.B1(n_1350),
.B2(n_1343),
.B3(n_1358),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1396),
.B(n_1357),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1381),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1381),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1394),
.B(n_1376),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1387),
.B(n_1361),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1387),
.B(n_1361),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1430),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1415),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1401),
.B(n_1392),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1420),
.B(n_1374),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1415),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1419),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1420),
.B(n_1374),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1404),
.Y(n_1441)
);

OAI31xp33_ASAP7_75t_L g1442 ( 
.A1(n_1429),
.A2(n_1397),
.A3(n_1422),
.B(n_1377),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1400),
.B(n_1385),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1400),
.B(n_1361),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1418),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1419),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1404),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1408),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1410),
.B(n_1389),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1408),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1417),
.Y(n_1453)
);

AND2x4_ASAP7_75t_SL g1454 ( 
.A(n_1407),
.B(n_1322),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1413),
.A2(n_1394),
.B(n_1397),
.C(n_1395),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1417),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1403),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_SL g1461 ( 
.A(n_1424),
.B(n_1391),
.C(n_1378),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1413),
.B(n_1295),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1427),
.Y(n_1464)
);

AOI32xp33_ASAP7_75t_L g1465 ( 
.A1(n_1430),
.A2(n_1382),
.A3(n_1398),
.B1(n_1399),
.B2(n_1380),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1430),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1425),
.A2(n_1368),
.B1(n_1398),
.B2(n_1380),
.C(n_1399),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1428),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1405),
.Y(n_1470)
);

NAND2x1_ASAP7_75t_L g1471 ( 
.A(n_1402),
.B(n_1374),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1403),
.B(n_1382),
.C(n_1362),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1432),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1450),
.B(n_1407),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1435),
.B(n_1409),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1450),
.B(n_1416),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1437),
.B(n_1416),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1433),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1439),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1460),
.B(n_1380),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1433),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1445),
.B(n_1470),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1434),
.B(n_1409),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1454),
.B(n_1426),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1437),
.B(n_1382),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1456),
.A2(n_1386),
.B1(n_1393),
.B2(n_1412),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1438),
.B(n_1380),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.B(n_1426),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1446),
.B(n_1431),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1422),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.Y(n_1493)
);

BUFx2_ASAP7_75t_SL g1494 ( 
.A(n_1447),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1451),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1436),
.B(n_1405),
.Y(n_1496)
);

XNOR2x2_ASAP7_75t_L g1497 ( 
.A(n_1473),
.B(n_1395),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1439),
.B(n_1402),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1451),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1442),
.A2(n_1424),
.B(n_1419),
.C(n_1378),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1452),
.B(n_1411),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1452),
.B(n_1411),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1436),
.B(n_1414),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1441),
.B(n_1384),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1455),
.B(n_1422),
.Y(n_1505)
);

INVx5_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1448),
.B(n_1384),
.Y(n_1508)
);

OAI31xp33_ASAP7_75t_L g1509 ( 
.A1(n_1500),
.A2(n_1456),
.A3(n_1422),
.B(n_1462),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1488),
.A2(n_1467),
.B(n_1465),
.C(n_1461),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1316),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1443),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1488),
.A2(n_1376),
.B(n_1455),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1485),
.B(n_1458),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1505),
.A2(n_1412),
.B1(n_1425),
.B2(n_1393),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1483),
.A2(n_1468),
.B(n_1464),
.C(n_1471),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1477),
.A2(n_1472),
.B1(n_1463),
.B2(n_1384),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1506),
.B(n_1462),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1494),
.B(n_1479),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1485),
.B(n_1423),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1492),
.A2(n_1486),
.B(n_1263),
.Y(n_1521)
);

NOR4xp25_ASAP7_75t_L g1522 ( 
.A(n_1497),
.B(n_1468),
.C(n_1469),
.D(n_1457),
.Y(n_1522)
);

AOI31xp33_ASAP7_75t_L g1523 ( 
.A1(n_1490),
.A2(n_1335),
.A3(n_1328),
.B(n_1462),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1476),
.B(n_1449),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1497),
.A2(n_1360),
.B1(n_1386),
.B2(n_1440),
.C(n_1431),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1479),
.A2(n_1471),
.B(n_1459),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1506),
.A2(n_1368),
.B1(n_1399),
.B2(n_1384),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1506),
.B(n_1406),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1476),
.B(n_1453),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1484),
.B(n_1440),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1477),
.A2(n_1398),
.B1(n_1399),
.B2(n_1368),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1495),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1528),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1511),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1533),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1494),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1522),
.B(n_1479),
.Y(n_1539)
);

AOI322xp5_ASAP7_75t_L g1540 ( 
.A1(n_1515),
.A2(n_1481),
.A3(n_1505),
.B1(n_1398),
.B2(n_1444),
.C1(n_1368),
.C2(n_1431),
.Y(n_1540)
);

AOI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1519),
.A2(n_1487),
.B(n_1482),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1524),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1530),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1531),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

NAND2x1_ASAP7_75t_L g1546 ( 
.A(n_1521),
.B(n_1490),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1509),
.B(n_1506),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1506),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1519),
.B(n_1498),
.Y(n_1550)
);

AOI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1513),
.A2(n_1487),
.B(n_1482),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1523),
.A2(n_1368),
.B1(n_1506),
.B2(n_1492),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1544),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1538),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1535),
.B(n_1537),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_1484),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1537),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1547),
.A2(n_1510),
.B1(n_1525),
.B2(n_1516),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1538),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1534),
.Y(n_1560)
);

OA22x2_ASAP7_75t_L g1561 ( 
.A1(n_1547),
.A2(n_1526),
.B1(n_1486),
.B2(n_1477),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1548),
.B(n_1482),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1548),
.B(n_1487),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1536),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1557),
.B(n_1550),
.Y(n_1565)
);

AOI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1556),
.A2(n_1541),
.B(n_1551),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1554),
.Y(n_1567)
);

NAND4xp25_ASAP7_75t_L g1568 ( 
.A(n_1555),
.B(n_1549),
.C(n_1545),
.D(n_1550),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1558),
.A2(n_1540),
.B(n_1546),
.C(n_1543),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1559),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1562),
.B(n_1546),
.Y(n_1571)
);

NOR3xp33_ASAP7_75t_L g1572 ( 
.A(n_1558),
.B(n_1542),
.C(n_1552),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1563),
.B(n_1493),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1565),
.Y(n_1574)
);

AOI311xp33_ASAP7_75t_L g1575 ( 
.A1(n_1572),
.A2(n_1553),
.A3(n_1560),
.B(n_1564),
.C(n_1561),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1569),
.B(n_1493),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_L g1577 ( 
.A(n_1571),
.B(n_1568),
.C(n_1566),
.D(n_1567),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_SL g1578 ( 
.A(n_1570),
.B(n_1518),
.C(n_1529),
.Y(n_1578)
);

AOI222xp33_ASAP7_75t_L g1579 ( 
.A1(n_1576),
.A2(n_1573),
.B1(n_1499),
.B2(n_1507),
.C1(n_1493),
.C2(n_1527),
.Y(n_1579)
);

AOI211xp5_ASAP7_75t_L g1580 ( 
.A1(n_1577),
.A2(n_1527),
.B(n_1517),
.C(n_1532),
.Y(n_1580)
);

AOI222xp33_ASAP7_75t_L g1581 ( 
.A1(n_1578),
.A2(n_1507),
.B1(n_1499),
.B2(n_1481),
.C1(n_1368),
.C2(n_1489),
.Y(n_1581)
);

NOR3xp33_ASAP7_75t_L g1582 ( 
.A(n_1574),
.B(n_1489),
.C(n_1486),
.Y(n_1582)
);

XNOR2xp5_ASAP7_75t_L g1583 ( 
.A(n_1575),
.B(n_1486),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1578),
.A2(n_1477),
.B(n_1475),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1583),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1584),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1582),
.B(n_1496),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1581),
.B(n_1579),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1580),
.A2(n_1492),
.B1(n_1475),
.B2(n_1478),
.Y(n_1589)
);

XNOR2x1_ASAP7_75t_L g1590 ( 
.A(n_1586),
.B(n_1492),
.Y(n_1590)
);

NOR3xp33_ASAP7_75t_SL g1591 ( 
.A(n_1588),
.B(n_1585),
.C(n_1587),
.Y(n_1591)
);

XOR2xp5_ASAP7_75t_L g1592 ( 
.A(n_1589),
.B(n_1373),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1591),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1593),
.Y(n_1594)
);

INVxp33_ASAP7_75t_SL g1595 ( 
.A(n_1594),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1594),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1595),
.B(n_1590),
.Y(n_1597)
);

OA22x2_ASAP7_75t_L g1598 ( 
.A1(n_1596),
.A2(n_1592),
.B1(n_1492),
.B2(n_1478),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1597),
.A2(n_1508),
.B(n_1504),
.Y(n_1599)
);

OAI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1598),
.A2(n_1503),
.B1(n_1496),
.B2(n_1508),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1599),
.A2(n_1504),
.B(n_1503),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1601),
.B(n_1600),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1602),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_R g1604 ( 
.A1(n_1603),
.A2(n_1478),
.B1(n_1491),
.B2(n_1501),
.C(n_1502),
.Y(n_1604)
);

AOI211xp5_ASAP7_75t_L g1605 ( 
.A1(n_1604),
.A2(n_1478),
.B(n_1299),
.C(n_1502),
.Y(n_1605)
);


endmodule