module fake_jpeg_12623_n_549 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_549);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_3),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_112),
.Y(n_132)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_65),
.Y(n_185)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_21),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_68),
.A2(n_107),
.B1(n_32),
.B2(n_38),
.Y(n_175)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_98),
.Y(n_130)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g174 ( 
.A(n_73),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_79),
.B(n_87),
.Y(n_176)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_8),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_90),
.B(n_100),
.Y(n_151)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_27),
.B(n_30),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_10),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_30),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_111),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_31),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_33),
.B(n_16),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_28),
.Y(n_155)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_126),
.B(n_142),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_66),
.A2(n_31),
.B1(n_43),
.B2(n_56),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_139),
.A2(n_145),
.B1(n_181),
.B2(n_184),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_89),
.A2(n_31),
.B1(n_96),
.B2(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_148),
.B(n_165),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_44),
.C(n_40),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_32),
.B(n_45),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_61),
.B(n_53),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_161),
.B(n_163),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_36),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_48),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_57),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_166),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_175),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_94),
.A2(n_56),
.B1(n_57),
.B2(n_28),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_99),
.A2(n_56),
.B1(n_50),
.B2(n_38),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_113),
.A2(n_28),
.B1(n_108),
.B2(n_117),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_187),
.A2(n_6),
.B1(n_16),
.B2(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_49),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_193),
.B(n_196),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_73),
.A2(n_49),
.B(n_58),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_48),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_65),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_63),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_85),
.A2(n_58),
.B1(n_36),
.B2(n_42),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_50),
.B1(n_45),
.B2(n_22),
.Y(n_226)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_206),
.Y(n_315)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_209),
.B(n_145),
.Y(n_284)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_130),
.B(n_42),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_77),
.B1(n_75),
.B2(n_74),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_216),
.A2(n_252),
.B1(n_260),
.B2(n_190),
.Y(n_294)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_217),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_132),
.A2(n_40),
.B(n_29),
.C(n_54),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_228),
.Y(n_277)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

BUFx6f_ASAP7_75t_SL g221 ( 
.A(n_156),
.Y(n_221)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_225),
.Y(n_296)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_151),
.A2(n_54),
.B1(n_52),
.B2(n_29),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_224),
.A2(n_235),
.B1(n_266),
.B2(n_268),
.Y(n_305)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_226),
.A2(n_183),
.B1(n_197),
.B2(n_149),
.Y(n_286)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_133),
.A2(n_52),
.B(n_22),
.C(n_28),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_146),
.Y(n_230)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_131),
.Y(n_231)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_0),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_232),
.B(n_249),
.Y(n_283)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_149),
.Y(n_234)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_167),
.A2(n_67),
.B1(n_59),
.B2(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_147),
.Y(n_240)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_137),
.Y(n_242)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_244),
.Y(n_274)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_245),
.A2(n_185),
.B1(n_268),
.B2(n_226),
.Y(n_307)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_6),
.A3(n_12),
.B1(n_16),
.B2(n_1),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_247),
.Y(n_293)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_248),
.A2(n_194),
.B1(n_189),
.B2(n_141),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_138),
.B(n_1),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_253),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_187),
.A2(n_6),
.B1(n_16),
.B2(n_4),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_128),
.B(n_1),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_129),
.B(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_256),
.Y(n_279)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_257),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_136),
.B(n_1),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_258),
.B(n_262),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_156),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_259),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_181),
.A2(n_3),
.B1(n_4),
.B2(n_139),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_154),
.B(n_3),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_269),
.Y(n_288)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_177),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_265),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_191),
.A2(n_4),
.B1(n_135),
.B2(n_140),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_267),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_188),
.B(n_173),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_191),
.A2(n_135),
.B1(n_140),
.B2(n_152),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_270),
.A2(n_271),
.B1(n_220),
.B2(n_217),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_152),
.A2(n_189),
.B1(n_171),
.B2(n_182),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_236),
.B(n_155),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_282),
.A2(n_292),
.B(n_281),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_208),
.C(n_243),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_307),
.B1(n_317),
.B2(n_208),
.Y(n_339)
);

AO21x2_ASAP7_75t_L g289 ( 
.A1(n_232),
.A2(n_215),
.B(n_216),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_236),
.A2(n_194),
.B(n_141),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_205),
.A2(n_160),
.B1(n_190),
.B2(n_199),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_171),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_299),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_199),
.B1(n_197),
.B2(n_183),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_218),
.B(n_143),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_241),
.B(n_178),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_302),
.B(n_244),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_259),
.B1(n_221),
.B2(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_228),
.B(n_160),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_320),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_245),
.A2(n_185),
.B1(n_209),
.B2(n_233),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_276),
.B1(n_309),
.B2(n_273),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_249),
.A2(n_229),
.B1(n_234),
.B2(n_207),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_255),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_204),
.C(n_211),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_300),
.C(n_313),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_326),
.A2(n_351),
.B1(n_301),
.B2(n_291),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_267),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_328),
.B(n_335),
.Y(n_379)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_289),
.A2(n_212),
.B1(n_227),
.B2(n_223),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_338),
.B1(n_353),
.B2(n_355),
.Y(n_369)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_321),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_334),
.B(n_340),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_277),
.B(n_206),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_213),
.B(n_210),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_337),
.A2(n_348),
.B(n_349),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_289),
.A2(n_265),
.B1(n_219),
.B2(n_250),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_339),
.A2(n_350),
.B1(n_357),
.B2(n_362),
.Y(n_390)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_258),
.B1(n_262),
.B2(n_240),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_247),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_342),
.B(n_318),
.Y(n_385)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_296),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_346),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_296),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_231),
.B(n_257),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_294),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_286),
.B1(n_304),
.B2(n_303),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

INVx11_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_289),
.A2(n_314),
.B1(n_277),
.B2(n_293),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_274),
.B(n_323),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_288),
.A2(n_305),
.B1(n_283),
.B2(n_279),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_288),
.A2(n_283),
.B1(n_279),
.B2(n_317),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_358),
.B1(n_359),
.B2(n_364),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_282),
.A2(n_308),
.B1(n_312),
.B2(n_278),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_278),
.A2(n_308),
.B1(n_312),
.B2(n_290),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_351),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_285),
.B(n_287),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_363),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_285),
.A2(n_290),
.B1(n_273),
.B2(n_287),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_272),
.A2(n_280),
.B1(n_319),
.B2(n_322),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_315),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_350),
.A2(n_272),
.B1(n_319),
.B2(n_311),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_327),
.B1(n_349),
.B2(n_332),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_368),
.B(n_389),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_361),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_335),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_311),
.B1(n_316),
.B2(n_300),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_393),
.B1(n_339),
.B2(n_362),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_386),
.C(n_387),
.Y(n_404)
);

XOR2x2_ASAP7_75t_L g384 ( 
.A(n_341),
.B(n_301),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_396),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_385),
.B(n_357),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_310),
.C(n_313),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_316),
.C(n_318),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_301),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_346),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_391),
.B(n_328),
.Y(n_407)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_327),
.A2(n_353),
.B1(n_338),
.B2(n_331),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_315),
.Y(n_394)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_395),
.A2(n_337),
.B(n_348),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_291),
.C(n_355),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_330),
.B(n_291),
.Y(n_398)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_398),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_347),
.C(n_354),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_363),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_392),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_409),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_421),
.B1(n_422),
.B2(n_371),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_407),
.B(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_384),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_408),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_366),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_411),
.A2(n_415),
.B1(n_418),
.B2(n_369),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_376),
.A2(n_347),
.B(n_342),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_419),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_329),
.B(n_354),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_424),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_390),
.A2(n_367),
.B1(n_399),
.B2(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_349),
.B1(n_340),
.B2(n_354),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_334),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_428),
.C(n_386),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_393),
.A2(n_340),
.B1(n_336),
.B2(n_344),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_369),
.A2(n_344),
.B1(n_343),
.B2(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_366),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_372),
.B(n_359),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_427),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_435),
.Y(n_464)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_427),
.B(n_396),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_434),
.B(n_410),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_389),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_436),
.A2(n_447),
.B1(n_448),
.B2(n_419),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_384),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_441),
.C(n_443),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_424),
.Y(n_439)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_415),
.A2(n_383),
.B1(n_370),
.B2(n_395),
.Y(n_442)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_382),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_387),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_449),
.C(n_450),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_418),
.A2(n_383),
.B1(n_380),
.B2(n_388),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_411),
.A2(n_380),
.B1(n_388),
.B2(n_394),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_398),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_381),
.C(n_365),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_403),
.B1(n_422),
.B2(n_413),
.Y(n_452)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_466),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_457),
.A2(n_471),
.B1(n_472),
.B2(n_459),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_430),
.A2(n_444),
.B(n_412),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_458),
.A2(n_469),
.B(n_470),
.Y(n_480)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_453),
.Y(n_462)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_385),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_467),
.Y(n_481)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_402),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_379),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_379),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_449),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_430),
.A2(n_414),
.B(n_405),
.Y(n_469)
);

XOR2x2_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_434),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_417),
.B(n_410),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_377),
.B(n_360),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_447),
.A2(n_413),
.B1(n_400),
.B2(n_417),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_451),
.A2(n_400),
.B1(n_423),
.B2(n_416),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_SL g473 ( 
.A(n_450),
.B(n_426),
.C(n_377),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_477),
.CI(n_466),
.CON(n_487),
.SN(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_476),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_397),
.C(n_374),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_474),
.C(n_441),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_479),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_480),
.A2(n_490),
.B(n_493),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_494),
.C(n_495),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_484),
.A2(n_485),
.B1(n_488),
.B2(n_491),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_452),
.B1(n_433),
.B2(n_448),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_443),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_487),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_454),
.B1(n_432),
.B2(n_438),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_457),
.A2(n_445),
.B1(n_431),
.B2(n_397),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_374),
.C(n_364),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_352),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_490),
.B(n_458),
.CI(n_459),
.CON(n_497),
.SN(n_497)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_497),
.B(n_490),
.CI(n_489),
.CON(n_520),
.SN(n_520)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_455),
.B1(n_460),
.B2(n_471),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_498),
.A2(n_508),
.B1(n_497),
.B2(n_507),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_464),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_502),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_475),
.C(n_464),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_504),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_456),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_481),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_485),
.A2(n_455),
.B1(n_460),
.B2(n_462),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_478),
.B1(n_472),
.B2(n_494),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_465),
.Y(n_507)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_507),
.Y(n_513)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_482),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_506),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_505),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_502),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_488),
.B(n_493),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_517),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_495),
.C(n_473),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_499),
.C(n_496),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_506),
.B(n_500),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_519),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_521),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_500),
.A2(n_467),
.B1(n_482),
.B2(n_492),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g522 ( 
.A1(n_515),
.A2(n_504),
.B(n_503),
.Y(n_522)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_522),
.A2(n_525),
.B(n_526),
.C(n_521),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_501),
.Y(n_523)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_523),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_503),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_524),
.B(n_513),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_529),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_498),
.Y(n_533)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_531),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_532),
.A2(n_537),
.B(n_526),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_534),
.C(n_535),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_529),
.B(n_514),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_514),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_538),
.A2(n_540),
.B(n_489),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_536),
.A2(n_525),
.B(n_512),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g544 ( 
.A(n_541),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_539),
.A2(n_533),
.B(n_492),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_542),
.A2(n_543),
.B(n_497),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_544),
.C(n_499),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_502),
.C(n_487),
.Y(n_547)
);

MAJx2_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_487),
.C(n_497),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_520),
.B(n_545),
.Y(n_549)
);


endmodule