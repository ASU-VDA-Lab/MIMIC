module fake_jpeg_20212_n_279 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_24),
.C(n_21),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_21),
.C(n_25),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_13),
.B1(n_16),
.B2(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_15),
.Y(n_55)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_34),
.B1(n_13),
.B2(n_16),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_14),
.B1(n_38),
.B2(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_28),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_69),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_71),
.B(n_21),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_45),
.B(n_24),
.C(n_16),
.Y(n_79)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_44),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_66),
.C(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_41),
.B1(n_48),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_83),
.B1(n_92),
.B2(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_66),
.B1(n_56),
.B2(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_48),
.B1(n_45),
.B2(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_88),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_37),
.B(n_14),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_55),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_69),
.Y(n_95)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_71),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_87),
.Y(n_98)
);

XNOR2x2_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_62),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_110),
.B1(n_79),
.B2(n_78),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_68),
.B1(n_67),
.B2(n_51),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_66),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_79),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_124),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_90),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_81),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_94),
.B1(n_104),
.B2(n_106),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_107),
.B(n_100),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_72),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_98),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_86),
.B(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_84),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_103),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_19),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_160),
.B1(n_38),
.B2(n_36),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_156),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_136),
.B(n_123),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_80),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_152),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_80),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_83),
.C(n_89),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_30),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_74),
.B(n_1),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_159),
.B(n_115),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_133),
.B(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_74),
.B1(n_67),
.B2(n_51),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_35),
.C(n_44),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_177),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_135),
.B(n_122),
.C(n_129),
.Y(n_165)
);

NOR4xp25_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_114),
.C(n_131),
.D(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_152),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_114),
.B(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_183),
.B1(n_20),
.B2(n_22),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_116),
.B(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_119),
.B1(n_116),
.B2(n_38),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_148),
.B1(n_146),
.B2(n_141),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_119),
.B1(n_31),
.B2(n_36),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_159),
.B1(n_146),
.B2(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_184),
.B1(n_29),
.B2(n_17),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_19),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_154),
.C(n_158),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_138),
.B(n_20),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_182),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_194),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_191),
.B1(n_206),
.B2(n_176),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_141),
.B1(n_148),
.B2(n_33),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_35),
.C(n_30),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_35),
.C(n_19),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_15),
.C(n_26),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_15),
.C(n_22),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_15),
.C(n_20),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_15),
.C(n_20),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_170),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_181),
.B1(n_165),
.B2(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_163),
.C(n_177),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_219),
.C(n_221),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_183),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_176),
.B1(n_168),
.B2(n_178),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_222),
.B1(n_187),
.B2(n_201),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_199),
.B(n_178),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_17),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_168),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_214),
.B1(n_215),
.B2(n_212),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_188),
.C(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_236),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_213),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_197),
.C(n_17),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_0),
.C(n_1),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_214),
.B(n_219),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_12),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_237),
.B1(n_225),
.B2(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_12),
.C(n_11),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_11),
.C(n_29),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_248),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_0),
.B(n_1),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_236),
.B(n_233),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_258),
.B(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_228),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_230),
.C(n_228),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_259),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_263),
.B(n_264),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_224),
.B(n_1),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_0),
.B(n_2),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_0),
.B(n_2),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_267)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_250),
.C(n_252),
.D(n_4),
.Y(n_266)
);

OAI321xp33_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_267),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_4),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.A3(n_268),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_6),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_269),
.B1(n_7),
.B2(n_9),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_6),
.B(n_9),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_278),
.Y(n_279)
);


endmodule